magic
tech sky130B
magscale 1 2
timestamp 1669668395
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 283834 700272 283840 700324
rect 283892 700312 283898 700324
rect 304994 700312 305000 700324
rect 283892 700284 305000 700312
rect 283892 700272 283898 700284
rect 304994 700272 305000 700284
rect 305052 700272 305058 700324
rect 340138 700272 340144 700324
rect 340196 700312 340202 700324
rect 348786 700312 348792 700324
rect 340196 700284 348792 700312
rect 340196 700272 340202 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 403618 700272 403624 700324
rect 403676 700312 403682 700324
rect 413646 700312 413652 700324
rect 403676 700284 413652 700312
rect 403676 700272 403682 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 414658 700272 414664 700324
rect 414716 700312 414722 700324
rect 478506 700312 478512 700324
rect 414716 700284 478512 700312
rect 414716 700272 414722 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 154114 700068 154120 700120
rect 154172 700108 154178 700120
rect 155218 700108 155224 700120
rect 154172 700080 155224 700108
rect 154172 700068 154178 700080
rect 155218 700068 155224 700080
rect 155276 700068 155282 700120
rect 8110 699660 8116 699712
rect 8168 699700 8174 699712
rect 10318 699700 10324 699712
rect 8168 699672 10324 699700
rect 8168 699660 8174 699672
rect 10318 699660 10324 699672
rect 10376 699660 10382 699712
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 26878 699700 26884 699712
rect 24360 699672 26884 699700
rect 24360 699660 24366 699672
rect 26878 699660 26884 699672
rect 26936 699660 26942 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 90358 699700 90364 699712
rect 89220 699672 90364 699700
rect 89220 699660 89226 699672
rect 90358 699660 90364 699672
rect 90416 699660 90422 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 526438 699660 526444 699712
rect 526496 699700 526502 699712
rect 527174 699700 527180 699712
rect 526496 699672 527180 699700
rect 526496 699660 526502 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 218974 698912 218980 698964
rect 219032 698952 219038 698964
rect 306374 698952 306380 698964
rect 219032 698924 306380 698952
rect 219032 698912 219038 698924
rect 306374 698912 306380 698924
rect 306432 698912 306438 698964
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 299658 696940 299664 696992
rect 299716 696980 299722 696992
rect 580166 696980 580172 696992
rect 299716 696952 580172 696980
rect 299716 696940 299722 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 300118 683204 300124 683256
rect 300176 683244 300182 683256
rect 580166 683244 580172 683256
rect 300176 683216 580172 683244
rect 300176 683204 300182 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 310514 683176 310520 683188
rect 3476 683148 310520 683176
rect 3476 683136 3482 683148
rect 310514 683136 310520 683148
rect 310572 683136 310578 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 310606 670732 310612 670744
rect 3568 670704 310612 670732
rect 3568 670692 3574 670704
rect 310606 670692 310612 670704
rect 310664 670692 310670 670744
rect 330478 670692 330484 670744
rect 330536 670732 330542 670744
rect 580166 670732 580172 670744
rect 330536 670704 580172 670732
rect 330536 670692 330542 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 310698 656928 310704 656940
rect 3476 656900 310704 656928
rect 3476 656888 3482 656900
rect 310698 656888 310704 656900
rect 310756 656888 310762 656940
rect 323578 643084 323584 643136
rect 323636 643124 323642 643136
rect 580166 643124 580172 643136
rect 323636 643096 580172 643124
rect 323636 643084 323642 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 289078 632108 289084 632120
rect 3476 632080 289084 632108
rect 3476 632068 3482 632080
rect 289078 632068 289084 632080
rect 289136 632068 289142 632120
rect 298738 630640 298744 630692
rect 298796 630680 298802 630692
rect 580166 630680 580172 630692
rect 298796 630652 580172 630680
rect 298796 630640 298802 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 302878 618304 302884 618316
rect 3200 618276 302884 618304
rect 3200 618264 3206 618276
rect 302878 618264 302884 618276
rect 302936 618264 302942 618316
rect 363598 616836 363604 616888
rect 363656 616876 363662 616888
rect 580166 616876 580172 616888
rect 363656 616848 580172 616876
rect 363656 616836 363662 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 291838 605860 291844 605872
rect 3292 605832 291844 605860
rect 3292 605820 3298 605832
rect 291838 605820 291844 605832
rect 291896 605820 291902 605872
rect 324958 590656 324964 590708
rect 325016 590696 325022 590708
rect 579798 590696 579804 590708
rect 325016 590668 579804 590696
rect 325016 590656 325022 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 334618 576852 334624 576904
rect 334676 576892 334682 576904
rect 580166 576892 580172 576904
rect 334676 576864 580172 576892
rect 334676 576852 334682 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 313274 565876 313280 565888
rect 3292 565848 313280 565876
rect 3292 565836 3298 565848
rect 313274 565836 313280 565848
rect 313332 565836 313338 565888
rect 319438 563048 319444 563100
rect 319496 563088 319502 563100
rect 579798 563088 579804 563100
rect 319496 563060 579804 563088
rect 319496 563048 319502 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 46198 553432 46204 553444
rect 3384 553404 46204 553432
rect 3384 553392 3390 553404
rect 46198 553392 46204 553404
rect 46256 553392 46262 553444
rect 320818 536800 320824 536852
rect 320876 536840 320882 536852
rect 580166 536840 580172 536852
rect 320876 536812 580172 536840
rect 320876 536800 320882 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2774 527144 2780 527196
rect 2832 527184 2838 527196
rect 4798 527184 4804 527196
rect 2832 527156 4804 527184
rect 2832 527144 2838 527156
rect 4798 527144 4804 527156
rect 4856 527144 4862 527196
rect 329098 524424 329104 524476
rect 329156 524464 329162 524476
rect 580166 524464 580172 524476
rect 329156 524436 580172 524464
rect 329156 524424 329162 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 250438 514808 250444 514820
rect 3568 514780 250444 514808
rect 3568 514768 3574 514780
rect 250438 514768 250444 514780
rect 250496 514768 250502 514820
rect 318058 510620 318064 510672
rect 318116 510660 318122 510672
rect 580166 510660 580172 510672
rect 318116 510632 580172 510660
rect 318116 510620 318122 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 14458 501004 14464 501016
rect 3108 500976 14464 501004
rect 3108 500964 3114 500976
rect 14458 500964 14464 500976
rect 14516 500964 14522 501016
rect 322198 484372 322204 484424
rect 322256 484412 322262 484424
rect 580166 484412 580172 484424
rect 322256 484384 580172 484412
rect 322256 484372 322262 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 7558 474756 7564 474768
rect 3108 474728 7564 474756
rect 3108 474716 3114 474728
rect 7558 474716 7564 474728
rect 7616 474716 7622 474768
rect 399478 470568 399484 470620
rect 399536 470608 399542 470620
rect 579982 470608 579988 470620
rect 399536 470580 579988 470608
rect 399536 470568 399542 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 314746 462380 314752 462392
rect 3568 462352 314752 462380
rect 3568 462340 3574 462352
rect 314746 462340 314752 462352
rect 314804 462340 314810 462392
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 15838 448576 15844 448588
rect 3200 448548 15844 448576
rect 3200 448536 3206 448548
rect 15838 448536 15844 448548
rect 15896 448536 15902 448588
rect 295978 447788 295984 447840
rect 296036 447828 296042 447840
rect 399478 447828 399484 447840
rect 296036 447800 399484 447828
rect 296036 447788 296042 447800
rect 399478 447788 399484 447800
rect 399536 447788 399542 447840
rect 294598 430584 294604 430636
rect 294656 430624 294662 430636
rect 579890 430624 579896 430636
rect 294656 430596 579896 430624
rect 294656 430584 294662 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 151078 422328 151084 422340
rect 3568 422300 151084 422328
rect 3568 422288 3574 422300
rect 151078 422288 151084 422300
rect 151136 422288 151142 422340
rect 294690 418140 294696 418192
rect 294748 418180 294754 418192
rect 580166 418180 580172 418192
rect 294748 418152 580172 418180
rect 294748 418140 294754 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 309594 409884 309600 409896
rect 2924 409856 309600 409884
rect 2924 409844 2930 409856
rect 309594 409844 309600 409856
rect 309652 409844 309658 409896
rect 26878 407736 26884 407788
rect 26936 407776 26942 407788
rect 309134 407776 309140 407788
rect 26936 407748 309140 407776
rect 26936 407736 26942 407748
rect 309134 407736 309140 407748
rect 309192 407736 309198 407788
rect 250438 406376 250444 406428
rect 250496 406416 250502 406428
rect 314838 406416 314844 406428
rect 250496 406388 314844 406416
rect 250496 406376 250502 406388
rect 314838 406376 314844 406388
rect 314896 406376 314902 406428
rect 294782 404336 294788 404388
rect 294840 404376 294846 404388
rect 580166 404376 580172 404388
rect 294840 404348 580172 404376
rect 294840 404336 294846 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 309594 403588 309600 403640
rect 309652 403628 309658 403640
rect 316034 403628 316040 403640
rect 309652 403600 316040 403628
rect 309652 403588 309658 403600
rect 316034 403588 316040 403600
rect 316092 403588 316098 403640
rect 304258 402228 304264 402280
rect 304316 402268 304322 402280
rect 340138 402268 340144 402280
rect 304316 402240 340144 402268
rect 304316 402228 304322 402240
rect 340138 402228 340144 402240
rect 340196 402228 340202 402280
rect 302970 400868 302976 400920
rect 303028 400908 303034 400920
rect 414658 400908 414664 400920
rect 303028 400880 414664 400908
rect 303028 400868 303034 400880
rect 414658 400868 414664 400880
rect 414716 400868 414722 400920
rect 298830 399440 298836 399492
rect 298888 399480 298894 399492
rect 334618 399480 334624 399492
rect 298888 399452 334624 399480
rect 298888 399440 298894 399452
rect 334618 399440 334624 399452
rect 334676 399440 334682 399492
rect 304350 398080 304356 398132
rect 304408 398120 304414 398132
rect 403618 398120 403624 398132
rect 304408 398092 403624 398120
rect 304408 398080 304414 398092
rect 403618 398080 403624 398092
rect 403676 398080 403682 398132
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 305638 397508 305644 397520
rect 3568 397480 305644 397508
rect 3568 397468 3574 397480
rect 305638 397468 305644 397480
rect 305696 397468 305702 397520
rect 297358 396720 297364 396772
rect 297416 396760 297422 396772
rect 329098 396760 329104 396772
rect 297416 396732 329104 396760
rect 297416 396720 297422 396732
rect 329098 396720 329104 396732
rect 329156 396720 329162 396772
rect 302878 395360 302884 395412
rect 302936 395400 302942 395412
rect 311894 395400 311900 395412
rect 302936 395372 311900 395400
rect 302936 395360 302942 395372
rect 311894 395360 311900 395372
rect 311952 395360 311958 395412
rect 14458 395292 14464 395344
rect 14516 395332 14522 395344
rect 313366 395332 313372 395344
rect 14516 395304 313372 395332
rect 14516 395292 14522 395304
rect 313366 395292 313372 395304
rect 313424 395292 313430 395344
rect 201494 394000 201500 394052
rect 201552 394040 201558 394052
rect 306466 394040 306472 394052
rect 201552 394012 306472 394040
rect 201552 394000 201558 394012
rect 306466 394000 306472 394012
rect 306524 394000 306530 394052
rect 301498 393932 301504 393984
rect 301556 393972 301562 393984
rect 542354 393972 542360 393984
rect 301556 393944 542360 393972
rect 301556 393932 301562 393944
rect 542354 393932 542360 393944
rect 542412 393932 542418 393984
rect 304442 392640 304448 392692
rect 304500 392680 304506 392692
rect 331214 392680 331220 392692
rect 304500 392652 331220 392680
rect 304500 392640 304506 392652
rect 331214 392640 331220 392652
rect 331272 392640 331278 392692
rect 155218 392572 155224 392624
rect 155276 392612 155282 392624
rect 307754 392612 307760 392624
rect 155276 392584 307760 392612
rect 155276 392572 155282 392584
rect 307754 392572 307760 392584
rect 307812 392572 307818 392624
rect 15838 391212 15844 391264
rect 15896 391252 15902 391264
rect 255314 391252 255320 391264
rect 15896 391224 255320 391252
rect 15896 391212 15902 391224
rect 255314 391212 255320 391224
rect 255372 391212 255378 391264
rect 302878 391212 302884 391264
rect 302936 391252 302942 391264
rect 396718 391252 396724 391264
rect 302936 391224 396724 391252
rect 302936 391212 302942 391224
rect 396718 391212 396724 391224
rect 396776 391212 396782 391264
rect 255314 390532 255320 390584
rect 255372 390572 255378 390584
rect 314930 390572 314936 390584
rect 255372 390544 314936 390572
rect 255372 390532 255378 390544
rect 314930 390532 314936 390544
rect 314988 390532 314994 390584
rect 303246 389784 303252 389836
rect 303304 389824 303310 389836
rect 462314 389824 462320 389836
rect 303304 389796 462320 389824
rect 303304 389784 303310 389796
rect 462314 389784 462320 389796
rect 462372 389784 462378 389836
rect 298922 388492 298928 388544
rect 298980 388532 298986 388544
rect 323578 388532 323584 388544
rect 298980 388504 323584 388532
rect 298980 388492 298986 388504
rect 323578 388492 323584 388504
rect 323636 388492 323642 388544
rect 10318 388424 10324 388476
rect 10376 388464 10382 388476
rect 309226 388464 309232 388476
rect 10376 388436 309232 388464
rect 10376 388424 10382 388436
rect 309226 388424 309232 388436
rect 309284 388424 309290 388476
rect 296070 387132 296076 387184
rect 296128 387172 296134 387184
rect 322198 387172 322204 387184
rect 296128 387144 322204 387172
rect 296128 387132 296134 387144
rect 322198 387132 322204 387144
rect 322256 387132 322262 387184
rect 136634 387064 136640 387116
rect 136692 387104 136698 387116
rect 307846 387104 307852 387116
rect 136692 387076 307852 387104
rect 136692 387064 136698 387076
rect 307846 387064 307852 387076
rect 307904 387064 307910 387116
rect 296714 385636 296720 385688
rect 296772 385676 296778 385688
rect 324958 385676 324964 385688
rect 296772 385648 324964 385676
rect 296772 385636 296778 385648
rect 324958 385636 324964 385648
rect 325016 385636 325022 385688
rect 151078 384344 151084 384396
rect 151136 384384 151142 384396
rect 316126 384384 316132 384396
rect 151136 384356 316132 384384
rect 151136 384344 151142 384356
rect 316126 384344 316132 384356
rect 316184 384344 316190 384396
rect 301038 384276 301044 384328
rect 301096 384316 301102 384328
rect 526438 384316 526444 384328
rect 301096 384288 526444 384316
rect 301096 384276 301102 384288
rect 526438 384276 526444 384288
rect 526496 384276 526502 384328
rect 305546 383092 305552 383104
rect 267706 383064 305552 383092
rect 245654 382984 245660 383036
rect 245712 383024 245718 383036
rect 266354 383024 266360 383036
rect 245712 382996 266360 383024
rect 245712 382984 245718 382996
rect 266354 382984 266360 382996
rect 266412 383024 266418 383036
rect 267706 383024 267734 383064
rect 305546 383052 305552 383064
rect 305604 383052 305610 383104
rect 266412 382996 267734 383024
rect 266412 382984 266418 382996
rect 303338 382984 303344 383036
rect 303396 383024 303402 383036
rect 429194 383024 429200 383036
rect 303396 382996 429200 383024
rect 303396 382984 303402 382996
rect 429194 382984 429200 382996
rect 429252 382984 429258 383036
rect 71774 382916 71780 382968
rect 71832 382956 71838 382968
rect 307938 382956 307944 382968
rect 71832 382928 307944 382956
rect 71832 382916 71838 382928
rect 307938 382916 307944 382928
rect 307996 382916 308002 382968
rect 301774 381488 301780 381540
rect 301832 381528 301838 381540
rect 494054 381528 494060 381540
rect 301832 381500 494060 381528
rect 301832 381488 301838 381500
rect 494054 381488 494060 381500
rect 494112 381488 494118 381540
rect 291838 380196 291844 380248
rect 291896 380236 291902 380248
rect 312078 380236 312084 380248
rect 291896 380208 312084 380236
rect 291896 380196 291902 380208
rect 312078 380196 312084 380208
rect 312136 380196 312142 380248
rect 299750 380128 299756 380180
rect 299808 380168 299814 380180
rect 330478 380168 330484 380180
rect 299808 380140 330484 380168
rect 299808 380128 299814 380140
rect 330478 380128 330484 380140
rect 330536 380128 330542 380180
rect 292574 378156 292580 378208
rect 292632 378196 292638 378208
rect 580166 378196 580172 378208
rect 292632 378168 580172 378196
rect 292632 378156 292638 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 297082 377476 297088 377528
rect 297140 377516 297146 377528
rect 320818 377516 320824 377528
rect 297140 377488 320824 377516
rect 297140 377476 297146 377488
rect 320818 377476 320824 377488
rect 320876 377476 320882 377528
rect 298922 377408 298928 377460
rect 298980 377448 298986 377460
rect 363598 377448 363604 377460
rect 298980 377420 363604 377448
rect 298980 377408 298986 377420
rect 363598 377408 363604 377420
rect 363656 377408 363662 377460
rect 262122 376728 262128 376780
rect 262180 376768 262186 376780
rect 322382 376768 322388 376780
rect 262180 376740 322388 376768
rect 262180 376728 262186 376740
rect 322382 376728 322388 376740
rect 322440 376728 322446 376780
rect 296622 376116 296628 376168
rect 296680 376156 296686 376168
rect 318058 376156 318064 376168
rect 296680 376128 318064 376156
rect 296680 376116 296686 376128
rect 318058 376116 318064 376128
rect 318116 376116 318122 376168
rect 303154 376048 303160 376100
rect 303212 376088 303218 376100
rect 558914 376088 558920 376100
rect 303212 376060 558920 376088
rect 303212 376048 303218 376060
rect 558914 376048 558920 376060
rect 558972 376048 558978 376100
rect 3418 375980 3424 376032
rect 3476 376020 3482 376032
rect 312814 376020 312820 376032
rect 3476 375992 312820 376020
rect 3476 375980 3482 375992
rect 312814 375980 312820 375992
rect 312872 375980 312878 376032
rect 275094 375844 275100 375896
rect 275152 375884 275158 375896
rect 306374 375884 306380 375896
rect 275152 375856 306380 375884
rect 275152 375844 275158 375856
rect 306374 375844 306380 375856
rect 306432 375844 306438 375896
rect 236638 375776 236644 375828
rect 236696 375816 236702 375828
rect 294690 375816 294696 375828
rect 236696 375788 294696 375816
rect 236696 375776 236702 375788
rect 294690 375776 294696 375788
rect 294748 375816 294754 375828
rect 294874 375816 294880 375828
rect 294748 375788 294880 375816
rect 294748 375776 294754 375788
rect 294874 375776 294880 375788
rect 294932 375776 294938 375828
rect 249794 375708 249800 375760
rect 249852 375748 249858 375760
rect 309134 375748 309140 375760
rect 249852 375720 309140 375748
rect 249852 375708 249858 375720
rect 309134 375708 309140 375720
rect 309192 375708 309198 375760
rect 239398 375640 239404 375692
rect 239456 375680 239462 375692
rect 298830 375680 298836 375692
rect 239456 375652 298836 375680
rect 239456 375640 239462 375652
rect 298830 375640 298836 375652
rect 298888 375640 298894 375692
rect 244274 375572 244280 375624
rect 244332 375612 244338 375624
rect 304258 375612 304264 375624
rect 244332 375584 304264 375612
rect 244332 375572 244338 375584
rect 304258 375572 304264 375584
rect 304316 375612 304322 375624
rect 304718 375612 304724 375624
rect 304316 375584 304724 375612
rect 304316 375572 304322 375584
rect 304718 375572 304724 375584
rect 304776 375572 304782 375624
rect 238754 375504 238760 375556
rect 238812 375544 238818 375556
rect 298738 375544 298744 375556
rect 238812 375516 298744 375544
rect 238812 375504 238818 375516
rect 298738 375504 298744 375516
rect 298796 375504 298802 375556
rect 240134 375436 240140 375488
rect 240192 375476 240198 375488
rect 300302 375476 300308 375488
rect 240192 375448 300308 375476
rect 240192 375436 240198 375448
rect 300302 375436 300308 375448
rect 300360 375436 300366 375488
rect 235994 375368 236000 375420
rect 236052 375408 236058 375420
rect 297358 375408 297364 375420
rect 236052 375380 297364 375408
rect 236052 375368 236058 375380
rect 297358 375368 297364 375380
rect 297416 375368 297422 375420
rect 298738 375368 298744 375420
rect 298796 375408 298802 375420
rect 299382 375408 299388 375420
rect 298796 375380 299388 375408
rect 298796 375368 298802 375380
rect 299382 375368 299388 375380
rect 299440 375368 299446 375420
rect 306374 375368 306380 375420
rect 306432 375408 306438 375420
rect 306926 375408 306932 375420
rect 306432 375380 306932 375408
rect 306432 375368 306438 375380
rect 306926 375368 306932 375380
rect 306984 375368 306990 375420
rect 309134 375368 309140 375420
rect 309192 375408 309198 375420
rect 310238 375408 310244 375420
rect 309192 375380 310244 375408
rect 309192 375368 309198 375380
rect 310238 375368 310244 375380
rect 310296 375368 310302 375420
rect 262490 374892 262496 374944
rect 262548 374932 262554 374944
rect 323118 374932 323124 374944
rect 262548 374904 323124 374932
rect 262548 374892 262554 374904
rect 323118 374892 323124 374904
rect 323176 374892 323182 374944
rect 278590 374824 278596 374876
rect 278648 374864 278654 374876
rect 296070 374864 296076 374876
rect 278648 374836 296076 374864
rect 278648 374824 278654 374836
rect 296070 374824 296076 374836
rect 296128 374824 296134 374876
rect 297818 374824 297824 374876
rect 297876 374864 297882 374876
rect 319438 374864 319444 374876
rect 297876 374836 319444 374864
rect 297876 374824 297882 374836
rect 319438 374824 319444 374836
rect 319496 374824 319502 374876
rect 277946 374756 277952 374808
rect 278004 374796 278010 374808
rect 304534 374796 304540 374808
rect 278004 374768 304540 374796
rect 278004 374756 278010 374768
rect 304534 374756 304540 374768
rect 304592 374756 304598 374808
rect 275738 374688 275744 374740
rect 275796 374728 275802 374740
rect 304350 374728 304356 374740
rect 275796 374700 304356 374728
rect 275796 374688 275802 374700
rect 304350 374688 304356 374700
rect 304408 374688 304414 374740
rect 278498 374620 278504 374672
rect 278556 374660 278562 374672
rect 295886 374660 295892 374672
rect 278556 374632 295892 374660
rect 278556 374620 278562 374632
rect 295886 374620 295892 374632
rect 295944 374620 295950 374672
rect 580258 374660 580264 374672
rect 299446 374632 580264 374660
rect 253198 374552 253204 374604
rect 253256 374592 253262 374604
rect 294782 374592 294788 374604
rect 253256 374564 294788 374592
rect 253256 374552 253262 374564
rect 294782 374552 294788 374564
rect 294840 374552 294846 374604
rect 295518 374552 295524 374604
rect 295576 374592 295582 374604
rect 299446 374592 299474 374632
rect 580258 374620 580264 374632
rect 580316 374620 580322 374672
rect 295576 374564 299474 374592
rect 295576 374552 295582 374564
rect 275186 374484 275192 374536
rect 275244 374524 275250 374536
rect 319070 374524 319076 374536
rect 275244 374496 319076 374524
rect 275244 374484 275250 374496
rect 319070 374484 319076 374496
rect 319128 374484 319134 374536
rect 255958 374416 255964 374468
rect 256016 374456 256022 374468
rect 299750 374456 299756 374468
rect 256016 374428 299756 374456
rect 256016 374416 256022 374428
rect 299750 374416 299756 374428
rect 299808 374416 299814 374468
rect 257338 374348 257344 374400
rect 257396 374388 257402 374400
rect 300762 374388 300768 374400
rect 257396 374360 300768 374388
rect 257396 374348 257402 374360
rect 300762 374348 300768 374360
rect 300820 374388 300826 374400
rect 303154 374388 303160 374400
rect 300820 374360 303160 374388
rect 300820 374348 300826 374360
rect 303154 374348 303160 374360
rect 303212 374348 303218 374400
rect 313274 374348 313280 374400
rect 313332 374388 313338 374400
rect 313458 374388 313464 374400
rect 313332 374360 313464 374388
rect 313332 374348 313338 374360
rect 313458 374348 313464 374360
rect 313516 374348 313522 374400
rect 259638 374280 259644 374332
rect 259696 374320 259702 374332
rect 319806 374320 319812 374332
rect 259696 374292 319812 374320
rect 259696 374280 259702 374292
rect 319806 374280 319812 374292
rect 319864 374280 319870 374332
rect 264882 374212 264888 374264
rect 264940 374252 264946 374264
rect 325326 374252 325332 374264
rect 264940 374224 325332 374252
rect 264940 374212 264946 374224
rect 325326 374212 325332 374224
rect 325384 374212 325390 374264
rect 234706 374144 234712 374196
rect 234764 374184 234770 374196
rect 294598 374184 294604 374196
rect 234764 374156 294604 374184
rect 234764 374144 234770 374156
rect 294598 374144 294604 374156
rect 294656 374144 294662 374196
rect 260098 374076 260104 374128
rect 260156 374116 260162 374128
rect 320174 374116 320180 374128
rect 260156 374088 320180 374116
rect 260156 374076 260162 374088
rect 320174 374076 320180 374088
rect 320232 374076 320238 374128
rect 281074 374008 281080 374060
rect 281132 374048 281138 374060
rect 297818 374048 297824 374060
rect 281132 374020 297824 374048
rect 281132 374008 281138 374020
rect 297818 374008 297824 374020
rect 297876 374008 297882 374060
rect 295794 373600 295800 373652
rect 295852 373640 295858 373652
rect 296070 373640 296076 373652
rect 295852 373612 296076 373640
rect 295852 373600 295858 373612
rect 296070 373600 296076 373612
rect 296128 373600 296134 373652
rect 294322 373532 294328 373584
rect 294380 373572 294386 373584
rect 294782 373572 294788 373584
rect 294380 373544 294788 373572
rect 294380 373532 294386 373544
rect 294782 373532 294788 373544
rect 294840 373532 294846 373584
rect 230474 373328 230480 373380
rect 230532 373368 230538 373380
rect 291562 373368 291568 373380
rect 230532 373340 291568 373368
rect 230532 373328 230538 373340
rect 291562 373328 291568 373340
rect 291620 373328 291626 373380
rect 304442 373328 304448 373380
rect 304500 373368 304506 373380
rect 364334 373368 364340 373380
rect 304500 373340 364340 373368
rect 304500 373328 304506 373340
rect 364334 373328 364340 373340
rect 364392 373328 364398 373380
rect 234614 373260 234620 373312
rect 234672 373300 234678 373312
rect 248414 373300 248420 373312
rect 234672 373272 248420 373300
rect 234672 373260 234678 373272
rect 248414 373260 248420 373272
rect 248472 373260 248478 373312
rect 262398 373192 262404 373244
rect 262456 373232 262462 373244
rect 313734 373232 313740 373244
rect 262456 373204 313740 373232
rect 262456 373192 262462 373204
rect 313734 373192 313740 373204
rect 313792 373192 313798 373244
rect 258810 373124 258816 373176
rect 258868 373164 258874 373176
rect 317322 373164 317328 373176
rect 258868 373136 317328 373164
rect 258868 373124 258874 373136
rect 317322 373124 317328 373136
rect 317380 373124 317386 373176
rect 257430 373056 257436 373108
rect 257488 373096 257494 373108
rect 317230 373096 317236 373108
rect 257488 373068 317236 373096
rect 257488 373056 257494 373068
rect 317230 373056 317236 373068
rect 317288 373056 317294 373108
rect 229094 372988 229100 373040
rect 229152 373028 229158 373040
rect 288986 373028 288992 373040
rect 229152 373000 288992 373028
rect 229152 372988 229158 373000
rect 288986 372988 288992 373000
rect 289044 373028 289050 373040
rect 577590 373028 577596 373040
rect 289044 373000 577596 373028
rect 289044 372988 289050 373000
rect 577590 372988 577596 373000
rect 577648 372988 577654 373040
rect 258718 372920 258724 372972
rect 258776 372960 258782 372972
rect 318794 372960 318800 372972
rect 258776 372932 318800 372960
rect 258776 372920 258782 372932
rect 318794 372920 318800 372932
rect 318852 372920 318858 372972
rect 262306 372852 262312 372904
rect 262364 372892 262370 372904
rect 322934 372892 322940 372904
rect 262364 372864 322940 372892
rect 262364 372852 262370 372864
rect 322934 372852 322940 372864
rect 322992 372852 322998 372904
rect 259546 372784 259552 372836
rect 259604 372824 259610 372836
rect 320542 372824 320548 372836
rect 259604 372796 320548 372824
rect 259604 372784 259610 372796
rect 320542 372784 320548 372796
rect 320600 372784 320606 372836
rect 261018 372716 261024 372768
rect 261076 372756 261082 372768
rect 321646 372756 321652 372768
rect 261076 372728 321652 372756
rect 261076 372716 261082 372728
rect 321646 372716 321652 372728
rect 321704 372716 321710 372768
rect 275922 372648 275928 372700
rect 275980 372688 275986 372700
rect 323486 372688 323492 372700
rect 275980 372660 323492 372688
rect 275980 372648 275986 372660
rect 323486 372648 323492 372660
rect 323544 372648 323550 372700
rect 3418 372580 3424 372632
rect 3476 372620 3482 372632
rect 256694 372620 256700 372632
rect 3476 372592 256700 372620
rect 3476 372580 3482 372592
rect 256694 372580 256700 372592
rect 256752 372620 256758 372632
rect 257430 372620 257436 372632
rect 256752 372592 257436 372620
rect 256752 372580 256758 372592
rect 257430 372580 257436 372592
rect 257488 372580 257494 372632
rect 281166 372580 281172 372632
rect 281224 372620 281230 372632
rect 295518 372620 295524 372632
rect 281224 372592 295524 372620
rect 281224 372580 281230 372592
rect 295518 372580 295524 372592
rect 295576 372580 295582 372632
rect 307754 372512 307760 372564
rect 307812 372552 307818 372564
rect 308030 372552 308036 372564
rect 307812 372524 308036 372552
rect 307812 372512 307818 372524
rect 308030 372512 308036 372524
rect 308088 372512 308094 372564
rect 245746 372172 245752 372224
rect 245804 372212 245810 372224
rect 304994 372212 305000 372224
rect 245804 372184 305000 372212
rect 245804 372172 245810 372184
rect 304994 372172 305000 372184
rect 305052 372212 305058 372224
rect 305822 372212 305828 372224
rect 305052 372184 305828 372212
rect 305052 372172 305058 372184
rect 305822 372172 305828 372184
rect 305880 372172 305886 372224
rect 245010 372104 245016 372156
rect 245068 372144 245074 372156
rect 292206 372144 292212 372156
rect 245068 372116 292212 372144
rect 245068 372104 245074 372116
rect 292206 372104 292212 372116
rect 292264 372144 292270 372156
rect 363598 372144 363604 372156
rect 292264 372116 363604 372144
rect 292264 372104 292270 372116
rect 363598 372104 363604 372116
rect 363656 372104 363662 372156
rect 243538 372036 243544 372088
rect 243596 372076 243602 372088
rect 288250 372076 288256 372088
rect 243596 372048 288256 372076
rect 243596 372036 243602 372048
rect 288250 372036 288256 372048
rect 288308 372036 288314 372088
rect 289262 372036 289268 372088
rect 289320 372076 289326 372088
rect 577498 372076 577504 372088
rect 289320 372048 577504 372076
rect 289320 372036 289326 372048
rect 577498 372036 577504 372048
rect 577556 372036 577562 372088
rect 279510 371968 279516 372020
rect 279568 372008 279574 372020
rect 290550 372008 290556 372020
rect 279568 371980 290556 372008
rect 279568 371968 279574 371980
rect 290550 371968 290556 371980
rect 290608 371968 290614 372020
rect 313734 371968 313740 372020
rect 313792 372008 313798 372020
rect 322014 372008 322020 372020
rect 313792 371980 322020 372008
rect 313792 371968 313798 371980
rect 322014 371968 322020 371980
rect 322072 371968 322078 372020
rect 280798 371900 280804 371952
rect 280856 371940 280862 371952
rect 314746 371940 314752 371952
rect 280856 371912 314752 371940
rect 280856 371900 280862 371912
rect 314746 371900 314752 371912
rect 314804 371940 314810 371952
rect 315758 371940 315764 371952
rect 314804 371912 315764 371940
rect 314804 371900 314810 371912
rect 315758 371900 315764 371912
rect 315816 371900 315822 371952
rect 280890 371832 280896 371884
rect 280948 371872 280954 371884
rect 316034 371872 316040 371884
rect 280948 371844 316040 371872
rect 280948 371832 280954 371844
rect 316034 371832 316040 371844
rect 316092 371872 316098 371884
rect 316862 371872 316868 371884
rect 316092 371844 316868 371872
rect 316092 371832 316098 371844
rect 316862 371832 316868 371844
rect 316920 371832 316926 371884
rect 280430 371764 280436 371816
rect 280488 371804 280494 371816
rect 317966 371804 317972 371816
rect 280488 371776 317972 371804
rect 280488 371764 280494 371776
rect 317966 371764 317972 371776
rect 318024 371764 318030 371816
rect 279418 371696 279424 371748
rect 279476 371736 279482 371748
rect 321278 371736 321284 371748
rect 279476 371708 321284 371736
rect 279476 371696 279482 371708
rect 321278 371696 321284 371708
rect 321336 371696 321342 371748
rect 280982 371628 280988 371680
rect 281040 371668 281046 371680
rect 313458 371668 313464 371680
rect 281040 371640 313464 371668
rect 281040 371628 281046 371640
rect 313458 371628 313464 371640
rect 313516 371628 313522 371680
rect 280246 371560 280252 371612
rect 280304 371600 280310 371612
rect 324590 371600 324596 371612
rect 280304 371572 324596 371600
rect 280304 371560 280310 371572
rect 324590 371560 324596 371572
rect 324648 371560 324654 371612
rect 247678 371492 247684 371544
rect 247736 371532 247742 371544
rect 293678 371532 293684 371544
rect 247736 371504 293684 371532
rect 247736 371492 247742 371504
rect 293678 371492 293684 371504
rect 293736 371492 293742 371544
rect 293954 371492 293960 371544
rect 294012 371532 294018 371544
rect 335998 371532 336004 371544
rect 294012 371504 336004 371532
rect 294012 371492 294018 371504
rect 335998 371492 336004 371504
rect 336056 371492 336062 371544
rect 250438 371424 250444 371476
rect 250496 371464 250502 371476
rect 308030 371464 308036 371476
rect 250496 371436 308036 371464
rect 250496 371424 250502 371436
rect 308030 371424 308036 371436
rect 308088 371424 308094 371476
rect 308858 371424 308864 371476
rect 308916 371464 308922 371476
rect 316126 371464 316132 371476
rect 308916 371436 316132 371464
rect 308916 371424 308922 371436
rect 316126 371424 316132 371436
rect 316184 371424 316190 371476
rect 317322 371424 317328 371476
rect 317380 371464 317386 371476
rect 318334 371464 318340 371476
rect 317380 371436 318340 371464
rect 317380 371424 317386 371436
rect 318334 371424 318340 371436
rect 318392 371424 318398 371476
rect 290550 371356 290556 371408
rect 290608 371396 290614 371408
rect 299474 371396 299480 371408
rect 290608 371368 299480 371396
rect 290608 371356 290614 371368
rect 299474 371356 299480 371368
rect 299532 371356 299538 371408
rect 314838 371396 314844 371408
rect 302206 371368 314844 371396
rect 281994 371288 282000 371340
rect 282052 371328 282058 371340
rect 291838 371328 291844 371340
rect 282052 371300 291844 371328
rect 282052 371288 282058 371300
rect 291838 371288 291844 371300
rect 291896 371288 291902 371340
rect 299290 371288 299296 371340
rect 299348 371328 299354 371340
rect 302206 371328 302234 371368
rect 314838 371356 314844 371368
rect 314896 371356 314902 371408
rect 299348 371300 302234 371328
rect 299348 371288 299354 371300
rect 242158 371220 242164 371272
rect 242216 371260 242222 371272
rect 289262 371260 289268 371272
rect 242216 371232 289268 371260
rect 242216 371220 242222 371232
rect 289262 371220 289268 371232
rect 289320 371220 289326 371272
rect 314562 371220 314568 371272
rect 314620 371260 314626 371272
rect 319438 371260 319444 371272
rect 314620 371232 319444 371260
rect 314620 371220 314626 371232
rect 319438 371220 319444 371232
rect 319496 371220 319502 371272
rect 319530 371220 319536 371272
rect 319588 371260 319594 371272
rect 323854 371260 323860 371272
rect 319588 371232 323860 371260
rect 319588 371220 319594 371232
rect 323854 371220 323860 371232
rect 323912 371220 323918 371272
rect 241514 370744 241520 370796
rect 241572 370784 241578 370796
rect 302234 370784 302240 370796
rect 241572 370756 302240 370784
rect 241572 370744 241578 370756
rect 302234 370744 302240 370756
rect 302292 370784 302298 370796
rect 303246 370784 303252 370796
rect 302292 370756 303252 370784
rect 302292 370744 302298 370756
rect 303246 370744 303252 370756
rect 303304 370744 303310 370796
rect 260190 370676 260196 370728
rect 260248 370716 260254 370728
rect 314562 370716 314568 370728
rect 260248 370688 314568 370716
rect 260248 370676 260254 370688
rect 314562 370676 314568 370688
rect 314620 370676 314626 370728
rect 229186 370608 229192 370660
rect 229244 370648 229250 370660
rect 289998 370648 290004 370660
rect 229244 370620 290004 370648
rect 229244 370608 229250 370620
rect 289998 370608 290004 370620
rect 290056 370608 290062 370660
rect 293678 370608 293684 370660
rect 293736 370648 293742 370660
rect 293736 370620 297220 370648
rect 293736 370608 293742 370620
rect 236086 370540 236092 370592
rect 236144 370580 236150 370592
rect 297082 370580 297088 370592
rect 236144 370552 297088 370580
rect 236144 370540 236150 370552
rect 297082 370540 297088 370552
rect 297140 370540 297146 370592
rect 231946 370472 231952 370524
rect 232004 370512 232010 370524
rect 292942 370512 292948 370524
rect 232004 370484 292948 370512
rect 232004 370472 232010 370484
rect 292942 370472 292948 370484
rect 293000 370512 293006 370524
rect 293770 370512 293776 370524
rect 293000 370484 293776 370512
rect 293000 370472 293006 370484
rect 293770 370472 293776 370484
rect 293828 370472 293834 370524
rect 297192 370512 297220 370620
rect 302326 370608 302332 370660
rect 302384 370648 302390 370660
rect 580350 370648 580356 370660
rect 302384 370620 580356 370648
rect 302384 370608 302390 370620
rect 580350 370608 580356 370620
rect 580408 370608 580414 370660
rect 299474 370540 299480 370592
rect 299532 370580 299538 370592
rect 580534 370580 580540 370592
rect 299532 370552 580540 370580
rect 299532 370540 299538 370552
rect 580534 370540 580540 370552
rect 580592 370540 580598 370592
rect 580166 370512 580172 370524
rect 297192 370484 580172 370512
rect 580166 370472 580172 370484
rect 580224 370472 580230 370524
rect 244918 370404 244924 370456
rect 244976 370444 244982 370456
rect 296622 370444 296628 370456
rect 244976 370416 296628 370444
rect 244976 370404 244982 370416
rect 296622 370404 296628 370416
rect 296680 370404 296686 370456
rect 231854 370336 231860 370388
rect 231912 370376 231918 370388
rect 292666 370376 292672 370388
rect 231912 370348 292672 370376
rect 231912 370336 231918 370348
rect 292666 370336 292672 370348
rect 292724 370376 292730 370388
rect 329098 370376 329104 370388
rect 292724 370348 329104 370376
rect 292724 370336 292730 370348
rect 329098 370336 329104 370348
rect 329156 370336 329162 370388
rect 242894 370268 242900 370320
rect 242952 370308 242958 370320
rect 302878 370308 302884 370320
rect 242952 370280 302884 370308
rect 242952 370268 242958 370280
rect 302878 370268 302884 370280
rect 302936 370268 302942 370320
rect 245838 370200 245844 370252
rect 245896 370240 245902 370252
rect 306558 370240 306564 370252
rect 245896 370212 306564 370240
rect 245896 370200 245902 370212
rect 306558 370200 306564 370212
rect 306616 370200 306622 370252
rect 247034 370132 247040 370184
rect 247092 370172 247098 370184
rect 307662 370172 307668 370184
rect 247092 370144 307668 370172
rect 247092 370132 247098 370144
rect 307662 370132 307668 370144
rect 307720 370132 307726 370184
rect 277854 370064 277860 370116
rect 277912 370104 277918 370116
rect 293172 370104 293178 370116
rect 277912 370076 293178 370104
rect 277912 370064 277918 370076
rect 293172 370064 293178 370076
rect 293230 370104 293236 370116
rect 329190 370104 329196 370116
rect 293230 370076 329196 370104
rect 293230 370064 293236 370076
rect 329190 370064 329196 370076
rect 329248 370064 329254 370116
rect 282270 369996 282276 370048
rect 282328 370036 282334 370048
rect 317598 370036 317604 370048
rect 282328 370008 317604 370036
rect 282328 369996 282334 370008
rect 317598 369996 317604 370008
rect 317656 369996 317662 370048
rect 281350 369928 281356 369980
rect 281408 369968 281414 369980
rect 281408 369940 290412 369968
rect 281408 369928 281414 369940
rect 281442 369860 281448 369912
rect 281500 369900 281506 369912
rect 288526 369900 288532 369912
rect 281500 369872 288532 369900
rect 281500 369860 281506 369872
rect 288526 369860 288532 369872
rect 288584 369860 288590 369912
rect 290384 369900 290412 369940
rect 291562 369928 291568 369980
rect 291620 369968 291626 369980
rect 330478 369968 330484 369980
rect 291620 369940 330484 369968
rect 291620 369928 291626 369940
rect 330478 369928 330484 369940
rect 330536 369928 330542 369980
rect 290734 369900 290740 369912
rect 290384 369872 290740 369900
rect 290734 369860 290740 369872
rect 290792 369860 290798 369912
rect 345658 369900 345664 369912
rect 299446 369872 345664 369900
rect 290458 369656 290464 369708
rect 290516 369696 290522 369708
rect 299446 369696 299474 369872
rect 345658 369860 345664 369872
rect 345716 369860 345722 369912
rect 290516 369668 299474 369696
rect 290516 369656 290522 369668
rect 291930 369588 291936 369640
rect 291988 369628 291994 369640
rect 292206 369628 292212 369640
rect 291988 369600 292212 369628
rect 291988 369588 291994 369600
rect 292206 369588 292212 369600
rect 292264 369588 292270 369640
rect 308858 369492 308864 369504
rect 290108 369464 308864 369492
rect 282362 369384 282368 369436
rect 282420 369424 282426 369436
rect 284110 369424 284116 369436
rect 282420 369396 284116 369424
rect 282420 369384 282426 369396
rect 284110 369384 284116 369396
rect 284168 369384 284174 369436
rect 289998 369424 290004 369436
rect 286428 369396 290004 369424
rect 282178 369316 282184 369368
rect 282236 369356 282242 369368
rect 286428 369356 286456 369396
rect 289998 369384 290004 369396
rect 290056 369384 290062 369436
rect 290108 369356 290136 369464
rect 308858 369452 308864 369464
rect 308916 369452 308922 369504
rect 292298 369424 292304 369436
rect 282236 369328 286456 369356
rect 289096 369328 290136 369356
rect 291166 369396 292304 369424
rect 282236 369316 282242 369328
rect 255406 369248 255412 369300
rect 255464 369288 255470 369300
rect 289096 369288 289124 369328
rect 255464 369260 289124 369288
rect 255464 369248 255470 369260
rect 245930 369180 245936 369232
rect 245988 369220 245994 369232
rect 248414 369220 248420 369232
rect 245988 369192 248420 369220
rect 245988 369180 245994 369192
rect 248414 369180 248420 369192
rect 248472 369220 248478 369232
rect 282454 369220 282460 369232
rect 248472 369192 282460 369220
rect 248472 369180 248478 369192
rect 282454 369180 282460 369192
rect 282512 369180 282518 369232
rect 229278 369112 229284 369164
rect 229336 369152 229342 369164
rect 282178 369152 282184 369164
rect 229336 369124 282184 369152
rect 229336 369112 229342 369124
rect 282178 369112 282184 369124
rect 282236 369112 282242 369164
rect 291166 369016 291194 369396
rect 292298 369384 292304 369396
rect 292356 369424 292362 369436
rect 293310 369424 293316 369436
rect 292356 369396 293316 369424
rect 292356 369384 292362 369396
rect 293310 369384 293316 369396
rect 293368 369384 293374 369436
rect 306282 369424 306288 369436
rect 302206 369396 306288 369424
rect 298066 369260 299474 369288
rect 298066 369016 298094 369260
rect 299446 369152 299474 369260
rect 302206 369152 302234 369396
rect 306282 369384 306288 369396
rect 306340 369384 306346 369436
rect 326246 369384 326252 369436
rect 326304 369424 326310 369436
rect 329006 369424 329012 369436
rect 326304 369396 329012 369424
rect 326304 369384 326310 369396
rect 329006 369384 329012 369396
rect 329064 369384 329070 369436
rect 299446 369124 302234 369152
rect 277366 368988 291194 369016
rect 293926 368988 298094 369016
rect 233234 368500 233240 368552
rect 233292 368540 233298 368552
rect 277366 368540 277394 368988
rect 282454 368772 282460 368824
rect 282512 368812 282518 368824
rect 293926 368812 293954 368988
rect 282512 368784 293954 368812
rect 282512 368772 282518 368784
rect 233292 368512 277394 368540
rect 233292 368500 233298 368512
rect 264238 366324 264244 366376
rect 264296 366364 264302 366376
rect 280246 366364 280252 366376
rect 264296 366336 280252 366364
rect 264296 366324 264302 366336
rect 280246 366324 280252 366336
rect 280304 366324 280310 366376
rect 258350 364352 258356 364404
rect 258408 364392 258414 364404
rect 280430 364392 280436 364404
rect 258408 364364 280436 364392
rect 258408 364352 258414 364364
rect 280430 364352 280436 364364
rect 280488 364352 280494 364404
rect 223758 360204 223764 360256
rect 223816 360244 223822 360256
rect 280706 360244 280712 360256
rect 223816 360216 280712 360244
rect 223816 360204 223822 360216
rect 280706 360204 280712 360216
rect 280764 360204 280770 360256
rect 226334 358776 226340 358828
rect 226392 358816 226398 358828
rect 280062 358816 280068 358828
rect 226392 358788 280068 358816
rect 226392 358776 226398 358788
rect 280062 358776 280068 358788
rect 280120 358816 280126 358828
rect 280706 358816 280712 358828
rect 280120 358788 280712 358816
rect 280120 358776 280126 358788
rect 280706 358776 280712 358788
rect 280764 358776 280770 358828
rect 3418 358028 3424 358080
rect 3476 358068 3482 358080
rect 258350 358068 258356 358080
rect 3476 358040 258356 358068
rect 3476 358028 3482 358040
rect 258350 358028 258356 358040
rect 258408 358028 258414 358080
rect 252554 356668 252560 356720
rect 252612 356708 252618 356720
rect 280982 356708 280988 356720
rect 252612 356680 280988 356708
rect 252612 356668 252618 356680
rect 280982 356668 280988 356680
rect 281040 356668 281046 356720
rect 329190 353200 329196 353252
rect 329248 353240 329254 353252
rect 579614 353240 579620 353252
rect 329248 353212 579620 353240
rect 329248 353200 329254 353212
rect 579614 353200 579620 353212
rect 579672 353200 579678 353252
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 256786 345080 256792 345092
rect 3384 345052 256792 345080
rect 3384 345040 3390 345052
rect 256786 345040 256792 345052
rect 256844 345040 256850 345092
rect 230566 327700 230572 327752
rect 230624 327740 230630 327752
rect 279510 327740 279516 327752
rect 230624 327712 279516 327740
rect 230624 327700 230630 327712
rect 279510 327700 279516 327712
rect 279568 327700 279574 327752
rect 261478 326340 261484 326392
rect 261536 326380 261542 326392
rect 279418 326380 279424 326392
rect 261536 326352 279424 326380
rect 261536 326340 261542 326352
rect 279418 326340 279424 326352
rect 279476 326340 279482 326392
rect 329098 325592 329104 325644
rect 329156 325632 329162 325644
rect 580166 325632 580172 325644
rect 329156 325604 580172 325632
rect 329156 325592 329162 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 256878 324912 256884 324964
rect 256936 324952 256942 324964
rect 280890 324952 280896 324964
rect 256936 324924 280896 324952
rect 256936 324912 256942 324924
rect 280890 324912 280896 324924
rect 280948 324912 280954 324964
rect 255498 323552 255504 323604
rect 255556 323592 255562 323604
rect 280798 323592 280804 323604
rect 255556 323564 280804 323592
rect 255556 323552 255562 323564
rect 280798 323552 280804 323564
rect 280856 323552 280862 323604
rect 225046 322192 225052 322244
rect 225104 322232 225110 322244
rect 279970 322232 279976 322244
rect 225104 322204 279976 322232
rect 225104 322192 225110 322204
rect 279970 322192 279976 322204
rect 280028 322232 280034 322244
rect 280798 322232 280804 322244
rect 280028 322204 280804 322232
rect 280028 322192 280034 322204
rect 280798 322192 280804 322204
rect 280856 322192 280862 322244
rect 314626 321048 325694 321076
rect 281902 320968 281908 321020
rect 281960 321008 281966 321020
rect 281960 320980 293954 321008
rect 281960 320968 281966 320980
rect 293926 320940 293954 320980
rect 293926 320912 296714 320940
rect 282270 320696 282276 320748
rect 282328 320736 282334 320748
rect 283696 320736 283702 320748
rect 282328 320708 283702 320736
rect 282328 320696 282334 320708
rect 283696 320696 283702 320708
rect 283754 320696 283760 320748
rect 283806 320708 293954 320736
rect 282178 320628 282184 320680
rect 282236 320668 282242 320680
rect 283806 320668 283834 320708
rect 293926 320668 293954 320708
rect 296686 320668 296714 320912
rect 302924 320668 302930 320680
rect 282236 320640 283834 320668
rect 288038 320640 288342 320668
rect 293926 320640 295334 320668
rect 296686 320640 302930 320668
rect 282236 320628 282242 320640
rect 211062 320560 211068 320612
rect 211120 320600 211126 320612
rect 285812 320600 285818 320612
rect 211120 320572 285818 320600
rect 211120 320560 211126 320572
rect 285812 320560 285818 320572
rect 285870 320560 285876 320612
rect 272610 320492 272616 320544
rect 272668 320532 272674 320544
rect 281902 320532 281908 320544
rect 272668 320504 281908 320532
rect 272668 320492 272674 320504
rect 281902 320492 281908 320504
rect 281960 320492 281966 320544
rect 288038 320532 288066 320640
rect 288314 320600 288342 320640
rect 295306 320600 295334 320640
rect 302924 320628 302930 320640
rect 302982 320628 302988 320680
rect 314626 320668 314654 321048
rect 325666 320872 325694 321048
rect 303034 320640 303614 320668
rect 303034 320600 303062 320640
rect 288314 320572 293954 320600
rect 295306 320572 303062 320600
rect 287900 320504 288066 320532
rect 293926 320532 293954 320572
rect 303586 320532 303614 320640
rect 309290 320640 314654 320668
rect 316006 320844 317184 320872
rect 325666 320844 328454 320872
rect 304966 320572 307754 320600
rect 304966 320532 304994 320572
rect 293926 320504 296714 320532
rect 303586 320504 304994 320532
rect 248506 320424 248512 320476
rect 248564 320464 248570 320476
rect 287900 320464 287928 320504
rect 248564 320436 287928 320464
rect 248564 320424 248570 320436
rect 249978 320356 249984 320408
rect 250036 320396 250042 320408
rect 282178 320396 282184 320408
rect 250036 320368 282184 320396
rect 250036 320356 250042 320368
rect 282178 320356 282184 320368
rect 282236 320356 282242 320408
rect 219158 320288 219164 320340
rect 219216 320328 219222 320340
rect 292436 320328 292442 320340
rect 219216 320300 292442 320328
rect 219216 320288 219222 320300
rect 292436 320288 292442 320300
rect 292494 320288 292500 320340
rect 296686 320328 296714 320504
rect 302206 320436 304994 320464
rect 302206 320328 302234 320436
rect 296686 320300 302234 320328
rect 275646 320220 275652 320272
rect 275704 320260 275710 320272
rect 275704 320232 295518 320260
rect 275704 320220 275710 320232
rect 219342 320152 219348 320204
rect 219400 320192 219406 320204
rect 295490 320192 295518 320232
rect 304966 320192 304994 320436
rect 307726 320260 307754 320572
rect 307726 320232 309226 320260
rect 219400 320164 295334 320192
rect 295490 320164 296346 320192
rect 304966 320164 307524 320192
rect 219400 320152 219406 320164
rect 280706 320084 280712 320136
rect 280764 320124 280770 320136
rect 280764 320096 288434 320124
rect 280764 320084 280770 320096
rect 284616 320056 284622 320068
rect 273226 320028 284622 320056
rect 224862 319676 224868 319728
rect 224920 319716 224926 319728
rect 273226 319716 273254 320028
rect 284616 320016 284622 320028
rect 284674 320016 284680 320068
rect 287008 320016 287014 320068
rect 287066 320016 287072 320068
rect 288406 320056 288434 320096
rect 295306 320056 295334 320164
rect 288406 320028 292758 320056
rect 295306 320028 295978 320056
rect 281994 319880 282000 319932
rect 282052 319920 282058 319932
rect 283328 319920 283334 319932
rect 282052 319892 283334 319920
rect 282052 319880 282058 319892
rect 283328 319880 283334 319892
rect 283386 319880 283392 319932
rect 283512 319880 283518 319932
rect 283570 319880 283576 319932
rect 283742 319880 283748 319932
rect 283800 319920 283806 319932
rect 283972 319920 283978 319932
rect 283800 319892 283978 319920
rect 283800 319880 283806 319892
rect 283972 319880 283978 319892
rect 284030 319880 284036 319932
rect 284340 319880 284346 319932
rect 284398 319880 284404 319932
rect 284800 319920 284806 319932
rect 284772 319880 284806 319920
rect 284858 319880 284864 319932
rect 284892 319880 284898 319932
rect 284950 319880 284956 319932
rect 281718 319812 281724 319864
rect 281776 319852 281782 319864
rect 282684 319852 282690 319864
rect 281776 319824 282690 319852
rect 281776 319812 281782 319824
rect 282684 319812 282690 319824
rect 282742 319812 282748 319864
rect 224920 319688 273254 319716
rect 224920 319676 224926 319688
rect 283190 319676 283196 319728
rect 283248 319716 283254 319728
rect 283530 319716 283558 319880
rect 283248 319688 283558 319716
rect 284358 319716 284386 319880
rect 284772 319796 284800 319880
rect 284754 319744 284760 319796
rect 284812 319744 284818 319796
rect 284478 319716 284484 319728
rect 284358 319688 284484 319716
rect 283248 319676 283254 319688
rect 284478 319676 284484 319688
rect 284536 319676 284542 319728
rect 284910 319716 284938 319880
rect 286364 319812 286370 319864
rect 286422 319852 286428 319864
rect 286422 319824 286548 319852
rect 286422 319812 286428 319824
rect 286520 319796 286548 319824
rect 286502 319744 286508 319796
rect 286560 319744 286566 319796
rect 285030 319716 285036 319728
rect 284910 319688 285036 319716
rect 285030 319676 285036 319688
rect 285088 319676 285094 319728
rect 285950 319676 285956 319728
rect 286008 319716 286014 319728
rect 287026 319716 287054 320016
rect 292730 319932 292758 320028
rect 293236 319960 295426 319988
rect 287468 319880 287474 319932
rect 287526 319920 287532 319932
rect 289492 319920 289498 319932
rect 287526 319880 287560 319920
rect 287532 319796 287560 319880
rect 289464 319880 289498 319920
rect 289550 319880 289556 319932
rect 290044 319920 290050 319932
rect 290016 319880 290050 319920
rect 290102 319880 290108 319932
rect 291608 319880 291614 319932
rect 291666 319880 291672 319932
rect 292712 319880 292718 319932
rect 292770 319880 292776 319932
rect 289464 319796 289492 319880
rect 290016 319796 290044 319880
rect 287514 319744 287520 319796
rect 287572 319744 287578 319796
rect 289446 319744 289452 319796
rect 289504 319744 289510 319796
rect 289998 319744 290004 319796
rect 290056 319744 290062 319796
rect 291626 319728 291654 319880
rect 286008 319688 287054 319716
rect 286008 319676 286014 319688
rect 291562 319676 291568 319728
rect 291620 319688 291654 319728
rect 291620 319676 291626 319688
rect 269758 319608 269764 319660
rect 269816 319648 269822 319660
rect 293236 319648 293264 319960
rect 293816 319920 293822 319932
rect 293788 319880 293822 319920
rect 293874 319880 293880 319932
rect 294552 319880 294558 319932
rect 294610 319880 294616 319932
rect 295196 319880 295202 319932
rect 295254 319880 295260 319932
rect 295288 319880 295294 319932
rect 295346 319880 295352 319932
rect 293788 319796 293816 319880
rect 293908 319812 293914 319864
rect 293966 319812 293972 319864
rect 294322 319812 294328 319864
rect 294380 319852 294386 319864
rect 294570 319852 294598 319880
rect 294380 319824 294598 319852
rect 294380 319812 294386 319824
rect 293770 319744 293776 319796
rect 293828 319744 293834 319796
rect 293926 319784 293954 319812
rect 293880 319756 293954 319784
rect 293880 319660 293908 319756
rect 295214 319728 295242 319880
rect 295150 319676 295156 319728
rect 295208 319688 295242 319728
rect 295208 319676 295214 319688
rect 269816 319620 293264 319648
rect 269816 319608 269822 319620
rect 293862 319608 293868 319660
rect 293920 319608 293926 319660
rect 293954 319608 293960 319660
rect 294012 319648 294018 319660
rect 295306 319648 295334 319880
rect 294012 319620 295334 319648
rect 295398 319648 295426 319960
rect 295748 319880 295754 319932
rect 295806 319880 295812 319932
rect 295518 319676 295524 319728
rect 295576 319716 295582 319728
rect 295766 319716 295794 319880
rect 295950 319852 295978 320028
rect 296318 319932 296346 320164
rect 296686 320028 303798 320056
rect 296300 319880 296306 319932
rect 296358 319880 296364 319932
rect 296576 319880 296582 319932
rect 296634 319880 296640 319932
rect 296594 319852 296622 319880
rect 295950 319824 296622 319852
rect 295576 319688 295794 319716
rect 295576 319676 295582 319688
rect 296686 319648 296714 320028
rect 295398 319620 296714 319648
rect 297054 319960 303614 319988
rect 294012 319608 294018 319620
rect 264330 319540 264336 319592
rect 264388 319580 264394 319592
rect 296530 319580 296536 319592
rect 264388 319552 296536 319580
rect 264388 319540 264394 319552
rect 296530 319540 296536 319552
rect 296588 319540 296594 319592
rect 252738 319472 252744 319524
rect 252796 319512 252802 319524
rect 297054 319512 297082 319960
rect 298324 319880 298330 319932
rect 298382 319880 298388 319932
rect 298692 319880 298698 319932
rect 298750 319880 298756 319932
rect 298784 319880 298790 319932
rect 298842 319880 298848 319932
rect 299244 319880 299250 319932
rect 299302 319880 299308 319932
rect 301268 319920 301274 319932
rect 300826 319892 301274 319920
rect 298342 319728 298370 319880
rect 298710 319784 298738 319880
rect 298278 319676 298284 319728
rect 298336 319688 298370 319728
rect 298572 319756 298738 319784
rect 298336 319676 298342 319688
rect 298572 319592 298600 319756
rect 298802 319660 298830 319880
rect 299152 319812 299158 319864
rect 299210 319812 299216 319864
rect 298738 319608 298744 319660
rect 298796 319620 298830 319660
rect 298796 319608 298802 319620
rect 298554 319540 298560 319592
rect 298612 319540 298618 319592
rect 252796 319484 297082 319512
rect 252796 319472 252802 319484
rect 237466 319404 237472 319456
rect 237524 319444 237530 319456
rect 295334 319444 295340 319456
rect 237524 319416 295340 319444
rect 237524 319404 237530 319416
rect 295334 319404 295340 319416
rect 295392 319404 295398 319456
rect 295702 319404 295708 319456
rect 295760 319444 295766 319456
rect 296070 319444 296076 319456
rect 295760 319416 296076 319444
rect 295760 319404 295766 319416
rect 296070 319404 296076 319416
rect 296128 319404 296134 319456
rect 299170 319444 299198 319812
rect 299262 319580 299290 319880
rect 300072 319812 300078 319864
rect 300130 319812 300136 319864
rect 299382 319580 299388 319592
rect 299262 319552 299388 319580
rect 299382 319540 299388 319552
rect 299440 319540 299446 319592
rect 300090 319580 300118 319812
rect 300826 319592 300854 319892
rect 301268 319880 301274 319892
rect 301326 319880 301332 319932
rect 301360 319880 301366 319932
rect 301418 319880 301424 319932
rect 301728 319880 301734 319932
rect 301786 319880 301792 319932
rect 301912 319880 301918 319932
rect 301970 319880 301976 319932
rect 303292 319880 303298 319932
rect 303350 319880 303356 319932
rect 303476 319880 303482 319932
rect 303534 319880 303540 319932
rect 301378 319796 301406 319880
rect 301452 319812 301458 319864
rect 301510 319812 301516 319864
rect 301314 319744 301320 319796
rect 301372 319756 301406 319796
rect 301372 319744 301378 319756
rect 301470 319728 301498 319812
rect 301406 319676 301412 319728
rect 301464 319688 301498 319728
rect 301464 319676 301470 319688
rect 300210 319580 300216 319592
rect 300090 319552 300216 319580
rect 300210 319540 300216 319552
rect 300268 319540 300274 319592
rect 300762 319540 300768 319592
rect 300820 319552 300854 319592
rect 300820 319540 300826 319552
rect 301590 319540 301596 319592
rect 301648 319580 301654 319592
rect 301746 319580 301774 319880
rect 301930 319728 301958 319880
rect 301866 319676 301872 319728
rect 301924 319688 301958 319728
rect 301924 319676 301930 319688
rect 302694 319676 302700 319728
rect 302752 319716 302758 319728
rect 303310 319716 303338 319880
rect 303494 319728 303522 319880
rect 303586 319852 303614 319960
rect 303770 319932 303798 320028
rect 303862 319960 305684 319988
rect 303752 319880 303758 319932
rect 303810 319880 303816 319932
rect 303862 319852 303890 319960
rect 304028 319880 304034 319932
rect 304086 319880 304092 319932
rect 304856 319920 304862 319932
rect 304644 319892 304862 319920
rect 303586 319824 303890 319852
rect 303798 319744 303804 319796
rect 303856 319784 303862 319796
rect 304046 319784 304074 319880
rect 303856 319756 304074 319784
rect 303856 319744 303862 319756
rect 302752 319688 303338 319716
rect 302752 319676 302758 319688
rect 303430 319676 303436 319728
rect 303488 319688 303522 319728
rect 303488 319676 303494 319688
rect 302418 319608 302424 319660
rect 302476 319648 302482 319660
rect 302602 319648 302608 319660
rect 302476 319620 302608 319648
rect 302476 319608 302482 319620
rect 302602 319608 302608 319620
rect 302660 319608 302666 319660
rect 301648 319552 301774 319580
rect 301648 319540 301654 319552
rect 301958 319540 301964 319592
rect 302016 319580 302022 319592
rect 302142 319580 302148 319592
rect 302016 319552 302148 319580
rect 302016 319540 302022 319552
rect 302142 319540 302148 319552
rect 302200 319540 302206 319592
rect 304258 319540 304264 319592
rect 304316 319580 304322 319592
rect 304644 319580 304672 319892
rect 304856 319880 304862 319892
rect 304914 319880 304920 319932
rect 305224 319920 305230 319932
rect 305196 319880 305230 319920
rect 305282 319880 305288 319932
rect 305316 319880 305322 319932
rect 305374 319880 305380 319932
rect 305500 319880 305506 319932
rect 305558 319880 305564 319932
rect 304764 319812 304770 319864
rect 304822 319812 304828 319864
rect 304782 319592 304810 319812
rect 305196 319796 305224 319880
rect 305334 319796 305362 319880
rect 305408 319812 305414 319864
rect 305466 319812 305472 319864
rect 305178 319744 305184 319796
rect 305236 319744 305242 319796
rect 305270 319744 305276 319796
rect 305328 319756 305362 319796
rect 305328 319744 305334 319756
rect 305426 319728 305454 319812
rect 305362 319676 305368 319728
rect 305420 319688 305454 319728
rect 305420 319676 305426 319688
rect 305518 319648 305546 319880
rect 305518 319620 305592 319648
rect 304316 319552 304672 319580
rect 304316 319540 304322 319552
rect 304718 319540 304724 319592
rect 304776 319552 304810 319592
rect 304776 319540 304782 319552
rect 299290 319444 299296 319456
rect 299170 319416 299296 319444
rect 299290 319404 299296 319416
rect 299348 319404 299354 319456
rect 300854 319404 300860 319456
rect 300912 319444 300918 319456
rect 301038 319444 301044 319456
rect 300912 319416 301044 319444
rect 300912 319404 300918 319416
rect 301038 319404 301044 319416
rect 301096 319404 301102 319456
rect 301314 319404 301320 319456
rect 301372 319444 301378 319456
rect 301590 319444 301596 319456
rect 301372 319416 301596 319444
rect 301372 319404 301378 319416
rect 301590 319404 301596 319416
rect 301648 319404 301654 319456
rect 305362 319404 305368 319456
rect 305420 319444 305426 319456
rect 305564 319444 305592 319620
rect 305656 319512 305684 319960
rect 305960 319880 305966 319932
rect 306018 319880 306024 319932
rect 306512 319880 306518 319932
rect 306570 319880 306576 319932
rect 306696 319880 306702 319932
rect 306754 319880 306760 319932
rect 305978 319660 306006 319880
rect 306530 319660 306558 319880
rect 305914 319608 305920 319660
rect 305972 319620 306006 319660
rect 305972 319608 305978 319620
rect 306466 319608 306472 319660
rect 306524 319620 306558 319660
rect 306524 319608 306530 319620
rect 306714 319580 306742 319880
rect 307496 319592 307524 320164
rect 308490 319920 308496 319932
rect 308324 319892 308496 319920
rect 308324 319864 308352 319892
rect 308490 319880 308496 319892
rect 308548 319880 308554 319932
rect 309088 319880 309094 319932
rect 309146 319880 309152 319932
rect 308306 319812 308312 319864
rect 308364 319812 308370 319864
rect 308950 319608 308956 319660
rect 309008 319648 309014 319660
rect 309106 319648 309134 319880
rect 309198 319716 309226 320232
rect 309290 319932 309318 320640
rect 309842 320572 314654 320600
rect 309842 319932 309870 320572
rect 314626 320464 314654 320572
rect 316006 320464 316034 320844
rect 317156 320804 317184 320844
rect 327626 320804 327632 320816
rect 317156 320776 327632 320804
rect 327626 320764 327632 320776
rect 327684 320764 327690 320816
rect 328178 320668 328184 320680
rect 316972 320640 328184 320668
rect 316972 320600 317000 320640
rect 328178 320628 328184 320640
rect 328236 320628 328242 320680
rect 314626 320436 316034 320464
rect 316880 320572 317000 320600
rect 328426 320600 328454 320844
rect 338574 320600 338580 320612
rect 328426 320572 338580 320600
rect 316880 320328 316908 320572
rect 338574 320560 338580 320572
rect 338632 320560 338638 320612
rect 314626 320300 316908 320328
rect 317064 320436 326982 320464
rect 314626 320124 314654 320300
rect 317064 320192 317092 320436
rect 326954 320396 326982 320436
rect 327718 320424 327724 320476
rect 327776 320464 327782 320476
rect 336734 320464 336740 320476
rect 327776 320436 336740 320464
rect 327776 320424 327782 320436
rect 336734 320424 336740 320436
rect 336792 320424 336798 320476
rect 338298 320396 338304 320408
rect 326954 320368 338304 320396
rect 338298 320356 338304 320368
rect 338356 320356 338362 320408
rect 336826 320328 336832 320340
rect 312280 320096 314654 320124
rect 314718 320164 317092 320192
rect 317156 320300 336832 320328
rect 310946 319960 312032 319988
rect 310946 319932 310974 319960
rect 309272 319880 309278 319932
rect 309330 319880 309336 319932
rect 309364 319880 309370 319932
rect 309422 319880 309428 319932
rect 309548 319880 309554 319932
rect 309606 319880 309612 319932
rect 309824 319880 309830 319932
rect 309882 319880 309888 319932
rect 310284 319880 310290 319932
rect 310342 319880 310348 319932
rect 310928 319880 310934 319932
rect 310986 319880 310992 319932
rect 311112 319880 311118 319932
rect 311170 319880 311176 319932
rect 311480 319880 311486 319932
rect 311538 319880 311544 319932
rect 309382 319796 309410 319880
rect 309318 319744 309324 319796
rect 309376 319756 309410 319796
rect 309566 319784 309594 319880
rect 309778 319784 309784 319796
rect 309566 319756 309784 319784
rect 309376 319744 309382 319756
rect 309778 319744 309784 319756
rect 309836 319744 309842 319796
rect 310302 319728 310330 319880
rect 309686 319716 309692 319728
rect 309198 319688 309692 319716
rect 309686 319676 309692 319688
rect 309744 319676 309750 319728
rect 310238 319676 310244 319728
rect 310296 319688 310330 319728
rect 311130 319716 311158 319880
rect 311250 319716 311256 319728
rect 311130 319688 311256 319716
rect 310296 319676 310302 319688
rect 311250 319676 311256 319688
rect 311308 319676 311314 319728
rect 309008 319620 309134 319648
rect 309008 319608 309014 319620
rect 309226 319608 309232 319660
rect 309284 319648 309290 319660
rect 309870 319648 309876 319660
rect 309284 319620 309876 319648
rect 309284 319608 309290 319620
rect 309870 319608 309876 319620
rect 309928 319608 309934 319660
rect 306926 319580 306932 319592
rect 306714 319552 306932 319580
rect 306926 319540 306932 319552
rect 306984 319540 306990 319592
rect 307478 319540 307484 319592
rect 307536 319540 307542 319592
rect 310882 319512 310888 319524
rect 305656 319484 310888 319512
rect 310882 319472 310888 319484
rect 310940 319472 310946 319524
rect 311498 319512 311526 319880
rect 311848 319812 311854 319864
rect 311906 319812 311912 319864
rect 311866 319592 311894 319812
rect 312004 319784 312032 319960
rect 312280 319932 312308 320096
rect 312464 320028 314654 320056
rect 312464 319988 312492 320028
rect 312418 319960 312492 319988
rect 312280 319892 312314 319932
rect 312308 319880 312314 319892
rect 312366 319880 312372 319932
rect 312418 319852 312446 319960
rect 313044 319880 313050 319932
rect 313102 319880 313108 319932
rect 313412 319880 313418 319932
rect 313470 319880 313476 319932
rect 313780 319880 313786 319932
rect 313838 319880 313844 319932
rect 312188 319824 312446 319852
rect 312188 319784 312216 319824
rect 312584 319812 312590 319864
rect 312642 319812 312648 319864
rect 312676 319812 312682 319864
rect 312734 319812 312740 319864
rect 312768 319812 312774 319864
rect 312826 319812 312832 319864
rect 312860 319812 312866 319864
rect 312918 319852 312924 319864
rect 312918 319824 312998 319852
rect 312918 319812 312924 319824
rect 312004 319756 312216 319784
rect 312262 319744 312268 319796
rect 312320 319784 312326 319796
rect 312320 319756 312400 319784
rect 312320 319744 312326 319756
rect 312372 319660 312400 319756
rect 312602 319728 312630 319812
rect 312538 319676 312544 319728
rect 312596 319688 312630 319728
rect 312596 319676 312602 319688
rect 312694 319660 312722 319812
rect 312786 319716 312814 319812
rect 312786 319688 312860 319716
rect 312354 319608 312360 319660
rect 312412 319608 312418 319660
rect 312694 319620 312728 319660
rect 312722 319608 312728 319620
rect 312780 319608 312786 319660
rect 312832 319592 312860 319688
rect 312970 319648 312998 319824
rect 313062 319716 313090 319880
rect 313430 319784 313458 319880
rect 313384 319756 313458 319784
rect 313062 319688 313228 319716
rect 313090 319648 313096 319660
rect 312970 319620 313096 319648
rect 313090 319608 313096 319620
rect 313148 319608 313154 319660
rect 311866 319552 311900 319592
rect 311894 319540 311900 319552
rect 311952 319540 311958 319592
rect 312814 319540 312820 319592
rect 312872 319540 312878 319592
rect 311498 319484 311664 319512
rect 311636 319456 311664 319484
rect 305420 319416 305592 319444
rect 305420 319404 305426 319416
rect 309962 319404 309968 319456
rect 310020 319444 310026 319456
rect 310146 319444 310152 319456
rect 310020 319416 310152 319444
rect 310020 319404 310026 319416
rect 310146 319404 310152 319416
rect 310204 319404 310210 319456
rect 310790 319404 310796 319456
rect 310848 319444 310854 319456
rect 310848 319416 311480 319444
rect 310848 319404 310854 319416
rect 251450 319336 251456 319388
rect 251508 319376 251514 319388
rect 311342 319376 311348 319388
rect 251508 319348 311348 319376
rect 251508 319336 251514 319348
rect 311342 319336 311348 319348
rect 311400 319336 311406 319388
rect 311452 319376 311480 319416
rect 311618 319404 311624 319456
rect 311676 319404 311682 319456
rect 312262 319404 312268 319456
rect 312320 319444 312326 319456
rect 312630 319444 312636 319456
rect 312320 319416 312636 319444
rect 312320 319404 312326 319416
rect 312630 319404 312636 319416
rect 312688 319404 312694 319456
rect 312906 319404 312912 319456
rect 312964 319444 312970 319456
rect 313200 319444 313228 319688
rect 313384 319580 313412 319756
rect 313292 319552 313412 319580
rect 313292 319456 313320 319552
rect 312964 319416 313228 319444
rect 312964 319404 312970 319416
rect 313274 319404 313280 319456
rect 313332 319404 313338 319456
rect 313458 319404 313464 319456
rect 313516 319444 313522 319456
rect 313798 319444 313826 319880
rect 313872 319812 313878 319864
rect 313930 319812 313936 319864
rect 314056 319812 314062 319864
rect 314114 319812 314120 319864
rect 314626 319852 314654 320028
rect 314718 319920 314746 320164
rect 317156 319988 317184 320300
rect 336826 320288 336832 320300
rect 336884 320288 336890 320340
rect 327626 320220 327632 320272
rect 327684 320260 327690 320272
rect 335814 320260 335820 320272
rect 327684 320232 335820 320260
rect 327684 320220 327690 320232
rect 335814 320220 335820 320232
rect 335872 320220 335878 320272
rect 327534 320152 327540 320204
rect 327592 320192 327598 320204
rect 335906 320192 335912 320204
rect 327592 320164 335912 320192
rect 327592 320152 327598 320164
rect 335906 320152 335912 320164
rect 335964 320152 335970 320204
rect 321692 320084 321698 320136
rect 321750 320124 321756 320136
rect 331398 320124 331404 320136
rect 321750 320096 331404 320124
rect 321750 320084 321756 320096
rect 331398 320084 331404 320096
rect 331456 320084 331462 320136
rect 320864 320016 320870 320068
rect 320922 320056 320928 320068
rect 332962 320056 332968 320068
rect 320922 320028 332968 320056
rect 320922 320016 320928 320028
rect 332962 320016 332968 320028
rect 333020 320016 333026 320068
rect 333054 319988 333060 320000
rect 314902 319960 317184 319988
rect 321710 319960 333060 319988
rect 314792 319920 314798 319932
rect 314718 319892 314798 319920
rect 314792 319880 314798 319892
rect 314850 319880 314856 319932
rect 314902 319852 314930 319960
rect 315436 319880 315442 319932
rect 315494 319880 315500 319932
rect 315620 319880 315626 319932
rect 315678 319880 315684 319932
rect 316908 319880 316914 319932
rect 316966 319880 316972 319932
rect 317000 319880 317006 319932
rect 317058 319880 317064 319932
rect 319576 319880 319582 319932
rect 319634 319880 319640 319932
rect 320680 319920 320686 319932
rect 320422 319892 320686 319920
rect 314626 319824 314930 319852
rect 313890 319580 313918 319812
rect 314074 319648 314102 319812
rect 314074 319620 314332 319648
rect 314194 319580 314200 319592
rect 313890 319552 314200 319580
rect 314194 319540 314200 319552
rect 314252 319540 314258 319592
rect 313918 319472 313924 319524
rect 313976 319512 313982 319524
rect 314304 319512 314332 319620
rect 315298 319608 315304 319660
rect 315356 319648 315362 319660
rect 315454 319648 315482 319880
rect 315356 319620 315482 319648
rect 315638 319660 315666 319880
rect 316402 319812 316408 319864
rect 316460 319852 316466 319864
rect 316632 319852 316638 319864
rect 316460 319824 316638 319852
rect 316460 319812 316466 319824
rect 316632 319812 316638 319824
rect 316690 319812 316696 319864
rect 316218 319676 316224 319728
rect 316276 319716 316282 319728
rect 316926 319716 316954 319880
rect 317018 319784 317046 319880
rect 317386 319824 317966 319852
rect 317138 319784 317144 319796
rect 317018 319756 317144 319784
rect 317138 319744 317144 319756
rect 317196 319744 317202 319796
rect 316276 319688 316954 319716
rect 316276 319676 316282 319688
rect 315638 319620 315672 319660
rect 315356 319608 315362 319620
rect 315666 319608 315672 319620
rect 315724 319608 315730 319660
rect 316034 319608 316040 319660
rect 316092 319648 316098 319660
rect 317386 319648 317414 319824
rect 316092 319620 317414 319648
rect 317938 319648 317966 319824
rect 318196 319812 318202 319864
rect 318254 319852 318260 319864
rect 318886 319852 318892 319864
rect 318254 319824 318892 319852
rect 318254 319812 318260 319824
rect 318886 319812 318892 319824
rect 318944 319812 318950 319864
rect 319254 319812 319260 319864
rect 319312 319852 319318 319864
rect 319594 319852 319622 319880
rect 319312 319824 319622 319852
rect 319312 319812 319318 319824
rect 320312 319812 320318 319864
rect 320370 319812 320376 319864
rect 320330 319784 320358 319812
rect 320284 319756 320358 319784
rect 320284 319728 320312 319756
rect 320422 319728 320450 319892
rect 320680 319880 320686 319892
rect 320738 319880 320744 319932
rect 320588 319812 320594 319864
rect 320646 319812 320652 319864
rect 320606 319784 320634 319812
rect 321710 319784 321738 319960
rect 333054 319948 333060 319960
rect 333112 319948 333118 320000
rect 323532 319880 323538 319932
rect 323590 319880 323596 319932
rect 320606 319756 321738 319784
rect 323210 319744 323216 319796
rect 323268 319784 323274 319796
rect 323550 319784 323578 319880
rect 338206 319784 338212 319796
rect 323268 319756 323578 319784
rect 328426 319756 338212 319784
rect 323268 319744 323274 319756
rect 320266 319676 320272 319728
rect 320324 319676 320330 319728
rect 320358 319676 320364 319728
rect 320416 319688 320450 319728
rect 328426 319716 328454 319756
rect 338206 319744 338212 319756
rect 338264 319744 338270 319796
rect 340874 319716 340880 319728
rect 320560 319688 328454 319716
rect 328564 319688 340880 319716
rect 320416 319676 320422 319688
rect 320560 319648 320588 319688
rect 317938 319620 320588 319648
rect 316092 319608 316098 319620
rect 320634 319608 320640 319660
rect 320692 319648 320698 319660
rect 328454 319648 328460 319660
rect 320692 319620 328460 319648
rect 320692 319608 320698 319620
rect 328454 319608 328460 319620
rect 328512 319608 328518 319660
rect 322106 319512 322112 319524
rect 313976 319484 314332 319512
rect 316420 319484 322112 319512
rect 313976 319472 313982 319484
rect 313516 319416 313826 319444
rect 313516 319404 313522 319416
rect 314654 319376 314660 319388
rect 311452 319348 314660 319376
rect 314654 319336 314660 319348
rect 314712 319336 314718 319388
rect 243078 319268 243084 319320
rect 243136 319308 243142 319320
rect 302510 319308 302516 319320
rect 243136 319280 302516 319308
rect 243136 319268 243142 319280
rect 302510 319268 302516 319280
rect 302568 319268 302574 319320
rect 309778 319268 309784 319320
rect 309836 319308 309842 319320
rect 316034 319308 316040 319320
rect 309836 319280 316040 319308
rect 309836 319268 309842 319280
rect 316034 319268 316040 319280
rect 316092 319268 316098 319320
rect 248690 319200 248696 319252
rect 248748 319240 248754 319252
rect 309318 319240 309324 319252
rect 248748 319212 309324 319240
rect 248748 319200 248754 319212
rect 309318 319200 309324 319212
rect 309376 319200 309382 319252
rect 311710 319200 311716 319252
rect 311768 319240 311774 319252
rect 311894 319240 311900 319252
rect 311768 319212 311900 319240
rect 311768 319200 311774 319212
rect 311894 319200 311900 319212
rect 311952 319200 311958 319252
rect 248598 319132 248604 319184
rect 248656 319172 248662 319184
rect 309226 319172 309232 319184
rect 248656 319144 309232 319172
rect 248656 319132 248662 319144
rect 309226 319132 309232 319144
rect 309284 319132 309290 319184
rect 316420 319172 316448 319484
rect 322106 319472 322112 319484
rect 322164 319472 322170 319524
rect 323026 319472 323032 319524
rect 323084 319512 323090 319524
rect 323486 319512 323492 319524
rect 323084 319484 323492 319512
rect 323084 319472 323090 319484
rect 323486 319472 323492 319484
rect 323544 319472 323550 319524
rect 328564 319512 328592 319688
rect 340874 319676 340880 319688
rect 340932 319676 340938 319728
rect 323596 319484 328592 319512
rect 316494 319404 316500 319456
rect 316552 319444 316558 319456
rect 323596 319444 323624 319484
rect 316552 319416 323624 319444
rect 316552 319404 316558 319416
rect 325878 319404 325884 319456
rect 325936 319444 325942 319456
rect 326062 319444 326068 319456
rect 325936 319416 326068 319444
rect 325936 319404 325942 319416
rect 326062 319404 326068 319416
rect 326120 319404 326126 319456
rect 328426 319416 331214 319444
rect 322382 319336 322388 319388
rect 322440 319376 322446 319388
rect 328426 319376 328454 319416
rect 322440 319348 328454 319376
rect 331186 319376 331214 319416
rect 335998 319404 336004 319456
rect 336056 319444 336062 319456
rect 580442 319444 580448 319456
rect 336056 319416 580448 319444
rect 336056 319404 336062 319416
rect 580442 319404 580448 319416
rect 580500 319404 580506 319456
rect 337010 319376 337016 319388
rect 331186 319348 337016 319376
rect 322440 319336 322446 319348
rect 337010 319336 337016 319348
rect 337068 319336 337074 319388
rect 338482 319308 338488 319320
rect 309336 319144 316448 319172
rect 316512 319280 338488 319308
rect 283466 319064 283472 319116
rect 283524 319104 283530 319116
rect 292114 319104 292120 319116
rect 283524 319076 292120 319104
rect 283524 319064 283530 319076
rect 292114 319064 292120 319076
rect 292172 319064 292178 319116
rect 275278 318996 275284 319048
rect 275336 319036 275342 319048
rect 294598 319036 294604 319048
rect 275336 319008 294604 319036
rect 275336 318996 275342 319008
rect 294598 318996 294604 319008
rect 294656 318996 294662 319048
rect 295702 318996 295708 319048
rect 295760 319036 295766 319048
rect 296438 319036 296444 319048
rect 295760 319008 296444 319036
rect 295760 318996 295766 319008
rect 296438 318996 296444 319008
rect 296496 318996 296502 319048
rect 296530 318996 296536 319048
rect 296588 319036 296594 319048
rect 309336 319036 309364 319144
rect 310698 319064 310704 319116
rect 310756 319104 310762 319116
rect 316512 319104 316540 319280
rect 338482 319268 338488 319280
rect 338540 319268 338546 319320
rect 321278 319200 321284 319252
rect 321336 319240 321342 319252
rect 331582 319240 331588 319252
rect 321336 319212 331588 319240
rect 321336 319200 321342 319212
rect 331582 319200 331588 319212
rect 331640 319200 331646 319252
rect 332870 319172 332876 319184
rect 310756 319076 316540 319104
rect 318352 319144 332876 319172
rect 310756 319064 310762 319076
rect 296588 319008 309364 319036
rect 296588 318996 296594 319008
rect 314286 318996 314292 319048
rect 314344 319036 314350 319048
rect 318352 319036 318380 319144
rect 332870 319132 332876 319144
rect 332928 319132 332934 319184
rect 331214 319104 331220 319116
rect 314344 319008 318380 319036
rect 321526 319076 331220 319104
rect 314344 318996 314350 319008
rect 272978 318928 272984 318980
rect 273036 318968 273042 318980
rect 297358 318968 297364 318980
rect 273036 318940 297364 318968
rect 273036 318928 273042 318940
rect 297358 318928 297364 318940
rect 297416 318928 297422 318980
rect 309042 318928 309048 318980
rect 309100 318968 309106 318980
rect 321526 318968 321554 319076
rect 331214 319064 331220 319076
rect 331272 319064 331278 319116
rect 325326 318996 325332 319048
rect 325384 319036 325390 319048
rect 325510 319036 325516 319048
rect 325384 319008 325516 319036
rect 325384 318996 325390 319008
rect 325510 318996 325516 319008
rect 325568 318996 325574 319048
rect 326062 318996 326068 319048
rect 326120 319036 326126 319048
rect 326614 319036 326620 319048
rect 326120 319008 326620 319036
rect 326120 318996 326126 319008
rect 326614 318996 326620 319008
rect 326672 318996 326678 319048
rect 309100 318940 321554 318968
rect 309100 318928 309106 318940
rect 322566 318928 322572 318980
rect 322624 318968 322630 318980
rect 331950 318968 331956 318980
rect 322624 318940 331956 318968
rect 322624 318928 322630 318940
rect 331950 318928 331956 318940
rect 332008 318928 332014 318980
rect 279878 318860 279884 318912
rect 279936 318900 279942 318912
rect 295518 318900 295524 318912
rect 279936 318872 295524 318900
rect 279936 318860 279942 318872
rect 295518 318860 295524 318872
rect 295576 318860 295582 318912
rect 318242 318860 318248 318912
rect 318300 318900 318306 318912
rect 318426 318900 318432 318912
rect 318300 318872 318432 318900
rect 318300 318860 318306 318872
rect 318426 318860 318432 318872
rect 318484 318860 318490 318912
rect 320266 318860 320272 318912
rect 320324 318900 320330 318912
rect 330386 318900 330392 318912
rect 320324 318872 330392 318900
rect 320324 318860 320330 318872
rect 330386 318860 330392 318872
rect 330444 318860 330450 318912
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 3476 318804 244320 318832
rect 3476 318792 3482 318804
rect 244292 318764 244320 318804
rect 278038 318792 278044 318844
rect 278096 318832 278102 318844
rect 284202 318832 284208 318844
rect 278096 318804 284208 318832
rect 278096 318792 278102 318804
rect 284202 318792 284208 318804
rect 284260 318792 284266 318844
rect 286686 318792 286692 318844
rect 286744 318832 286750 318844
rect 286870 318832 286876 318844
rect 286744 318804 286876 318832
rect 286744 318792 286750 318804
rect 286870 318792 286876 318804
rect 286928 318792 286934 318844
rect 288710 318792 288716 318844
rect 288768 318832 288774 318844
rect 289722 318832 289728 318844
rect 288768 318804 289728 318832
rect 288768 318792 288774 318804
rect 289722 318792 289728 318804
rect 289780 318792 289786 318844
rect 290918 318792 290924 318844
rect 290976 318832 290982 318844
rect 291102 318832 291108 318844
rect 290976 318804 291108 318832
rect 290976 318792 290982 318804
rect 291102 318792 291108 318804
rect 291160 318792 291166 318844
rect 292114 318792 292120 318844
rect 292172 318832 292178 318844
rect 292172 318804 292574 318832
rect 292172 318792 292178 318804
rect 258166 318764 258172 318776
rect 244292 318736 258172 318764
rect 258166 318724 258172 318736
rect 258224 318764 258230 318776
rect 258810 318764 258816 318776
rect 258224 318736 258816 318764
rect 258224 318724 258230 318736
rect 258810 318724 258816 318736
rect 258868 318724 258874 318776
rect 285030 318724 285036 318776
rect 285088 318764 285094 318776
rect 285214 318764 285220 318776
rect 285088 318736 285220 318764
rect 285088 318724 285094 318736
rect 285214 318724 285220 318736
rect 285272 318724 285278 318776
rect 286318 318724 286324 318776
rect 286376 318764 286382 318776
rect 287514 318764 287520 318776
rect 286376 318736 287520 318764
rect 286376 318724 286382 318736
rect 287514 318724 287520 318736
rect 287572 318724 287578 318776
rect 289446 318724 289452 318776
rect 289504 318764 289510 318776
rect 289630 318764 289636 318776
rect 289504 318736 289636 318764
rect 289504 318724 289510 318736
rect 289630 318724 289636 318736
rect 289688 318724 289694 318776
rect 292546 318764 292574 318804
rect 292942 318792 292948 318844
rect 293000 318832 293006 318844
rect 293862 318832 293868 318844
rect 293000 318804 293868 318832
rect 293000 318792 293006 318804
rect 293862 318792 293868 318804
rect 293920 318792 293926 318844
rect 298094 318792 298100 318844
rect 298152 318832 298158 318844
rect 298278 318832 298284 318844
rect 298152 318804 298284 318832
rect 298152 318792 298158 318804
rect 298278 318792 298284 318804
rect 298336 318792 298342 318844
rect 302970 318792 302976 318844
rect 303028 318832 303034 318844
rect 303246 318832 303252 318844
rect 303028 318804 303252 318832
rect 303028 318792 303034 318804
rect 303246 318792 303252 318804
rect 303304 318792 303310 318844
rect 322198 318792 322204 318844
rect 322256 318832 322262 318844
rect 330018 318832 330024 318844
rect 322256 318804 330024 318832
rect 322256 318792 322262 318804
rect 330018 318792 330024 318804
rect 330076 318792 330082 318844
rect 293034 318764 293040 318776
rect 292546 318736 293040 318764
rect 293034 318724 293040 318736
rect 293092 318724 293098 318776
rect 293310 318724 293316 318776
rect 293368 318764 293374 318776
rect 293678 318764 293684 318776
rect 293368 318736 293684 318764
rect 293368 318724 293374 318736
rect 293678 318724 293684 318736
rect 293736 318724 293742 318776
rect 301038 318764 301044 318776
rect 293972 318736 301044 318764
rect 279602 318656 279608 318708
rect 279660 318696 279666 318708
rect 293972 318696 294000 318736
rect 301038 318724 301044 318736
rect 301096 318724 301102 318776
rect 318426 318724 318432 318776
rect 318484 318764 318490 318776
rect 318794 318764 318800 318776
rect 318484 318736 318800 318764
rect 318484 318724 318490 318736
rect 318794 318724 318800 318736
rect 318852 318724 318858 318776
rect 319898 318724 319904 318776
rect 319956 318764 319962 318776
rect 329834 318764 329840 318776
rect 319956 318736 329840 318764
rect 319956 318724 319962 318736
rect 329834 318724 329840 318736
rect 329892 318724 329898 318776
rect 279660 318668 294000 318696
rect 279660 318656 279666 318668
rect 294046 318656 294052 318708
rect 294104 318696 294110 318708
rect 294782 318696 294788 318708
rect 294104 318668 294788 318696
rect 294104 318656 294110 318668
rect 294782 318656 294788 318668
rect 294840 318656 294846 318708
rect 295886 318656 295892 318708
rect 295944 318696 295950 318708
rect 300762 318696 300768 318708
rect 295944 318668 300768 318696
rect 295944 318656 295950 318668
rect 300762 318656 300768 318668
rect 300820 318656 300826 318708
rect 319990 318656 319996 318708
rect 320048 318696 320054 318708
rect 330110 318696 330116 318708
rect 320048 318668 330116 318696
rect 320048 318656 320054 318668
rect 330110 318656 330116 318668
rect 330168 318656 330174 318708
rect 277578 318588 277584 318640
rect 277636 318628 277642 318640
rect 278406 318628 278412 318640
rect 277636 318600 278412 318628
rect 277636 318588 277642 318600
rect 278406 318588 278412 318600
rect 278464 318588 278470 318640
rect 282178 318588 282184 318640
rect 282236 318628 282242 318640
rect 285398 318628 285404 318640
rect 282236 318600 285404 318628
rect 282236 318588 282242 318600
rect 285398 318588 285404 318600
rect 285456 318588 285462 318640
rect 287790 318588 287796 318640
rect 287848 318628 287854 318640
rect 294966 318628 294972 318640
rect 287848 318600 294972 318628
rect 287848 318588 287854 318600
rect 294966 318588 294972 318600
rect 295024 318588 295030 318640
rect 298278 318588 298284 318640
rect 298336 318628 298342 318640
rect 299382 318628 299388 318640
rect 298336 318600 299388 318628
rect 298336 318588 298342 318600
rect 299382 318588 299388 318600
rect 299440 318588 299446 318640
rect 301038 318588 301044 318640
rect 301096 318628 301102 318640
rect 303798 318628 303804 318640
rect 301096 318600 303804 318628
rect 301096 318588 301102 318600
rect 303798 318588 303804 318600
rect 303856 318588 303862 318640
rect 312078 318588 312084 318640
rect 312136 318628 312142 318640
rect 323486 318628 323492 318640
rect 312136 318600 323492 318628
rect 312136 318588 312142 318600
rect 323486 318588 323492 318600
rect 323544 318588 323550 318640
rect 324958 318588 324964 318640
rect 325016 318628 325022 318640
rect 325602 318628 325608 318640
rect 325016 318600 325608 318628
rect 325016 318588 325022 318600
rect 325602 318588 325608 318600
rect 325660 318588 325666 318640
rect 326338 318588 326344 318640
rect 326396 318628 326402 318640
rect 334526 318628 334532 318640
rect 326396 318600 334532 318628
rect 326396 318588 326402 318600
rect 334526 318588 334532 318600
rect 334584 318588 334590 318640
rect 272886 318520 272892 318572
rect 272944 318560 272950 318572
rect 294046 318560 294052 318572
rect 272944 318532 294052 318560
rect 272944 318520 272950 318532
rect 294046 318520 294052 318532
rect 294104 318520 294110 318572
rect 295150 318520 295156 318572
rect 295208 318520 295214 318572
rect 295610 318520 295616 318572
rect 295668 318560 295674 318572
rect 300854 318560 300860 318572
rect 295668 318532 300860 318560
rect 295668 318520 295674 318532
rect 300854 318520 300860 318532
rect 300912 318520 300918 318572
rect 317322 318520 317328 318572
rect 317380 318560 317386 318572
rect 329098 318560 329104 318572
rect 317380 318532 329104 318560
rect 317380 318520 317386 318532
rect 329098 318520 329104 318532
rect 329156 318520 329162 318572
rect 247218 318452 247224 318504
rect 247276 318492 247282 318504
rect 282822 318492 282828 318504
rect 247276 318464 282828 318492
rect 247276 318452 247282 318464
rect 282822 318452 282828 318464
rect 282880 318452 282886 318504
rect 295168 318492 295196 318520
rect 286152 318464 295196 318492
rect 238846 318384 238852 318436
rect 238904 318424 238910 318436
rect 282270 318424 282276 318436
rect 238904 318396 282276 318424
rect 238904 318384 238910 318396
rect 282270 318384 282276 318396
rect 282328 318384 282334 318436
rect 282638 318384 282644 318436
rect 282696 318424 282702 318436
rect 286152 318424 286180 318464
rect 296622 318452 296628 318504
rect 296680 318492 296686 318504
rect 302050 318492 302056 318504
rect 296680 318464 302056 318492
rect 296680 318452 296686 318464
rect 302050 318452 302056 318464
rect 302108 318452 302114 318504
rect 317966 318452 317972 318504
rect 318024 318492 318030 318504
rect 325602 318492 325608 318504
rect 318024 318464 325608 318492
rect 318024 318452 318030 318464
rect 325602 318452 325608 318464
rect 325660 318452 325666 318504
rect 325786 318452 325792 318504
rect 325844 318492 325850 318504
rect 335722 318492 335728 318504
rect 325844 318464 335728 318492
rect 325844 318452 325850 318464
rect 335722 318452 335728 318464
rect 335780 318452 335786 318504
rect 282696 318396 286180 318424
rect 282696 318384 282702 318396
rect 289446 318384 289452 318436
rect 289504 318424 289510 318436
rect 289504 318396 294874 318424
rect 289504 318384 289510 318396
rect 209682 318316 209688 318368
rect 209740 318356 209746 318368
rect 283742 318356 283748 318368
rect 209740 318328 283748 318356
rect 209740 318316 209746 318328
rect 283742 318316 283748 318328
rect 283800 318316 283806 318368
rect 284846 318316 284852 318368
rect 284904 318356 284910 318368
rect 285122 318356 285128 318368
rect 284904 318328 285128 318356
rect 284904 318316 284910 318328
rect 285122 318316 285128 318328
rect 285180 318316 285186 318368
rect 291930 318316 291936 318368
rect 291988 318356 291994 318368
rect 294414 318356 294420 318368
rect 291988 318328 294420 318356
rect 291988 318316 291994 318328
rect 294414 318316 294420 318328
rect 294472 318316 294478 318368
rect 294846 318356 294874 318396
rect 295150 318384 295156 318436
rect 295208 318424 295214 318436
rect 303430 318424 303436 318436
rect 295208 318396 303436 318424
rect 295208 318384 295214 318396
rect 303430 318384 303436 318396
rect 303488 318384 303494 318436
rect 317414 318384 317420 318436
rect 317472 318424 317478 318436
rect 326522 318424 326528 318436
rect 317472 318396 326528 318424
rect 317472 318384 317478 318396
rect 326522 318384 326528 318396
rect 326580 318384 326586 318436
rect 297082 318356 297088 318368
rect 294846 318328 297088 318356
rect 297082 318316 297088 318328
rect 297140 318316 297146 318368
rect 300854 318316 300860 318368
rect 300912 318356 300918 318368
rect 302234 318356 302240 318368
rect 300912 318328 302240 318356
rect 300912 318316 300918 318328
rect 302234 318316 302240 318328
rect 302292 318316 302298 318368
rect 318886 318316 318892 318368
rect 318944 318356 318950 318368
rect 335538 318356 335544 318368
rect 318944 318328 335544 318356
rect 318944 318316 318950 318328
rect 335538 318316 335544 318328
rect 335596 318316 335602 318368
rect 212258 318248 212264 318300
rect 212316 318288 212322 318300
rect 286226 318288 286232 318300
rect 212316 318260 286232 318288
rect 212316 318248 212322 318260
rect 286226 318248 286232 318260
rect 286284 318248 286290 318300
rect 292114 318248 292120 318300
rect 292172 318288 292178 318300
rect 299934 318288 299940 318300
rect 292172 318260 299940 318288
rect 292172 318248 292178 318260
rect 299934 318248 299940 318260
rect 299992 318248 299998 318300
rect 300210 318248 300216 318300
rect 300268 318288 300274 318300
rect 300762 318288 300768 318300
rect 300268 318260 300768 318288
rect 300268 318248 300274 318260
rect 300762 318248 300768 318260
rect 300820 318248 300826 318300
rect 311802 318248 311808 318300
rect 311860 318288 311866 318300
rect 326338 318288 326344 318300
rect 311860 318260 326344 318288
rect 311860 318248 311866 318260
rect 326338 318248 326344 318260
rect 326396 318248 326402 318300
rect 287238 318220 287244 318232
rect 273226 318192 287244 318220
rect 218974 318112 218980 318164
rect 219032 318152 219038 318164
rect 273226 318152 273254 318192
rect 287238 318180 287244 318192
rect 287296 318180 287302 318232
rect 288802 318180 288808 318232
rect 288860 318220 288866 318232
rect 289262 318220 289268 318232
rect 288860 318192 289268 318220
rect 288860 318180 288866 318192
rect 289262 318180 289268 318192
rect 289320 318180 289326 318232
rect 290734 318180 290740 318232
rect 290792 318220 290798 318232
rect 298094 318220 298100 318232
rect 290792 318192 298100 318220
rect 290792 318180 290798 318192
rect 298094 318180 298100 318192
rect 298152 318180 298158 318232
rect 299290 318180 299296 318232
rect 299348 318220 299354 318232
rect 306650 318220 306656 318232
rect 299348 318192 306656 318220
rect 299348 318180 299354 318192
rect 306650 318180 306656 318192
rect 306708 318180 306714 318232
rect 319346 318180 319352 318232
rect 319404 318220 319410 318232
rect 319404 318192 323808 318220
rect 319404 318180 319410 318192
rect 219032 318124 273254 318152
rect 219032 318112 219038 318124
rect 286226 318112 286232 318164
rect 286284 318152 286290 318164
rect 286778 318152 286784 318164
rect 286284 318124 286784 318152
rect 286284 318112 286290 318124
rect 286778 318112 286784 318124
rect 286836 318112 286842 318164
rect 295978 318152 295984 318164
rect 287900 318124 295984 318152
rect 219066 318044 219072 318096
rect 219124 318084 219130 318096
rect 287790 318084 287796 318096
rect 219124 318056 287796 318084
rect 219124 318044 219130 318056
rect 287790 318044 287796 318056
rect 287848 318044 287854 318096
rect 287238 317976 287244 318028
rect 287296 318016 287302 318028
rect 287900 318016 287928 318124
rect 295978 318112 295984 318124
rect 296036 318112 296042 318164
rect 300210 318112 300216 318164
rect 300268 318152 300274 318164
rect 302786 318152 302792 318164
rect 300268 318124 302792 318152
rect 300268 318112 300274 318124
rect 302786 318112 302792 318124
rect 302844 318112 302850 318164
rect 316586 318112 316592 318164
rect 316644 318152 316650 318164
rect 316644 318124 323624 318152
rect 316644 318112 316650 318124
rect 294046 318044 294052 318096
rect 294104 318084 294110 318096
rect 301774 318084 301780 318096
rect 294104 318056 301780 318084
rect 294104 318044 294110 318056
rect 301774 318044 301780 318056
rect 301832 318044 301838 318096
rect 287296 317988 287928 318016
rect 287296 317976 287302 317988
rect 288802 317976 288808 318028
rect 288860 318016 288866 318028
rect 289078 318016 289084 318028
rect 288860 317988 289084 318016
rect 288860 317976 288866 317988
rect 289078 317976 289084 317988
rect 289136 317976 289142 318028
rect 295334 317976 295340 318028
rect 295392 318016 295398 318028
rect 301498 318016 301504 318028
rect 295392 317988 301504 318016
rect 295392 317976 295398 317988
rect 301498 317976 301504 317988
rect 301556 317976 301562 318028
rect 309778 317976 309784 318028
rect 309836 318016 309842 318028
rect 312538 318016 312544 318028
rect 309836 317988 312544 318016
rect 309836 317976 309842 317988
rect 312538 317976 312544 317988
rect 312596 317976 312602 318028
rect 313366 317976 313372 318028
rect 313424 318016 313430 318028
rect 313424 317988 321554 318016
rect 313424 317976 313430 317988
rect 278130 317908 278136 317960
rect 278188 317948 278194 317960
rect 295426 317948 295432 317960
rect 278188 317920 295432 317948
rect 278188 317908 278194 317920
rect 295426 317908 295432 317920
rect 295484 317908 295490 317960
rect 303430 317908 303436 317960
rect 303488 317948 303494 317960
rect 304350 317948 304356 317960
rect 303488 317920 304356 317948
rect 303488 317908 303494 317920
rect 304350 317908 304356 317920
rect 304408 317908 304414 317960
rect 311802 317908 311808 317960
rect 311860 317948 311866 317960
rect 314010 317948 314016 317960
rect 311860 317920 314016 317948
rect 311860 317908 311866 317920
rect 314010 317908 314016 317920
rect 314068 317908 314074 317960
rect 321526 317948 321554 317988
rect 322382 317948 322388 317960
rect 321526 317920 322388 317948
rect 322382 317908 322388 317920
rect 322440 317908 322446 317960
rect 323596 317948 323624 318124
rect 323780 318084 323808 318192
rect 326430 318180 326436 318232
rect 326488 318220 326494 318232
rect 340966 318220 340972 318232
rect 326488 318192 340972 318220
rect 326488 318180 326494 318192
rect 340966 318180 340972 318192
rect 341024 318180 341030 318232
rect 326522 318112 326528 318164
rect 326580 318152 326586 318164
rect 349246 318152 349252 318164
rect 326580 318124 349252 318152
rect 326580 318112 326586 318124
rect 349246 318112 349252 318124
rect 349304 318112 349310 318164
rect 354674 318084 354680 318096
rect 323780 318056 354680 318084
rect 354674 318044 354680 318056
rect 354732 318044 354738 318096
rect 325602 317976 325608 318028
rect 325660 318016 325666 318028
rect 330570 318016 330576 318028
rect 325660 317988 330576 318016
rect 325660 317976 325666 317988
rect 330570 317976 330576 317988
rect 330628 317976 330634 318028
rect 326430 317948 326436 317960
rect 323596 317920 326436 317948
rect 326430 317908 326436 317920
rect 326488 317908 326494 317960
rect 286778 317840 286784 317892
rect 286836 317880 286842 317892
rect 293402 317880 293408 317892
rect 286836 317852 293408 317880
rect 286836 317840 286842 317852
rect 293402 317840 293408 317852
rect 293460 317840 293466 317892
rect 293862 317840 293868 317892
rect 293920 317880 293926 317892
rect 298462 317880 298468 317892
rect 293920 317852 298468 317880
rect 293920 317840 293926 317852
rect 298462 317840 298468 317852
rect 298520 317840 298526 317892
rect 312262 317840 312268 317892
rect 312320 317880 312326 317892
rect 326522 317880 326528 317892
rect 312320 317852 326528 317880
rect 312320 317840 312326 317852
rect 326522 317840 326528 317852
rect 326580 317840 326586 317892
rect 283742 317772 283748 317824
rect 283800 317812 283806 317824
rect 292298 317812 292304 317824
rect 283800 317784 292304 317812
rect 283800 317772 283806 317784
rect 292298 317772 292304 317784
rect 292356 317772 292362 317824
rect 294782 317772 294788 317824
rect 294840 317812 294846 317824
rect 298738 317812 298744 317824
rect 294840 317784 298744 317812
rect 294840 317772 294846 317784
rect 298738 317772 298744 317784
rect 298796 317772 298802 317824
rect 300026 317772 300032 317824
rect 300084 317812 300090 317824
rect 300302 317812 300308 317824
rect 300084 317784 300308 317812
rect 300084 317772 300090 317784
rect 300302 317772 300308 317784
rect 300360 317772 300366 317824
rect 301406 317772 301412 317824
rect 301464 317812 301470 317824
rect 302878 317812 302884 317824
rect 301464 317784 302884 317812
rect 301464 317772 301470 317784
rect 302878 317772 302884 317784
rect 302936 317772 302942 317824
rect 303798 317812 303804 317824
rect 302988 317784 303804 317812
rect 221734 317704 221740 317756
rect 221792 317744 221798 317756
rect 296622 317744 296628 317756
rect 221792 317716 296628 317744
rect 221792 317704 221798 317716
rect 296622 317704 296628 317716
rect 296680 317704 296686 317756
rect 297358 317704 297364 317756
rect 297416 317744 297422 317756
rect 301130 317744 301136 317756
rect 297416 317716 301136 317744
rect 297416 317704 297422 317716
rect 301130 317704 301136 317716
rect 301188 317704 301194 317756
rect 301222 317704 301228 317756
rect 301280 317744 301286 317756
rect 302988 317744 303016 317784
rect 303798 317772 303804 317784
rect 303856 317772 303862 317824
rect 307110 317744 307116 317756
rect 301280 317716 303016 317744
rect 303908 317716 307116 317744
rect 301280 317704 301286 317716
rect 276934 317636 276940 317688
rect 276992 317676 276998 317688
rect 295334 317676 295340 317688
rect 276992 317648 295340 317676
rect 276992 317636 276998 317648
rect 295334 317636 295340 317648
rect 295392 317636 295398 317688
rect 296254 317636 296260 317688
rect 296312 317676 296318 317688
rect 299566 317676 299572 317688
rect 296312 317648 299572 317676
rect 296312 317636 296318 317648
rect 299566 317636 299572 317648
rect 299624 317636 299630 317688
rect 301958 317636 301964 317688
rect 302016 317676 302022 317688
rect 303908 317676 303936 317716
rect 307110 317704 307116 317716
rect 307168 317704 307174 317756
rect 302016 317648 303936 317676
rect 302016 317636 302022 317648
rect 303982 317636 303988 317688
rect 304040 317676 304046 317688
rect 305270 317676 305276 317688
rect 304040 317648 305276 317676
rect 304040 317636 304046 317648
rect 305270 317636 305276 317648
rect 305328 317636 305334 317688
rect 305822 317636 305828 317688
rect 305880 317636 305886 317688
rect 320726 317636 320732 317688
rect 320784 317676 320790 317688
rect 321370 317676 321376 317688
rect 320784 317648 321376 317676
rect 320784 317636 320790 317648
rect 321370 317636 321376 317648
rect 321428 317636 321434 317688
rect 280614 317568 280620 317620
rect 280672 317608 280678 317620
rect 283742 317608 283748 317620
rect 280672 317580 283748 317608
rect 280672 317568 280678 317580
rect 283742 317568 283748 317580
rect 283800 317568 283806 317620
rect 283926 317568 283932 317620
rect 283984 317608 283990 317620
rect 290642 317608 290648 317620
rect 283984 317580 290648 317608
rect 283984 317568 283990 317580
rect 290642 317568 290648 317580
rect 290700 317568 290706 317620
rect 293402 317568 293408 317620
rect 293460 317608 293466 317620
rect 295058 317608 295064 317620
rect 293460 317580 295064 317608
rect 293460 317568 293466 317580
rect 295058 317568 295064 317580
rect 295116 317568 295122 317620
rect 296070 317568 296076 317620
rect 296128 317608 296134 317620
rect 298370 317608 298376 317620
rect 296128 317580 298376 317608
rect 296128 317568 296134 317580
rect 298370 317568 298376 317580
rect 298428 317568 298434 317620
rect 300302 317568 300308 317620
rect 300360 317608 300366 317620
rect 305840 317608 305868 317636
rect 300360 317580 305868 317608
rect 300360 317568 300366 317580
rect 306098 317568 306104 317620
rect 306156 317608 306162 317620
rect 306282 317608 306288 317620
rect 306156 317580 306288 317608
rect 306156 317568 306162 317580
rect 306282 317568 306288 317580
rect 306340 317568 306346 317620
rect 308490 317568 308496 317620
rect 308548 317608 308554 317620
rect 308950 317608 308956 317620
rect 308548 317580 308956 317608
rect 308548 317568 308554 317580
rect 308950 317568 308956 317580
rect 309008 317568 309014 317620
rect 323394 317568 323400 317620
rect 323452 317608 323458 317620
rect 327810 317608 327816 317620
rect 323452 317580 327816 317608
rect 323452 317568 323458 317580
rect 327810 317568 327816 317580
rect 327868 317568 327874 317620
rect 283650 317500 283656 317552
rect 283708 317540 283714 317552
rect 289538 317540 289544 317552
rect 283708 317512 289544 317540
rect 283708 317500 283714 317512
rect 289538 317500 289544 317512
rect 289596 317500 289602 317552
rect 295886 317540 295892 317552
rect 292546 317512 295892 317540
rect 272794 317432 272800 317484
rect 272852 317472 272858 317484
rect 292546 317472 292574 317512
rect 295886 317500 295892 317512
rect 295944 317500 295950 317552
rect 298186 317500 298192 317552
rect 298244 317540 298250 317552
rect 300118 317540 300124 317552
rect 298244 317512 300124 317540
rect 298244 317500 298250 317512
rect 300118 317500 300124 317512
rect 300176 317500 300182 317552
rect 303062 317500 303068 317552
rect 303120 317540 303126 317552
rect 305454 317540 305460 317552
rect 303120 317512 305460 317540
rect 303120 317500 303126 317512
rect 305454 317500 305460 317512
rect 305512 317500 305518 317552
rect 305822 317500 305828 317552
rect 305880 317540 305886 317552
rect 308030 317540 308036 317552
rect 305880 317512 308036 317540
rect 305880 317500 305886 317512
rect 308030 317500 308036 317512
rect 308088 317500 308094 317552
rect 313274 317500 313280 317552
rect 313332 317540 313338 317552
rect 320726 317540 320732 317552
rect 313332 317512 320732 317540
rect 313332 317500 313338 317512
rect 320726 317500 320732 317512
rect 320784 317500 320790 317552
rect 324406 317500 324412 317552
rect 324464 317540 324470 317552
rect 327626 317540 327632 317552
rect 324464 317512 327632 317540
rect 324464 317500 324470 317512
rect 327626 317500 327632 317512
rect 327684 317500 327690 317552
rect 272852 317444 292574 317472
rect 272852 317432 272858 317444
rect 295334 317432 295340 317484
rect 295392 317472 295398 317484
rect 297266 317472 297272 317484
rect 295392 317444 297272 317472
rect 295392 317432 295398 317444
rect 297266 317432 297272 317444
rect 297324 317432 297330 317484
rect 298830 317432 298836 317484
rect 298888 317472 298894 317484
rect 300486 317472 300492 317484
rect 298888 317444 300492 317472
rect 298888 317432 298894 317444
rect 300486 317432 300492 317444
rect 300544 317432 300550 317484
rect 303798 317432 303804 317484
rect 303856 317472 303862 317484
rect 303982 317472 303988 317484
rect 303856 317444 303988 317472
rect 303856 317432 303862 317444
rect 303982 317432 303988 317444
rect 304040 317432 304046 317484
rect 307570 317432 307576 317484
rect 307628 317472 307634 317484
rect 308214 317472 308220 317484
rect 307628 317444 308220 317472
rect 307628 317432 307634 317444
rect 308214 317432 308220 317444
rect 308272 317432 308278 317484
rect 308950 317432 308956 317484
rect 309008 317472 309014 317484
rect 309594 317472 309600 317484
rect 309008 317444 309600 317472
rect 309008 317432 309014 317444
rect 309594 317432 309600 317444
rect 309652 317432 309658 317484
rect 314562 317432 314568 317484
rect 314620 317472 314626 317484
rect 315114 317472 315120 317484
rect 314620 317444 315120 317472
rect 314620 317432 314626 317444
rect 315114 317432 315120 317444
rect 315172 317432 315178 317484
rect 315666 317432 315672 317484
rect 315724 317472 315730 317484
rect 317966 317472 317972 317484
rect 315724 317444 317972 317472
rect 315724 317432 315730 317444
rect 317966 317432 317972 317444
rect 318024 317432 318030 317484
rect 326154 317432 326160 317484
rect 326212 317472 326218 317484
rect 327534 317472 327540 317484
rect 326212 317444 327540 317472
rect 326212 317432 326218 317444
rect 327534 317432 327540 317444
rect 327592 317432 327598 317484
rect 279786 317364 279792 317416
rect 279844 317404 279850 317416
rect 302142 317404 302148 317416
rect 279844 317376 302148 317404
rect 279844 317364 279850 317376
rect 302142 317364 302148 317376
rect 302200 317364 302206 317416
rect 318702 317364 318708 317416
rect 318760 317404 318766 317416
rect 323394 317404 323400 317416
rect 318760 317376 323400 317404
rect 318760 317364 318766 317376
rect 323394 317364 323400 317376
rect 323452 317364 323458 317416
rect 274174 317296 274180 317348
rect 274232 317336 274238 317348
rect 296346 317336 296352 317348
rect 274232 317308 296352 317336
rect 274232 317296 274238 317308
rect 296346 317296 296352 317308
rect 296404 317296 296410 317348
rect 322934 317296 322940 317348
rect 322992 317336 322998 317348
rect 328730 317336 328736 317348
rect 322992 317308 328736 317336
rect 322992 317296 322998 317308
rect 328730 317296 328736 317308
rect 328788 317296 328794 317348
rect 274266 317228 274272 317280
rect 274324 317268 274330 317280
rect 296806 317268 296812 317280
rect 274324 317240 296812 317268
rect 274324 317228 274330 317240
rect 296806 317228 296812 317240
rect 296864 317228 296870 317280
rect 271414 317092 271420 317144
rect 271472 317132 271478 317144
rect 295794 317132 295800 317144
rect 271472 317104 295800 317132
rect 271472 317092 271478 317104
rect 295794 317092 295800 317104
rect 295852 317092 295858 317144
rect 295978 317092 295984 317144
rect 296036 317132 296042 317144
rect 305638 317132 305644 317144
rect 296036 317104 305644 317132
rect 296036 317092 296042 317104
rect 305638 317092 305644 317104
rect 305696 317092 305702 317144
rect 273990 317024 273996 317076
rect 274048 317064 274054 317076
rect 303614 317064 303620 317076
rect 274048 317036 303620 317064
rect 274048 317024 274054 317036
rect 303614 317024 303620 317036
rect 303672 317024 303678 317076
rect 317690 317024 317696 317076
rect 317748 317064 317754 317076
rect 334066 317064 334072 317076
rect 317748 317036 334072 317064
rect 317748 317024 317754 317036
rect 334066 317024 334072 317036
rect 334124 317024 334130 317076
rect 273162 316956 273168 317008
rect 273220 316996 273226 317008
rect 303706 316996 303712 317008
rect 273220 316968 303712 316996
rect 273220 316956 273226 316968
rect 303706 316956 303712 316968
rect 303764 316956 303770 317008
rect 308858 316956 308864 317008
rect 308916 316996 308922 317008
rect 328822 316996 328828 317008
rect 308916 316968 328828 316996
rect 308916 316956 308922 316968
rect 328822 316956 328828 316968
rect 328880 316956 328886 317008
rect 271506 316888 271512 316940
rect 271564 316928 271570 316940
rect 302602 316928 302608 316940
rect 271564 316900 302608 316928
rect 271564 316888 271570 316900
rect 302602 316888 302608 316900
rect 302660 316888 302666 316940
rect 308306 316888 308312 316940
rect 308364 316928 308370 316940
rect 329926 316928 329932 316940
rect 308364 316900 329932 316928
rect 308364 316888 308370 316900
rect 329926 316888 329932 316900
rect 329984 316888 329990 316940
rect 277302 316820 277308 316872
rect 277360 316860 277366 316872
rect 313734 316860 313740 316872
rect 277360 316832 313740 316860
rect 277360 316820 277366 316832
rect 313734 316820 313740 316832
rect 313792 316820 313798 316872
rect 316678 316820 316684 316872
rect 316736 316860 316742 316872
rect 336918 316860 336924 316872
rect 316736 316832 336924 316860
rect 316736 316820 316742 316832
rect 336918 316820 336924 316832
rect 336976 316820 336982 316872
rect 218790 316752 218796 316804
rect 218848 316792 218854 316804
rect 294598 316792 294604 316804
rect 218848 316764 294604 316792
rect 218848 316752 218854 316764
rect 294598 316752 294604 316764
rect 294656 316752 294662 316804
rect 295242 316752 295248 316804
rect 295300 316792 295306 316804
rect 304994 316792 305000 316804
rect 295300 316764 305000 316792
rect 295300 316752 295306 316764
rect 304994 316752 305000 316764
rect 305052 316752 305058 316804
rect 364334 316792 364340 316804
rect 311866 316764 364340 316792
rect 213362 316684 213368 316736
rect 213420 316724 213426 316736
rect 293862 316724 293868 316736
rect 213420 316696 293868 316724
rect 213420 316684 213426 316696
rect 293862 316684 293868 316696
rect 293920 316684 293926 316736
rect 296622 316684 296628 316736
rect 296680 316724 296686 316736
rect 296680 316696 304350 316724
rect 296680 316684 296686 316696
rect 282822 316616 282828 316668
rect 282880 316656 282886 316668
rect 303430 316656 303436 316668
rect 282880 316628 303436 316656
rect 282880 316616 282886 316628
rect 303430 316616 303436 316628
rect 303488 316616 303494 316668
rect 304322 316656 304350 316696
rect 308306 316684 308312 316736
rect 308364 316724 308370 316736
rect 310790 316724 310796 316736
rect 308364 316696 310796 316724
rect 308364 316684 308370 316696
rect 310790 316684 310796 316696
rect 310848 316724 310854 316736
rect 311866 316724 311894 316764
rect 364334 316752 364340 316764
rect 364392 316752 364398 316804
rect 310848 316696 311894 316724
rect 310848 316684 310854 316696
rect 323578 316684 323584 316736
rect 323636 316724 323642 316736
rect 400858 316724 400864 316736
rect 323636 316696 400864 316724
rect 323636 316684 323642 316696
rect 400858 316684 400864 316696
rect 400916 316684 400922 316736
rect 320450 316656 320456 316668
rect 304322 316628 320456 316656
rect 320450 316616 320456 316628
rect 320508 316616 320514 316668
rect 276842 316548 276848 316600
rect 276900 316588 276906 316600
rect 293954 316588 293960 316600
rect 276900 316560 293960 316588
rect 276900 316548 276906 316560
rect 293954 316548 293960 316560
rect 294012 316548 294018 316600
rect 280982 316480 280988 316532
rect 281040 316520 281046 316532
rect 292390 316520 292396 316532
rect 281040 316492 292396 316520
rect 281040 316480 281046 316492
rect 292390 316480 292396 316492
rect 292448 316480 292454 316532
rect 271322 316412 271328 316464
rect 271380 316452 271386 316464
rect 294322 316452 294328 316464
rect 271380 316424 294328 316452
rect 271380 316412 271386 316424
rect 294322 316412 294328 316424
rect 294380 316412 294386 316464
rect 325234 316412 325240 316464
rect 325292 316452 325298 316464
rect 325292 316424 331214 316452
rect 325292 316412 325298 316424
rect 324958 316276 324964 316328
rect 325016 316316 325022 316328
rect 327902 316316 327908 316328
rect 325016 316288 327908 316316
rect 325016 316276 325022 316288
rect 327902 316276 327908 316288
rect 327960 316276 327966 316328
rect 284294 316208 284300 316260
rect 284352 316248 284358 316260
rect 284846 316248 284852 316260
rect 284352 316220 284852 316248
rect 284352 316208 284358 316220
rect 284846 316208 284852 316220
rect 284904 316208 284910 316260
rect 309594 316208 309600 316260
rect 309652 316248 309658 316260
rect 310238 316248 310244 316260
rect 309652 316220 310244 316248
rect 309652 316208 309658 316220
rect 310238 316208 310244 316220
rect 310296 316208 310302 316260
rect 322198 316208 322204 316260
rect 322256 316248 322262 316260
rect 323578 316248 323584 316260
rect 322256 316220 323584 316248
rect 322256 316208 322262 316220
rect 323578 316208 323584 316220
rect 323636 316208 323642 316260
rect 324038 316208 324044 316260
rect 324096 316248 324102 316260
rect 331186 316248 331214 316424
rect 493318 316248 493324 316260
rect 324096 316220 326292 316248
rect 331186 316220 493324 316248
rect 324096 316208 324102 316220
rect 284754 316140 284760 316192
rect 284812 316180 284818 316192
rect 285490 316180 285496 316192
rect 284812 316152 285496 316180
rect 284812 316140 284818 316152
rect 285490 316140 285496 316152
rect 285548 316140 285554 316192
rect 306834 316140 306840 316192
rect 306892 316180 306898 316192
rect 307018 316180 307024 316192
rect 306892 316152 307024 316180
rect 306892 316140 306898 316152
rect 307018 316140 307024 316152
rect 307076 316140 307082 316192
rect 323854 316140 323860 316192
rect 323912 316180 323918 316192
rect 324130 316180 324136 316192
rect 323912 316152 324136 316180
rect 323912 316140 323918 316152
rect 324130 316140 324136 316152
rect 324188 316140 324194 316192
rect 325050 316140 325056 316192
rect 325108 316180 325114 316192
rect 325234 316180 325240 316192
rect 325108 316152 325240 316180
rect 325108 316140 325114 316152
rect 325234 316140 325240 316152
rect 325292 316140 325298 316192
rect 326264 316180 326292 316220
rect 493318 316208 493324 316220
rect 493376 316208 493382 316260
rect 534074 316180 534080 316192
rect 326264 316152 534080 316180
rect 534074 316140 534080 316152
rect 534132 316140 534138 316192
rect 283098 316072 283104 316124
rect 283156 316112 283162 316124
rect 284110 316112 284116 316124
rect 283156 316084 284116 316112
rect 283156 316072 283162 316084
rect 284110 316072 284116 316084
rect 284168 316072 284174 316124
rect 284662 316072 284668 316124
rect 284720 316112 284726 316124
rect 285582 316112 285588 316124
rect 284720 316084 285588 316112
rect 284720 316072 284726 316084
rect 285582 316072 285588 316084
rect 285640 316072 285646 316124
rect 287330 316072 287336 316124
rect 287388 316112 287394 316124
rect 287882 316112 287888 316124
rect 287388 316084 287888 316112
rect 287388 316072 287394 316084
rect 287882 316072 287888 316084
rect 287940 316072 287946 316124
rect 288526 316072 288532 316124
rect 288584 316112 288590 316124
rect 289354 316112 289360 316124
rect 288584 316084 289360 316112
rect 288584 316072 288590 316084
rect 289354 316072 289360 316084
rect 289412 316072 289418 316124
rect 290182 316072 290188 316124
rect 290240 316112 290246 316124
rect 290458 316112 290464 316124
rect 290240 316084 290464 316112
rect 290240 316072 290246 316084
rect 290458 316072 290464 316084
rect 290516 316072 290522 316124
rect 295610 316112 295616 316124
rect 292408 316084 295616 316112
rect 283006 316004 283012 316056
rect 283064 316044 283070 316056
rect 283834 316044 283840 316056
rect 283064 316016 283840 316044
rect 283064 316004 283070 316016
rect 283834 316004 283840 316016
rect 283892 316004 283898 316056
rect 284846 316004 284852 316056
rect 284904 316044 284910 316056
rect 285306 316044 285312 316056
rect 284904 316016 285312 316044
rect 284904 316004 284910 316016
rect 285306 316004 285312 316016
rect 285364 316004 285370 316056
rect 285674 316004 285680 316056
rect 285732 316044 285738 316056
rect 286870 316044 286876 316056
rect 285732 316016 286876 316044
rect 285732 316004 285738 316016
rect 286870 316004 286876 316016
rect 286928 316004 286934 316056
rect 287238 316004 287244 316056
rect 287296 316044 287302 316056
rect 288158 316044 288164 316056
rect 287296 316016 288164 316044
rect 287296 316004 287302 316016
rect 288158 316004 288164 316016
rect 288216 316004 288222 316056
rect 288618 316004 288624 316056
rect 288676 316044 288682 316056
rect 289170 316044 289176 316056
rect 288676 316016 289176 316044
rect 288676 316004 288682 316016
rect 289170 316004 289176 316016
rect 289228 316004 289234 316056
rect 289906 316004 289912 316056
rect 289964 316044 289970 316056
rect 290734 316044 290740 316056
rect 289964 316016 290740 316044
rect 289964 316004 289970 316016
rect 290734 316004 290740 316016
rect 290792 316004 290798 316056
rect 291470 316004 291476 316056
rect 291528 316044 291534 316056
rect 292022 316044 292028 316056
rect 291528 316016 292028 316044
rect 291528 316004 291534 316016
rect 292022 316004 292028 316016
rect 292080 316004 292086 316056
rect 275554 315936 275560 315988
rect 275612 315976 275618 315988
rect 290642 315976 290648 315988
rect 275612 315948 290648 315976
rect 275612 315936 275618 315948
rect 290642 315936 290648 315948
rect 290700 315936 290706 315988
rect 276750 315868 276756 315920
rect 276808 315908 276814 315920
rect 292408 315908 292436 316084
rect 295610 316072 295616 316084
rect 295668 316072 295674 316124
rect 309410 316072 309416 316124
rect 309468 316112 309474 316124
rect 310238 316112 310244 316124
rect 309468 316084 310244 316112
rect 309468 316072 309474 316084
rect 310238 316072 310244 316084
rect 310296 316072 310302 316124
rect 311526 316072 311532 316124
rect 311584 316112 311590 316124
rect 311710 316112 311716 316124
rect 311584 316084 311716 316112
rect 311584 316072 311590 316084
rect 311710 316072 311716 316084
rect 311768 316072 311774 316124
rect 315482 316072 315488 316124
rect 315540 316112 315546 316124
rect 315758 316112 315764 316124
rect 315540 316084 315764 316112
rect 315540 316072 315546 316084
rect 315758 316072 315764 316084
rect 315816 316072 315822 316124
rect 323578 316072 323584 316124
rect 323636 316112 323642 316124
rect 324038 316112 324044 316124
rect 323636 316084 324044 316112
rect 323636 316072 323642 316084
rect 324038 316072 324044 316084
rect 324096 316072 324102 316124
rect 325142 316072 325148 316124
rect 325200 316112 325206 316124
rect 547966 316112 547972 316124
rect 325200 316084 547972 316112
rect 325200 316072 325206 316084
rect 547966 316072 547972 316084
rect 548024 316072 548030 316124
rect 294230 316004 294236 316056
rect 294288 316044 294294 316056
rect 294506 316044 294512 316056
rect 294288 316016 294512 316044
rect 294288 316004 294294 316016
rect 294506 316004 294512 316016
rect 294564 316004 294570 316056
rect 294598 316004 294604 316056
rect 294656 316044 294662 316056
rect 301038 316044 301044 316056
rect 294656 316016 301044 316044
rect 294656 316004 294662 316016
rect 301038 316004 301044 316016
rect 301096 316004 301102 316056
rect 303890 316004 303896 316056
rect 303948 316044 303954 316056
rect 304810 316044 304816 316056
rect 303948 316016 304816 316044
rect 303948 316004 303954 316016
rect 304810 316004 304816 316016
rect 304868 316004 304874 316056
rect 306558 316004 306564 316056
rect 306616 316004 306622 316056
rect 306834 316004 306840 316056
rect 306892 316044 306898 316056
rect 307662 316044 307668 316056
rect 306892 316016 307668 316044
rect 306892 316004 306898 316016
rect 307662 316004 307668 316016
rect 307720 316004 307726 316056
rect 310790 316004 310796 316056
rect 310848 316044 310854 316056
rect 311158 316044 311164 316056
rect 310848 316016 311164 316044
rect 310848 316004 310854 316016
rect 311158 316004 311164 316016
rect 311216 316004 311222 316056
rect 318794 316004 318800 316056
rect 318852 316044 318858 316056
rect 319438 316044 319444 316056
rect 318852 316016 319444 316044
rect 318852 316004 318858 316016
rect 319438 316004 319444 316016
rect 319496 316004 319502 316056
rect 320174 316004 320180 316056
rect 320232 316044 320238 316056
rect 320634 316044 320640 316056
rect 320232 316016 320640 316044
rect 320232 316004 320238 316016
rect 320634 316004 320640 316016
rect 320692 316004 320698 316056
rect 321646 316004 321652 316056
rect 321704 316044 321710 316056
rect 322474 316044 322480 316056
rect 321704 316016 322480 316044
rect 321704 316004 321710 316016
rect 322474 316004 322480 316016
rect 322532 316004 322538 316056
rect 322842 316004 322848 316056
rect 322900 316044 322906 316056
rect 327442 316044 327448 316056
rect 322900 316016 327448 316044
rect 322900 316004 322906 316016
rect 327442 316004 327448 316016
rect 327500 316004 327506 316056
rect 327902 316004 327908 316056
rect 327960 316044 327966 316056
rect 554038 316044 554044 316056
rect 327960 316016 554044 316044
rect 327960 316004 327966 316016
rect 554038 316004 554044 316016
rect 554096 316004 554102 316056
rect 292850 315936 292856 315988
rect 292908 315976 292914 315988
rect 293770 315976 293776 315988
rect 292908 315948 293776 315976
rect 292908 315936 292914 315948
rect 293770 315936 293776 315948
rect 293828 315936 293834 315988
rect 299750 315936 299756 315988
rect 299808 315976 299814 315988
rect 300486 315976 300492 315988
rect 299808 315948 300492 315976
rect 299808 315936 299814 315948
rect 300486 315936 300492 315948
rect 300544 315936 300550 315988
rect 302510 315936 302516 315988
rect 302568 315976 302574 315988
rect 303154 315976 303160 315988
rect 302568 315948 303160 315976
rect 302568 315936 302574 315948
rect 303154 315936 303160 315948
rect 303212 315936 303218 315988
rect 303798 315936 303804 315988
rect 303856 315976 303862 315988
rect 304626 315976 304632 315988
rect 303856 315948 304632 315976
rect 303856 315936 303862 315948
rect 304626 315936 304632 315948
rect 304684 315936 304690 315988
rect 306374 315936 306380 315988
rect 306432 315976 306438 315988
rect 306576 315976 306604 316004
rect 306432 315948 306604 315976
rect 306432 315936 306438 315948
rect 306650 315936 306656 315988
rect 306708 315976 306714 315988
rect 307386 315976 307392 315988
rect 306708 315948 307392 315976
rect 306708 315936 306714 315948
rect 307386 315936 307392 315948
rect 307444 315936 307450 315988
rect 308398 315936 308404 315988
rect 308456 315976 308462 315988
rect 308858 315976 308864 315988
rect 308456 315948 308864 315976
rect 308456 315936 308462 315948
rect 308858 315936 308864 315948
rect 308916 315936 308922 315988
rect 310514 315936 310520 315988
rect 310572 315976 310578 315988
rect 311526 315976 311532 315988
rect 310572 315948 311532 315976
rect 310572 315936 310578 315948
rect 311526 315936 311532 315948
rect 311584 315936 311590 315988
rect 312078 315936 312084 315988
rect 312136 315976 312142 315988
rect 312446 315976 312452 315988
rect 312136 315948 312452 315976
rect 312136 315936 312142 315948
rect 312446 315936 312452 315948
rect 312504 315936 312510 315988
rect 312722 315936 312728 315988
rect 312780 315976 312786 315988
rect 312998 315976 313004 315988
rect 312780 315948 313004 315976
rect 312780 315936 312786 315948
rect 312998 315936 313004 315948
rect 313056 315936 313062 315988
rect 313642 315936 313648 315988
rect 313700 315976 313706 315988
rect 314286 315976 314292 315988
rect 313700 315948 314292 315976
rect 313700 315936 313706 315948
rect 314286 315936 314292 315948
rect 314344 315936 314350 315988
rect 315390 315936 315396 315988
rect 315448 315976 315454 315988
rect 315758 315976 315764 315988
rect 315448 315948 315764 315976
rect 315448 315936 315454 315948
rect 315758 315936 315764 315948
rect 315816 315936 315822 315988
rect 319162 315936 319168 315988
rect 319220 315976 319226 315988
rect 319714 315976 319720 315988
rect 319220 315948 319720 315976
rect 319220 315936 319226 315948
rect 319714 315936 319720 315948
rect 319772 315936 319778 315988
rect 320450 315936 320456 315988
rect 320508 315976 320514 315988
rect 321002 315976 321008 315988
rect 320508 315948 321008 315976
rect 320508 315936 320514 315948
rect 321002 315936 321008 315948
rect 321060 315936 321066 315988
rect 321554 315936 321560 315988
rect 321612 315976 321618 315988
rect 322750 315976 322756 315988
rect 321612 315948 322756 315976
rect 321612 315936 321618 315948
rect 322750 315936 322756 315948
rect 322808 315936 322814 315988
rect 324682 315936 324688 315988
rect 324740 315976 324746 315988
rect 324866 315976 324872 315988
rect 324740 315948 324872 315976
rect 324740 315936 324746 315948
rect 324866 315936 324872 315948
rect 324924 315936 324930 315988
rect 325786 315936 325792 315988
rect 325844 315976 325850 315988
rect 326246 315976 326252 315988
rect 325844 315948 326252 315976
rect 325844 315936 325850 315948
rect 326246 315936 326252 315948
rect 326304 315936 326310 315988
rect 327074 315936 327080 315988
rect 327132 315976 327138 315988
rect 327258 315976 327264 315988
rect 327132 315948 327264 315976
rect 327132 315936 327138 315948
rect 327258 315936 327264 315948
rect 327316 315936 327322 315988
rect 276808 315880 292436 315908
rect 276808 315868 276814 315880
rect 306558 315868 306564 315920
rect 306616 315908 306622 315920
rect 307294 315908 307300 315920
rect 306616 315880 307300 315908
rect 306616 315868 306622 315880
rect 307294 315868 307300 315880
rect 307352 315868 307358 315920
rect 308122 315868 308128 315920
rect 308180 315908 308186 315920
rect 308766 315908 308772 315920
rect 308180 315880 308772 315908
rect 308180 315868 308186 315880
rect 308766 315868 308772 315880
rect 308824 315868 308830 315920
rect 309318 315868 309324 315920
rect 309376 315908 309382 315920
rect 310330 315908 310336 315920
rect 309376 315880 310336 315908
rect 309376 315868 309382 315880
rect 310330 315868 310336 315880
rect 310388 315868 310394 315920
rect 321738 315868 321744 315920
rect 321796 315908 321802 315920
rect 321922 315908 321928 315920
rect 321796 315880 321928 315908
rect 321796 315868 321802 315880
rect 321922 315868 321928 315880
rect 321980 315868 321986 315920
rect 323302 315868 323308 315920
rect 323360 315908 323366 315920
rect 323946 315908 323952 315920
rect 323360 315880 323952 315908
rect 323360 315868 323366 315880
rect 323946 315868 323952 315880
rect 324004 315868 324010 315920
rect 274358 315800 274364 315852
rect 274416 315840 274422 315852
rect 274416 315812 292712 315840
rect 274416 315800 274422 315812
rect 272702 315732 272708 315784
rect 272760 315772 272766 315784
rect 292574 315772 292580 315784
rect 272760 315744 292580 315772
rect 272760 315732 272766 315744
rect 292574 315732 292580 315744
rect 292632 315732 292638 315784
rect 292684 315772 292712 315812
rect 292758 315800 292764 315852
rect 292816 315840 292822 315852
rect 293218 315840 293224 315852
rect 292816 315812 293224 315840
rect 292816 315800 292822 315812
rect 293218 315800 293224 315812
rect 293276 315800 293282 315852
rect 294414 315800 294420 315852
rect 294472 315840 294478 315852
rect 294874 315840 294880 315852
rect 294472 315812 294880 315840
rect 294472 315800 294478 315812
rect 294874 315800 294880 315812
rect 294932 315800 294938 315852
rect 306190 315800 306196 315852
rect 306248 315840 306254 315852
rect 307938 315840 307944 315852
rect 306248 315812 307944 315840
rect 306248 315800 306254 315812
rect 307938 315800 307944 315812
rect 307996 315800 308002 315852
rect 312446 315800 312452 315852
rect 312504 315840 312510 315852
rect 312722 315840 312728 315852
rect 312504 315812 312728 315840
rect 312504 315800 312510 315812
rect 312722 315800 312728 315812
rect 312780 315800 312786 315852
rect 313458 315800 313464 315852
rect 313516 315840 313522 315852
rect 314102 315840 314108 315852
rect 313516 315812 314108 315840
rect 313516 315800 313522 315812
rect 314102 315800 314108 315812
rect 314160 315800 314166 315852
rect 315206 315800 315212 315852
rect 315264 315840 315270 315852
rect 315574 315840 315580 315852
rect 315264 315812 315580 315840
rect 315264 315800 315270 315812
rect 315574 315800 315580 315812
rect 315632 315800 315638 315852
rect 320542 315800 320548 315852
rect 320600 315840 320606 315852
rect 321186 315840 321192 315852
rect 320600 315812 321192 315840
rect 320600 315800 320606 315812
rect 321186 315800 321192 315812
rect 321244 315800 321250 315852
rect 294046 315772 294052 315784
rect 292684 315744 294052 315772
rect 294046 315732 294052 315744
rect 294104 315732 294110 315784
rect 294322 315732 294328 315784
rect 294380 315772 294386 315784
rect 294690 315772 294696 315784
rect 294380 315744 294696 315772
rect 294380 315732 294386 315744
rect 294690 315732 294696 315744
rect 294748 315732 294754 315784
rect 307018 315732 307024 315784
rect 307076 315772 307082 315784
rect 309410 315772 309416 315784
rect 307076 315744 309416 315772
rect 307076 315732 307082 315744
rect 309410 315732 309416 315744
rect 309468 315732 309474 315784
rect 312354 315732 312360 315784
rect 312412 315772 312418 315784
rect 313182 315772 313188 315784
rect 312412 315744 313188 315772
rect 312412 315732 312418 315744
rect 313182 315732 313188 315744
rect 313240 315732 313246 315784
rect 274082 315664 274088 315716
rect 274140 315704 274146 315716
rect 292390 315704 292396 315716
rect 274140 315676 292396 315704
rect 274140 315664 274146 315676
rect 292390 315664 292396 315676
rect 292448 315664 292454 315716
rect 293034 315664 293040 315716
rect 293092 315704 293098 315716
rect 301682 315704 301688 315716
rect 293092 315676 301688 315704
rect 293092 315664 293098 315676
rect 301682 315664 301688 315676
rect 301740 315664 301746 315716
rect 306374 315664 306380 315716
rect 306432 315704 306438 315716
rect 310882 315704 310888 315716
rect 306432 315676 310888 315704
rect 306432 315664 306438 315676
rect 310882 315664 310888 315676
rect 310940 315664 310946 315716
rect 317782 315704 317788 315716
rect 311866 315676 317788 315704
rect 271230 315596 271236 315648
rect 271288 315636 271294 315648
rect 292298 315636 292304 315648
rect 271288 315608 292304 315636
rect 271288 315596 271294 315608
rect 292298 315596 292304 315608
rect 292356 315596 292362 315648
rect 294690 315596 294696 315648
rect 294748 315636 294754 315648
rect 303522 315636 303528 315648
rect 294748 315608 303528 315636
rect 294748 315596 294754 315608
rect 303522 315596 303528 315608
rect 303580 315596 303586 315648
rect 307662 315596 307668 315648
rect 307720 315636 307726 315648
rect 311866 315636 311894 315676
rect 317782 315664 317788 315676
rect 317840 315664 317846 315716
rect 307720 315608 311894 315636
rect 307720 315596 307726 315608
rect 311986 315596 311992 315648
rect 312044 315636 312050 315648
rect 313182 315636 313188 315648
rect 312044 315608 313188 315636
rect 312044 315596 312050 315608
rect 313182 315596 313188 315608
rect 313240 315596 313246 315648
rect 268378 315528 268384 315580
rect 268436 315568 268442 315580
rect 293954 315568 293960 315580
rect 268436 315540 293960 315568
rect 268436 315528 268442 315540
rect 293954 315528 293960 315540
rect 294012 315528 294018 315580
rect 294046 315528 294052 315580
rect 294104 315568 294110 315580
rect 299934 315568 299940 315580
rect 294104 315540 299940 315568
rect 294104 315528 294110 315540
rect 299934 315528 299940 315540
rect 299992 315528 299998 315580
rect 302878 315528 302884 315580
rect 302936 315568 302942 315580
rect 314838 315568 314844 315580
rect 302936 315540 314844 315568
rect 302936 315528 302942 315540
rect 314838 315528 314844 315540
rect 314896 315528 314902 315580
rect 272518 315460 272524 315512
rect 272576 315500 272582 315512
rect 316770 315500 316776 315512
rect 272576 315472 292528 315500
rect 272576 315460 272582 315472
rect 233050 315392 233056 315444
rect 233108 315432 233114 315444
rect 282914 315432 282920 315444
rect 233108 315404 282920 315432
rect 233108 315392 233114 315404
rect 282914 315392 282920 315404
rect 282972 315392 282978 315444
rect 283558 315392 283564 315444
rect 283616 315432 283622 315444
rect 284386 315432 284392 315444
rect 283616 315404 284392 315432
rect 283616 315392 283622 315404
rect 284386 315392 284392 315404
rect 284444 315392 284450 315444
rect 287606 315392 287612 315444
rect 287664 315432 287670 315444
rect 288250 315432 288256 315444
rect 287664 315404 288256 315432
rect 287664 315392 287670 315404
rect 288250 315392 288256 315404
rect 288308 315392 288314 315444
rect 289998 315392 290004 315444
rect 290056 315432 290062 315444
rect 290366 315432 290372 315444
rect 290056 315404 290372 315432
rect 290056 315392 290062 315404
rect 290366 315392 290372 315404
rect 290424 315392 290430 315444
rect 292500 315432 292528 315472
rect 292776 315472 316776 315500
rect 292776 315432 292804 315472
rect 316770 315460 316776 315472
rect 316828 315460 316834 315512
rect 292500 315404 292804 315432
rect 293954 315392 293960 315444
rect 294012 315432 294018 315444
rect 302050 315432 302056 315444
rect 294012 315404 302056 315432
rect 294012 315392 294018 315404
rect 302050 315392 302056 315404
rect 302108 315392 302114 315444
rect 308490 315392 308496 315444
rect 308548 315432 308554 315444
rect 331306 315432 331312 315444
rect 308548 315404 331312 315432
rect 308548 315392 308554 315404
rect 331306 315392 331312 315404
rect 331364 315392 331370 315444
rect 217686 315324 217692 315376
rect 217744 315364 217750 315376
rect 280154 315364 280160 315376
rect 217744 315336 280160 315364
rect 217744 315324 217750 315336
rect 280154 315324 280160 315336
rect 280212 315324 280218 315376
rect 287698 315324 287704 315376
rect 287756 315364 287762 315376
rect 287974 315364 287980 315376
rect 287756 315336 287980 315364
rect 287756 315324 287762 315336
rect 287974 315324 287980 315336
rect 288032 315324 288038 315376
rect 288342 315324 288348 315376
rect 288400 315364 288406 315376
rect 290274 315364 290280 315376
rect 288400 315336 290280 315364
rect 288400 315324 288406 315336
rect 290274 315324 290280 315336
rect 290332 315324 290338 315376
rect 292298 315324 292304 315376
rect 292356 315364 292362 315376
rect 294690 315364 294696 315376
rect 292356 315336 294696 315364
rect 292356 315324 292362 315336
rect 294690 315324 294696 315336
rect 294748 315324 294754 315376
rect 309962 315324 309968 315376
rect 310020 315364 310026 315376
rect 335998 315364 336004 315376
rect 310020 315336 336004 315364
rect 310020 315324 310026 315336
rect 335998 315324 336004 315336
rect 336056 315324 336062 315376
rect 215018 315256 215024 315308
rect 215076 315296 215082 315308
rect 284294 315296 284300 315308
rect 215076 315268 284300 315296
rect 215076 315256 215082 315268
rect 284294 315256 284300 315268
rect 284352 315256 284358 315308
rect 284386 315256 284392 315308
rect 284444 315296 284450 315308
rect 285030 315296 285036 315308
rect 284444 315268 285036 315296
rect 284444 315256 284450 315268
rect 285030 315256 285036 315268
rect 285088 315256 285094 315308
rect 287146 315256 287152 315308
rect 287204 315296 287210 315308
rect 288250 315296 288256 315308
rect 287204 315268 288256 315296
rect 287204 315256 287210 315268
rect 288250 315256 288256 315268
rect 288308 315256 288314 315308
rect 288434 315256 288440 315308
rect 288492 315296 288498 315308
rect 289538 315296 289544 315308
rect 288492 315268 289544 315296
rect 288492 315256 288498 315268
rect 289538 315256 289544 315268
rect 289596 315256 289602 315308
rect 291838 315256 291844 315308
rect 291896 315296 291902 315308
rect 306098 315296 306104 315308
rect 291896 315268 306104 315296
rect 291896 315256 291902 315268
rect 306098 315256 306104 315268
rect 306156 315256 306162 315308
rect 367094 315296 367100 315308
rect 311866 315268 367100 315296
rect 279694 315188 279700 315240
rect 279752 315228 279758 315240
rect 300670 315228 300676 315240
rect 279752 315200 300676 315228
rect 279752 315188 279758 315200
rect 300670 315188 300676 315200
rect 300728 315188 300734 315240
rect 303154 315188 303160 315240
rect 303212 315228 303218 315240
rect 311066 315228 311072 315240
rect 303212 315200 311072 315228
rect 303212 315188 303218 315200
rect 311066 315188 311072 315200
rect 311124 315228 311130 315240
rect 311866 315228 311894 315268
rect 367094 315256 367100 315268
rect 367152 315256 367158 315308
rect 311124 315200 311894 315228
rect 311124 315188 311130 315200
rect 278682 315120 278688 315172
rect 278740 315160 278746 315172
rect 295150 315160 295156 315172
rect 278740 315132 295156 315160
rect 278740 315120 278746 315132
rect 295150 315120 295156 315132
rect 295208 315120 295214 315172
rect 282914 315052 282920 315104
rect 282972 315092 282978 315104
rect 288894 315092 288900 315104
rect 282972 315064 288900 315092
rect 282972 315052 282978 315064
rect 288894 315052 288900 315064
rect 288952 315052 288958 315104
rect 292574 315052 292580 315104
rect 292632 315092 292638 315104
rect 299382 315092 299388 315104
rect 292632 315064 299388 315092
rect 292632 315052 292638 315064
rect 299382 315052 299388 315064
rect 299440 315052 299446 315104
rect 286410 314984 286416 315036
rect 286468 315024 286474 315036
rect 287882 315024 287888 315036
rect 286468 314996 287888 315024
rect 286468 314984 286474 314996
rect 287882 314984 287888 314996
rect 287940 314984 287946 315036
rect 312630 314712 312636 314764
rect 312688 314752 312694 314764
rect 396074 314752 396080 314764
rect 312688 314724 396080 314752
rect 312688 314712 312694 314724
rect 396074 314712 396080 314724
rect 396132 314712 396138 314764
rect 313918 314644 313924 314696
rect 313976 314684 313982 314696
rect 407114 314684 407120 314696
rect 313976 314656 407120 314684
rect 313976 314644 313982 314656
rect 407114 314644 407120 314656
rect 407172 314644 407178 314696
rect 276658 314576 276664 314628
rect 276716 314616 276722 314628
rect 290550 314616 290556 314628
rect 276716 314588 290556 314616
rect 276716 314576 276722 314588
rect 290550 314576 290556 314588
rect 290608 314576 290614 314628
rect 269850 314508 269856 314560
rect 269908 314548 269914 314560
rect 290458 314548 290464 314560
rect 269908 314520 290464 314548
rect 269908 314508 269914 314520
rect 290458 314508 290464 314520
rect 290516 314508 290522 314560
rect 299106 314508 299112 314560
rect 299164 314548 299170 314560
rect 299290 314548 299296 314560
rect 299164 314520 299296 314548
rect 299164 314508 299170 314520
rect 299290 314508 299296 314520
rect 299348 314508 299354 314560
rect 274542 314440 274548 314492
rect 274600 314480 274606 314492
rect 295242 314480 295248 314492
rect 274600 314452 295248 314480
rect 274600 314440 274606 314452
rect 295242 314440 295248 314452
rect 295300 314440 295306 314492
rect 279418 314372 279424 314424
rect 279476 314412 279482 314424
rect 304258 314412 304264 314424
rect 279476 314384 304264 314412
rect 279476 314372 279482 314384
rect 304258 314372 304264 314384
rect 304316 314372 304322 314424
rect 320910 314372 320916 314424
rect 320968 314412 320974 314424
rect 328914 314412 328920 314424
rect 320968 314384 328920 314412
rect 320968 314372 320974 314384
rect 328914 314372 328920 314384
rect 328972 314372 328978 314424
rect 280890 314304 280896 314356
rect 280948 314344 280954 314356
rect 315942 314344 315948 314356
rect 280948 314316 315948 314344
rect 280948 314304 280954 314316
rect 315942 314304 315948 314316
rect 316000 314344 316006 314356
rect 316000 314316 319392 314344
rect 316000 314304 316006 314316
rect 270034 314236 270040 314288
rect 270092 314276 270098 314288
rect 319254 314276 319260 314288
rect 270092 314248 319260 314276
rect 270092 314236 270098 314248
rect 319254 314236 319260 314248
rect 319312 314236 319318 314288
rect 286870 314168 286876 314220
rect 286928 314208 286934 314220
rect 298738 314208 298744 314220
rect 286928 314180 298744 314208
rect 286928 314168 286934 314180
rect 298738 314168 298744 314180
rect 298796 314168 298802 314220
rect 220538 314100 220544 314152
rect 220596 314140 220602 314152
rect 292206 314140 292212 314152
rect 220596 314112 292212 314140
rect 220596 314100 220602 314112
rect 292206 314100 292212 314112
rect 292264 314100 292270 314152
rect 218882 314032 218888 314084
rect 218940 314072 218946 314084
rect 291930 314072 291936 314084
rect 218940 314044 291936 314072
rect 218940 314032 218946 314044
rect 291930 314032 291936 314044
rect 291988 314032 291994 314084
rect 216306 313964 216312 314016
rect 216364 314004 216370 314016
rect 297818 314004 297824 314016
rect 216364 313976 297824 314004
rect 216364 313964 216370 313976
rect 297818 313964 297824 313976
rect 297876 313964 297882 314016
rect 319364 314004 319392 314316
rect 319622 314032 319628 314084
rect 319680 314072 319686 314084
rect 330294 314072 330300 314084
rect 319680 314044 330300 314072
rect 319680 314032 319686 314044
rect 330294 314032 330300 314044
rect 330352 314032 330358 314084
rect 431954 314004 431960 314016
rect 319364 313976 431960 314004
rect 431954 313964 431960 313976
rect 432012 313964 432018 314016
rect 216398 313896 216404 313948
rect 216456 313936 216462 313948
rect 216456 313908 287744 313936
rect 216456 313896 216462 313908
rect 221826 313828 221832 313880
rect 221884 313868 221890 313880
rect 286686 313868 286692 313880
rect 221884 313840 286692 313868
rect 221884 313828 221890 313840
rect 286686 313828 286692 313840
rect 286744 313828 286750 313880
rect 287716 313800 287744 313908
rect 291654 313896 291660 313948
rect 291712 313936 291718 313948
rect 292482 313936 292488 313948
rect 291712 313908 292488 313936
rect 291712 313896 291718 313908
rect 292482 313896 292488 313908
rect 292540 313896 292546 313948
rect 316954 313896 316960 313948
rect 317012 313936 317018 313948
rect 441614 313936 441620 313948
rect 317012 313908 441620 313936
rect 317012 313896 317018 313908
rect 441614 313896 441620 313908
rect 441672 313896 441678 313948
rect 297726 313800 297732 313812
rect 287716 313772 297732 313800
rect 297726 313760 297732 313772
rect 297784 313760 297790 313812
rect 315482 313760 315488 313812
rect 315540 313800 315546 313812
rect 316954 313800 316960 313812
rect 315540 313772 316960 313800
rect 315540 313760 315546 313772
rect 316954 313760 316960 313772
rect 317012 313760 317018 313812
rect 290642 313624 290648 313676
rect 290700 313664 290706 313676
rect 291194 313664 291200 313676
rect 290700 313636 291200 313664
rect 290700 313624 290706 313636
rect 291194 313624 291200 313636
rect 291252 313624 291258 313676
rect 300118 313352 300124 313404
rect 300176 313392 300182 313404
rect 306006 313392 306012 313404
rect 300176 313364 306012 313392
rect 300176 313352 300182 313364
rect 306006 313352 306012 313364
rect 306064 313352 306070 313404
rect 315298 313352 315304 313404
rect 315356 313392 315362 313404
rect 422938 313392 422944 313404
rect 315356 313364 422944 313392
rect 315356 313352 315362 313364
rect 422938 313352 422944 313364
rect 422996 313352 423002 313404
rect 268562 313284 268568 313336
rect 268620 313324 268626 313336
rect 314102 313324 314108 313336
rect 268620 313296 314108 313324
rect 268620 313284 268626 313296
rect 314102 313284 314108 313296
rect 314160 313284 314166 313336
rect 315390 313284 315396 313336
rect 315448 313324 315454 313336
rect 427814 313324 427820 313336
rect 315448 313296 427820 313324
rect 315448 313284 315454 313296
rect 427814 313284 427820 313296
rect 427872 313284 427878 313336
rect 293218 313216 293224 313268
rect 293276 313256 293282 313268
rect 296530 313256 296536 313268
rect 293276 313228 296536 313256
rect 293276 313216 293282 313228
rect 296530 313216 296536 313228
rect 296588 313216 296594 313268
rect 313274 313216 313280 313268
rect 313332 313256 313338 313268
rect 313826 313256 313832 313268
rect 313332 313228 313832 313256
rect 313332 313216 313338 313228
rect 313826 313216 313832 313228
rect 313884 313216 313890 313268
rect 296162 313148 296168 313200
rect 296220 313188 296226 313200
rect 300026 313188 300032 313200
rect 296220 313160 300032 313188
rect 296220 313148 296226 313160
rect 300026 313148 300032 313160
rect 300084 313148 300090 313200
rect 271690 313080 271696 313132
rect 271748 313120 271754 313132
rect 304534 313120 304540 313132
rect 271748 313092 304540 313120
rect 271748 313080 271754 313092
rect 304534 313080 304540 313092
rect 304592 313080 304598 313132
rect 278406 313012 278412 313064
rect 278464 313052 278470 313064
rect 312814 313052 312820 313064
rect 278464 313024 312820 313052
rect 278464 313012 278470 313024
rect 312814 313012 312820 313024
rect 312872 313012 312878 313064
rect 275370 312944 275376 312996
rect 275428 312984 275434 312996
rect 318058 312984 318064 312996
rect 275428 312956 318064 312984
rect 275428 312944 275434 312956
rect 318058 312944 318064 312956
rect 318116 312944 318122 312996
rect 252462 312876 252468 312928
rect 252520 312916 252526 312928
rect 311342 312916 311348 312928
rect 252520 312888 311348 312916
rect 252520 312876 252526 312888
rect 311342 312876 311348 312888
rect 311400 312876 311406 312928
rect 235626 312808 235632 312860
rect 235684 312848 235690 312860
rect 296438 312848 296444 312860
rect 235684 312820 296444 312848
rect 235684 312808 235690 312820
rect 296438 312808 296444 312820
rect 296496 312808 296502 312860
rect 297450 312808 297456 312860
rect 297508 312848 297514 312860
rect 321094 312848 321100 312860
rect 297508 312820 321100 312848
rect 297508 312808 297514 312820
rect 321094 312808 321100 312820
rect 321152 312808 321158 312860
rect 235902 312740 235908 312792
rect 235960 312780 235966 312792
rect 295886 312780 295892 312792
rect 235960 312752 295892 312780
rect 235960 312740 235966 312752
rect 295886 312740 295892 312752
rect 295944 312740 295950 312792
rect 309686 312740 309692 312792
rect 309744 312780 309750 312792
rect 342254 312780 342260 312792
rect 309744 312752 342260 312780
rect 309744 312740 309750 312752
rect 342254 312740 342260 312752
rect 342312 312740 342318 312792
rect 216030 312672 216036 312724
rect 216088 312712 216094 312724
rect 282546 312712 282552 312724
rect 216088 312684 282552 312712
rect 216088 312672 216094 312684
rect 282546 312672 282552 312684
rect 282604 312672 282610 312724
rect 315022 312712 315028 312724
rect 292546 312684 315028 312712
rect 216122 312604 216128 312656
rect 216180 312644 216186 312656
rect 284018 312644 284024 312656
rect 216180 312616 284024 312644
rect 216180 312604 216186 312616
rect 284018 312604 284024 312616
rect 284076 312604 284082 312656
rect 215938 312536 215944 312588
rect 215996 312576 216002 312588
rect 215996 312548 273254 312576
rect 215996 312536 216002 312548
rect 273226 312508 273254 312548
rect 282546 312536 282552 312588
rect 282604 312576 282610 312588
rect 292546 312576 292574 312684
rect 315022 312672 315028 312684
rect 315080 312672 315086 312724
rect 321094 312672 321100 312724
rect 321152 312712 321158 312724
rect 500218 312712 500224 312724
rect 321152 312684 500224 312712
rect 321152 312672 321158 312684
rect 500218 312672 500224 312684
rect 500276 312672 500282 312724
rect 322290 312604 322296 312656
rect 322348 312644 322354 312656
rect 511258 312644 511264 312656
rect 322348 312616 511264 312644
rect 322348 312604 322354 312616
rect 511258 312604 511264 312616
rect 511316 312604 511322 312656
rect 282604 312548 292574 312576
rect 282604 312536 282610 312548
rect 320910 312536 320916 312588
rect 320968 312576 320974 312588
rect 323026 312576 323032 312588
rect 320968 312548 323032 312576
rect 320968 312536 320974 312548
rect 323026 312536 323032 312548
rect 323084 312576 323090 312588
rect 526438 312576 526444 312588
rect 323084 312548 526444 312576
rect 323084 312536 323090 312548
rect 526438 312536 526444 312548
rect 526496 312536 526502 312588
rect 286502 312508 286508 312520
rect 273226 312480 286508 312508
rect 286502 312468 286508 312480
rect 286560 312468 286566 312520
rect 302970 312060 302976 312112
rect 303028 312100 303034 312112
rect 303154 312100 303160 312112
rect 303028 312072 303160 312100
rect 303028 312060 303034 312072
rect 303154 312060 303160 312072
rect 303212 312060 303218 312112
rect 288434 312032 288440 312044
rect 273226 312004 288440 312032
rect 213822 311924 213828 311976
rect 213880 311964 213886 311976
rect 273226 311964 273254 312004
rect 288434 311992 288440 312004
rect 288492 311992 288498 312044
rect 292574 311964 292580 311976
rect 213880 311936 273254 311964
rect 287716 311936 292580 311964
rect 213880 311924 213886 311936
rect 217502 311856 217508 311908
rect 217560 311896 217566 311908
rect 287716 311896 287744 311936
rect 292574 311924 292580 311936
rect 292632 311924 292638 311976
rect 320818 311924 320824 311976
rect 320876 311964 320882 311976
rect 322290 311964 322296 311976
rect 320876 311936 322296 311964
rect 320876 311924 320882 311936
rect 322290 311924 322296 311936
rect 322348 311924 322354 311976
rect 217560 311868 287744 311896
rect 217560 311856 217566 311868
rect 291930 311856 291936 311908
rect 291988 311896 291994 311908
rect 293586 311896 293592 311908
rect 291988 311868 293592 311896
rect 291988 311856 291994 311868
rect 293586 311856 293592 311868
rect 293644 311856 293650 311908
rect 313274 311856 313280 311908
rect 313332 311896 313338 311908
rect 409874 311896 409880 311908
rect 313332 311868 409880 311896
rect 313332 311856 313338 311868
rect 409874 311856 409880 311868
rect 409932 311856 409938 311908
rect 279510 311584 279516 311636
rect 279568 311624 279574 311636
rect 288250 311624 288256 311636
rect 279568 311596 288256 311624
rect 279568 311584 279574 311596
rect 288250 311584 288256 311596
rect 288308 311584 288314 311636
rect 277210 311516 277216 311568
rect 277268 311556 277274 311568
rect 303062 311556 303068 311568
rect 277268 311528 303068 311556
rect 277268 311516 277274 311528
rect 303062 311516 303068 311528
rect 303120 311516 303126 311568
rect 224586 311448 224592 311500
rect 224644 311488 224650 311500
rect 283006 311488 283012 311500
rect 224644 311460 283012 311488
rect 224644 311448 224650 311460
rect 283006 311448 283012 311460
rect 283064 311448 283070 311500
rect 300118 311448 300124 311500
rect 300176 311488 300182 311500
rect 300302 311488 300308 311500
rect 300176 311460 300308 311488
rect 300176 311448 300182 311460
rect 300302 311448 300308 311460
rect 300360 311448 300366 311500
rect 251082 311380 251088 311432
rect 251140 311420 251146 311432
rect 309502 311420 309508 311432
rect 251140 311392 309508 311420
rect 251140 311380 251146 311392
rect 309502 311380 309508 311392
rect 309560 311380 309566 311432
rect 249610 311312 249616 311364
rect 249668 311352 249674 311364
rect 309226 311352 309232 311364
rect 249668 311324 309232 311352
rect 249668 311312 249674 311324
rect 309226 311312 309232 311324
rect 309284 311312 309290 311364
rect 250990 311244 250996 311296
rect 251048 311284 251054 311296
rect 310606 311284 310612 311296
rect 251048 311256 310612 311284
rect 251048 311244 251054 311256
rect 310606 311244 310612 311256
rect 310664 311244 310670 311296
rect 250714 311176 250720 311228
rect 250772 311216 250778 311228
rect 311526 311216 311532 311228
rect 250772 311188 311532 311216
rect 250772 311176 250778 311188
rect 311526 311176 311532 311188
rect 311584 311176 311590 311228
rect 221642 311108 221648 311160
rect 221700 311148 221706 311160
rect 221700 311120 277394 311148
rect 221700 311108 221706 311120
rect 277366 311080 277394 311120
rect 280982 311108 280988 311160
rect 281040 311148 281046 311160
rect 281258 311148 281264 311160
rect 281040 311120 281264 311148
rect 281040 311108 281046 311120
rect 281258 311108 281264 311120
rect 281316 311108 281322 311160
rect 282638 311108 282644 311160
rect 282696 311148 282702 311160
rect 289446 311148 289452 311160
rect 282696 311120 289452 311148
rect 282696 311108 282702 311120
rect 289446 311108 289452 311120
rect 289504 311108 289510 311160
rect 294598 311108 294604 311160
rect 294656 311148 294662 311160
rect 294782 311148 294788 311160
rect 294656 311120 294788 311148
rect 294656 311108 294662 311120
rect 294782 311108 294788 311120
rect 294840 311108 294846 311160
rect 298738 311108 298744 311160
rect 298796 311148 298802 311160
rect 299106 311148 299112 311160
rect 298796 311120 299112 311148
rect 298796 311108 298802 311120
rect 299106 311108 299112 311120
rect 299164 311108 299170 311160
rect 300946 311108 300952 311160
rect 301004 311148 301010 311160
rect 301958 311148 301964 311160
rect 301004 311120 301964 311148
rect 301004 311108 301010 311120
rect 301958 311108 301964 311120
rect 302016 311108 302022 311160
rect 314102 311108 314108 311160
rect 314160 311148 314166 311160
rect 414014 311148 414020 311160
rect 314160 311120 414020 311148
rect 314160 311108 314166 311120
rect 414014 311108 414020 311120
rect 414072 311108 414078 311160
rect 284662 311080 284668 311092
rect 277366 311052 284668 311080
rect 284662 311040 284668 311052
rect 284720 311040 284726 311092
rect 312354 310564 312360 310616
rect 312412 310604 312418 310616
rect 312630 310604 312636 310616
rect 312412 310576 312636 310604
rect 312412 310564 312418 310576
rect 312630 310564 312636 310576
rect 312688 310604 312694 310616
rect 391934 310604 391940 310616
rect 312688 310576 391940 310604
rect 312688 310564 312694 310576
rect 391934 310564 391940 310576
rect 391992 310564 391998 310616
rect 324406 310496 324412 310548
rect 324464 310536 324470 310548
rect 324774 310536 324780 310548
rect 324464 310508 324780 310536
rect 324464 310496 324470 310508
rect 324774 310496 324780 310508
rect 324832 310536 324838 310548
rect 542998 310536 543004 310548
rect 324832 310508 543004 310536
rect 324832 310496 324838 310508
rect 542998 310496 543004 310508
rect 543056 310496 543062 310548
rect 289170 310428 289176 310480
rect 289228 310468 289234 310480
rect 293310 310468 293316 310480
rect 289228 310440 293316 310468
rect 289228 310428 289234 310440
rect 293310 310428 293316 310440
rect 293368 310428 293374 310480
rect 289262 310360 289268 310412
rect 289320 310400 289326 310412
rect 295334 310400 295340 310412
rect 289320 310372 295340 310400
rect 289320 310360 289326 310372
rect 295334 310360 295340 310372
rect 295392 310360 295398 310412
rect 276014 310292 276020 310344
rect 276072 310332 276078 310344
rect 285674 310332 285680 310344
rect 276072 310304 285680 310332
rect 276072 310292 276078 310304
rect 285674 310292 285680 310304
rect 285732 310292 285738 310344
rect 278222 310224 278228 310276
rect 278280 310264 278286 310276
rect 288618 310264 288624 310276
rect 278280 310236 288624 310264
rect 278280 310224 278286 310236
rect 288618 310224 288624 310236
rect 288676 310224 288682 310276
rect 256510 310156 256516 310208
rect 256568 310196 256574 310208
rect 314746 310196 314752 310208
rect 256568 310168 314752 310196
rect 256568 310156 256574 310168
rect 314746 310156 314752 310168
rect 314804 310156 314810 310208
rect 256602 310088 256608 310140
rect 256660 310128 256666 310140
rect 317230 310128 317236 310140
rect 256660 310100 317236 310128
rect 256660 310088 256666 310100
rect 317230 310088 317236 310100
rect 317288 310088 317294 310140
rect 256234 310020 256240 310072
rect 256292 310060 256298 310072
rect 316126 310060 316132 310072
rect 256292 310032 316132 310060
rect 256292 310020 256298 310032
rect 316126 310020 316132 310032
rect 316184 310020 316190 310072
rect 215754 309952 215760 310004
rect 215812 309992 215818 310004
rect 281718 309992 281724 310004
rect 215812 309964 281724 309992
rect 215812 309952 215818 309964
rect 281718 309952 281724 309964
rect 281776 309952 281782 310004
rect 285030 309952 285036 310004
rect 285088 309992 285094 310004
rect 318242 309992 318248 310004
rect 285088 309964 318248 309992
rect 285088 309952 285094 309964
rect 318242 309952 318248 309964
rect 318300 309952 318306 310004
rect 214926 309884 214932 309936
rect 214984 309924 214990 309936
rect 284386 309924 284392 309936
rect 214984 309896 284392 309924
rect 214984 309884 214990 309896
rect 284386 309884 284392 309896
rect 284444 309884 284450 309936
rect 286502 309884 286508 309936
rect 286560 309924 286566 309936
rect 318886 309924 318892 309936
rect 286560 309896 318892 309924
rect 286560 309884 286566 309896
rect 318886 309884 318892 309896
rect 318944 309884 318950 309936
rect 218606 309816 218612 309868
rect 218664 309856 218670 309868
rect 291102 309856 291108 309868
rect 218664 309828 291108 309856
rect 218664 309816 218670 309828
rect 291102 309816 291108 309828
rect 291160 309816 291166 309868
rect 214558 309748 214564 309800
rect 214616 309788 214622 309800
rect 290182 309788 290188 309800
rect 214616 309760 290188 309788
rect 214616 309748 214622 309760
rect 290182 309748 290188 309760
rect 290240 309748 290246 309800
rect 315574 309748 315580 309800
rect 315632 309788 315638 309800
rect 327350 309788 327356 309800
rect 315632 309760 327356 309788
rect 315632 309748 315638 309760
rect 327350 309748 327356 309760
rect 327408 309788 327414 309800
rect 565814 309788 565820 309800
rect 327408 309760 565820 309788
rect 327408 309748 327414 309760
rect 565814 309748 565820 309760
rect 565872 309748 565878 309800
rect 282270 309476 282276 309528
rect 282328 309516 282334 309528
rect 282546 309516 282552 309528
rect 282328 309488 282552 309516
rect 282328 309476 282334 309488
rect 282546 309476 282552 309488
rect 282604 309476 282610 309528
rect 281994 309340 282000 309392
rect 282052 309380 282058 309392
rect 282546 309380 282552 309392
rect 282052 309352 282552 309380
rect 282052 309340 282058 309352
rect 282546 309340 282552 309352
rect 282604 309340 282610 309392
rect 217410 309204 217416 309256
rect 217468 309244 217474 309256
rect 287146 309244 287152 309256
rect 217468 309216 287152 309244
rect 217468 309204 217474 309216
rect 287146 309204 287152 309216
rect 287204 309204 287210 309256
rect 213270 309136 213276 309188
rect 213328 309176 213334 309188
rect 285674 309176 285680 309188
rect 213328 309148 285680 309176
rect 213328 309136 213334 309148
rect 285674 309136 285680 309148
rect 285732 309136 285738 309188
rect 327718 309136 327724 309188
rect 327776 309176 327782 309188
rect 558914 309176 558920 309188
rect 327776 309148 558920 309176
rect 327776 309136 327782 309148
rect 558914 309136 558920 309148
rect 558972 309136 558978 309188
rect 214650 308456 214656 308508
rect 214708 308496 214714 308508
rect 288802 308496 288808 308508
rect 214708 308468 288808 308496
rect 214708 308456 214714 308468
rect 288802 308456 288808 308468
rect 288860 308456 288866 308508
rect 289446 308456 289452 308508
rect 289504 308496 289510 308508
rect 324406 308496 324412 308508
rect 289504 308468 324412 308496
rect 289504 308456 289510 308468
rect 324406 308456 324412 308468
rect 324464 308456 324470 308508
rect 210970 308388 210976 308440
rect 211028 308428 211034 308440
rect 285950 308428 285956 308440
rect 211028 308400 285956 308428
rect 211028 308388 211034 308400
rect 285950 308388 285956 308400
rect 286008 308388 286014 308440
rect 313918 308388 313924 308440
rect 313976 308428 313982 308440
rect 314930 308428 314936 308440
rect 313976 308400 314936 308428
rect 313976 308388 313982 308400
rect 314930 308388 314936 308400
rect 314988 308428 314994 308440
rect 416774 308428 416780 308440
rect 314988 308400 416780 308428
rect 314988 308388 314994 308400
rect 416774 308388 416780 308400
rect 416832 308388 416838 308440
rect 327810 307776 327816 307828
rect 327868 307816 327874 307828
rect 523034 307816 523040 307828
rect 327868 307788 523040 307816
rect 327868 307776 327874 307788
rect 523034 307776 523040 307788
rect 523092 307776 523098 307828
rect 287882 307572 287888 307624
rect 287940 307612 287946 307624
rect 296990 307612 296996 307624
rect 287940 307584 296996 307612
rect 287940 307572 287946 307584
rect 296990 307572 296996 307584
rect 297048 307572 297054 307624
rect 275830 307504 275836 307556
rect 275888 307544 275894 307556
rect 288710 307544 288716 307556
rect 275888 307516 288716 307544
rect 275888 307504 275894 307516
rect 288710 307504 288716 307516
rect 288768 307504 288774 307556
rect 290550 307504 290556 307556
rect 290608 307544 290614 307556
rect 293402 307544 293408 307556
rect 290608 307516 293408 307544
rect 290608 307504 290614 307516
rect 293402 307504 293408 307516
rect 293460 307504 293466 307556
rect 288342 307436 288348 307488
rect 288400 307476 288406 307488
rect 303890 307476 303896 307488
rect 288400 307448 303896 307476
rect 288400 307436 288406 307448
rect 303890 307436 303896 307448
rect 303948 307436 303954 307488
rect 285582 307368 285588 307420
rect 285640 307408 285646 307420
rect 303798 307408 303804 307420
rect 285640 307380 303804 307408
rect 285640 307368 285646 307380
rect 303798 307368 303804 307380
rect 303856 307368 303862 307420
rect 217318 307300 217324 307352
rect 217376 307340 217382 307352
rect 276014 307340 276020 307352
rect 217376 307312 276020 307340
rect 217376 307300 217382 307312
rect 276014 307300 276020 307312
rect 276072 307300 276078 307352
rect 284202 307300 284208 307352
rect 284260 307340 284266 307352
rect 304258 307340 304264 307352
rect 284260 307312 304264 307340
rect 284260 307300 284266 307312
rect 304258 307300 304264 307312
rect 304316 307300 304322 307352
rect 222194 307232 222200 307284
rect 222252 307272 222258 307284
rect 283190 307272 283196 307284
rect 222252 307244 283196 307272
rect 222252 307232 222258 307244
rect 283190 307232 283196 307244
rect 283248 307232 283254 307284
rect 290458 307232 290464 307284
rect 290516 307272 290522 307284
rect 315666 307272 315672 307284
rect 290516 307244 315672 307272
rect 290516 307232 290522 307244
rect 315666 307232 315672 307244
rect 315724 307232 315730 307284
rect 214742 307164 214748 307216
rect 214800 307204 214806 307216
rect 285122 307204 285128 307216
rect 214800 307176 285128 307204
rect 214800 307164 214806 307176
rect 285122 307164 285128 307176
rect 285180 307164 285186 307216
rect 289354 307164 289360 307216
rect 289412 307204 289418 307216
rect 313274 307204 313280 307216
rect 289412 307176 313280 307204
rect 289412 307164 289418 307176
rect 313274 307164 313280 307176
rect 313332 307164 313338 307216
rect 215846 307096 215852 307148
rect 215904 307136 215910 307148
rect 285858 307136 285864 307148
rect 215904 307108 285864 307136
rect 215904 307096 215910 307108
rect 285858 307096 285864 307108
rect 285916 307096 285922 307148
rect 286686 307096 286692 307148
rect 286744 307136 286750 307148
rect 321554 307136 321560 307148
rect 286744 307108 321560 307136
rect 286744 307096 286750 307108
rect 321554 307096 321560 307108
rect 321612 307096 321618 307148
rect 220354 307028 220360 307080
rect 220412 307068 220418 307080
rect 294874 307068 294880 307080
rect 220412 307040 294880 307068
rect 220412 307028 220418 307040
rect 294874 307028 294880 307040
rect 294932 307028 294938 307080
rect 287790 306960 287796 307012
rect 287848 307000 287854 307012
rect 294414 307000 294420 307012
rect 287848 306972 294420 307000
rect 287848 306960 287854 306972
rect 294414 306960 294420 306972
rect 294472 306960 294478 307012
rect 280890 306348 280896 306400
rect 280948 306388 280954 306400
rect 289630 306388 289636 306400
rect 280948 306360 289636 306388
rect 280948 306348 280954 306360
rect 289630 306348 289636 306360
rect 289688 306348 289694 306400
rect 580442 306388 580448 306400
rect 292500 306360 580448 306388
rect 282086 306280 282092 306332
rect 282144 306320 282150 306332
rect 292500 306320 292528 306360
rect 580442 306348 580448 306360
rect 580500 306348 580506 306400
rect 282144 306292 292528 306320
rect 282144 306280 282150 306292
rect 260282 305668 260288 305720
rect 260340 305708 260346 305720
rect 282086 305708 282092 305720
rect 260340 305680 282092 305708
rect 260340 305668 260346 305680
rect 282086 305668 282092 305680
rect 282144 305668 282150 305720
rect 283742 305668 283748 305720
rect 283800 305708 283806 305720
rect 304166 305708 304172 305720
rect 283800 305680 304172 305708
rect 283800 305668 283806 305680
rect 304166 305668 304172 305680
rect 304224 305668 304230 305720
rect 268654 305600 268660 305652
rect 268712 305640 268718 305652
rect 327626 305640 327632 305652
rect 268712 305612 327632 305640
rect 268712 305600 268718 305612
rect 327626 305600 327632 305612
rect 327684 305640 327690 305652
rect 540974 305640 540980 305652
rect 327684 305612 540980 305640
rect 327684 305600 327690 305612
rect 540974 305600 540980 305612
rect 541032 305600 541038 305652
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 253106 305028 253112 305040
rect 3292 305000 253112 305028
rect 3292 304988 3298 305000
rect 253106 304988 253112 305000
rect 253164 304988 253170 305040
rect 247126 304444 247132 304496
rect 247184 304484 247190 304496
rect 275094 304484 275100 304496
rect 247184 304456 275100 304484
rect 247184 304444 247190 304456
rect 275094 304444 275100 304456
rect 275152 304444 275158 304496
rect 218698 304376 218704 304428
rect 218756 304416 218762 304428
rect 280614 304416 280620 304428
rect 218756 304388 280620 304416
rect 218756 304376 218762 304388
rect 280614 304376 280620 304388
rect 280672 304376 280678 304428
rect 220262 304308 220268 304360
rect 220320 304348 220326 304360
rect 296898 304348 296904 304360
rect 220320 304320 296904 304348
rect 220320 304308 220326 304320
rect 296898 304308 296904 304320
rect 296956 304308 296962 304360
rect 220170 304240 220176 304292
rect 220228 304280 220234 304292
rect 297542 304280 297548 304292
rect 220228 304252 297548 304280
rect 220228 304240 220234 304252
rect 297542 304240 297548 304252
rect 297600 304240 297606 304292
rect 314102 304240 314108 304292
rect 314160 304280 314166 304292
rect 327534 304280 327540 304292
rect 314160 304252 327540 304280
rect 314160 304240 314166 304252
rect 327534 304240 327540 304252
rect 327592 304280 327598 304292
rect 563054 304280 563060 304292
rect 327592 304252 563060 304280
rect 327592 304240 327598 304252
rect 563054 304240 563060 304252
rect 563112 304240 563118 304292
rect 274450 302880 274456 302932
rect 274508 302920 274514 302932
rect 318610 302920 318616 302932
rect 274508 302892 318616 302920
rect 274508 302880 274514 302892
rect 318610 302880 318616 302892
rect 318668 302920 318674 302932
rect 329650 302920 329656 302932
rect 318668 302892 329656 302920
rect 318668 302880 318674 302892
rect 329650 302880 329656 302892
rect 329708 302880 329714 302932
rect 245838 301928 245844 301980
rect 245896 301928 245902 301980
rect 245746 301724 245752 301776
rect 245804 301764 245810 301776
rect 245856 301764 245884 301928
rect 245804 301736 245884 301764
rect 245804 301724 245810 301736
rect 253106 301724 253112 301776
rect 253164 301764 253170 301776
rect 258810 301764 258816 301776
rect 253164 301736 258816 301764
rect 253164 301724 253170 301736
rect 258810 301724 258816 301736
rect 258868 301724 258874 301776
rect 240134 301520 240140 301572
rect 240192 301560 240198 301572
rect 240318 301560 240324 301572
rect 240192 301532 240324 301560
rect 240192 301520 240198 301532
rect 240318 301520 240324 301532
rect 240376 301520 240382 301572
rect 221550 301452 221556 301504
rect 221608 301492 221614 301504
rect 302510 301492 302516 301504
rect 221608 301464 302516 301492
rect 221608 301452 221614 301464
rect 302510 301452 302516 301464
rect 302568 301452 302574 301504
rect 329098 300840 329104 300892
rect 329156 300880 329162 300892
rect 445754 300880 445760 300892
rect 329156 300852 445760 300880
rect 329156 300840 329162 300852
rect 445754 300840 445760 300852
rect 445812 300840 445818 300892
rect 258810 300772 258816 300824
rect 258868 300812 258874 300824
rect 259086 300812 259092 300824
rect 258868 300784 259092 300812
rect 258868 300772 258874 300784
rect 259086 300772 259092 300784
rect 259144 300812 259150 300824
rect 275186 300812 275192 300824
rect 259144 300784 275192 300812
rect 259144 300772 259150 300784
rect 275186 300772 275192 300784
rect 275244 300772 275250 300824
rect 304258 300364 304264 300416
rect 304316 300404 304322 300416
rect 305546 300404 305552 300416
rect 304316 300376 305552 300404
rect 304316 300364 304322 300376
rect 305546 300364 305552 300376
rect 305604 300364 305610 300416
rect 329650 300092 329656 300144
rect 329708 300132 329714 300144
rect 452654 300132 452660 300144
rect 329708 300104 452660 300132
rect 329708 300092 329714 300104
rect 452654 300092 452660 300104
rect 452712 300092 452718 300144
rect 256786 299480 256792 299532
rect 256844 299520 256850 299532
rect 257614 299520 257620 299532
rect 256844 299492 257620 299520
rect 256844 299480 256850 299492
rect 257614 299480 257620 299492
rect 257672 299480 257678 299532
rect 253934 298868 253940 298920
rect 253992 298908 253998 298920
rect 254670 298908 254676 298920
rect 253992 298880 254676 298908
rect 253992 298868 253998 298880
rect 254670 298868 254676 298880
rect 254728 298868 254734 298920
rect 229462 298800 229468 298852
rect 229520 298840 229526 298852
rect 242158 298840 242164 298852
rect 229520 298812 242164 298840
rect 229520 298800 229526 298812
rect 242158 298800 242164 298812
rect 242216 298800 242222 298852
rect 221458 298732 221464 298784
rect 221516 298772 221522 298784
rect 302418 298772 302424 298784
rect 221516 298744 302424 298772
rect 221516 298732 221522 298744
rect 302418 298732 302424 298744
rect 302476 298732 302482 298784
rect 332042 298732 332048 298784
rect 332100 298772 332106 298784
rect 572806 298772 572812 298784
rect 332100 298744 572812 298772
rect 332100 298732 332106 298744
rect 572806 298732 572812 298744
rect 572864 298732 572870 298784
rect 256694 297440 256700 297492
rect 256752 297480 256758 297492
rect 257246 297480 257252 297492
rect 256752 297452 257252 297480
rect 256752 297440 256758 297452
rect 257246 297440 257252 297452
rect 257304 297440 257310 297492
rect 232958 297372 232964 297424
rect 233016 297412 233022 297424
rect 277854 297412 277860 297424
rect 233016 297384 277860 297412
rect 233016 297372 233022 297384
rect 277854 297372 277860 297384
rect 277912 297372 277918 297424
rect 316678 297372 316684 297424
rect 316736 297412 316742 297424
rect 330570 297412 330576 297424
rect 316736 297384 330576 297412
rect 316736 297372 316742 297384
rect 330570 297372 330576 297384
rect 330628 297412 330634 297424
rect 456794 297412 456800 297424
rect 330628 297384 456800 297412
rect 330628 297372 330634 297384
rect 456794 297372 456800 297384
rect 456852 297372 456858 297424
rect 255406 297304 255412 297356
rect 255464 297344 255470 297356
rect 256326 297344 256332 297356
rect 255464 297316 256332 297344
rect 255464 297304 255470 297316
rect 256326 297304 256332 297316
rect 256384 297304 256390 297356
rect 256878 297304 256884 297356
rect 256936 297344 256942 297356
rect 257062 297344 257068 297356
rect 256936 297316 257068 297344
rect 256936 297304 256942 297316
rect 257062 297304 257068 297316
rect 257120 297304 257126 297356
rect 226886 296692 226892 296744
rect 226944 296732 226950 296744
rect 231118 296732 231124 296744
rect 226944 296704 231124 296732
rect 226944 296692 226950 296704
rect 231118 296692 231124 296704
rect 231176 296692 231182 296744
rect 244550 296012 244556 296064
rect 244608 296052 244614 296064
rect 277946 296052 277952 296064
rect 244608 296024 277952 296052
rect 244608 296012 244614 296024
rect 277946 296012 277952 296024
rect 278004 296012 278010 296064
rect 222286 295944 222292 295996
rect 222344 295984 222350 295996
rect 283374 295984 283380 295996
rect 222344 295956 283380 295984
rect 222344 295944 222350 295956
rect 283374 295944 283380 295956
rect 283432 295944 283438 295996
rect 258166 294652 258172 294704
rect 258224 294692 258230 294704
rect 258534 294692 258540 294704
rect 258224 294664 258540 294692
rect 258224 294652 258230 294664
rect 258534 294652 258540 294664
rect 258592 294652 258598 294704
rect 235718 294584 235724 294636
rect 235776 294624 235782 294636
rect 278590 294624 278596 294636
rect 235776 294596 278596 294624
rect 235776 294584 235782 294596
rect 278590 294584 278596 294596
rect 278648 294584 278654 294636
rect 318058 294584 318064 294636
rect 318116 294624 318122 294636
rect 329190 294624 329196 294636
rect 318116 294596 329196 294624
rect 318116 294584 318122 294596
rect 329190 294584 329196 294596
rect 329248 294624 329254 294636
rect 463694 294624 463700 294636
rect 329248 294596 463700 294624
rect 329248 294584 329254 294596
rect 463694 294584 463700 294596
rect 463752 294584 463758 294636
rect 312170 293972 312176 294024
rect 312228 294012 312234 294024
rect 312722 294012 312728 294024
rect 312228 293984 312728 294012
rect 312228 293972 312234 293984
rect 312722 293972 312728 293984
rect 312780 294012 312786 294024
rect 382274 294012 382280 294024
rect 312780 293984 382280 294012
rect 312780 293972 312786 293984
rect 382274 293972 382280 293984
rect 382332 293972 382338 294024
rect 248230 293904 248236 293956
rect 248288 293944 248294 293956
rect 250438 293944 250444 293956
rect 248288 293916 250444 293944
rect 248288 293904 248294 293916
rect 250438 293904 250444 293916
rect 250496 293904 250502 293956
rect 233878 293564 233884 293616
rect 233936 293604 233942 293616
rect 247586 293604 247592 293616
rect 233936 293576 247592 293604
rect 233936 293564 233942 293576
rect 247586 293564 247592 293576
rect 247644 293564 247650 293616
rect 231670 293496 231676 293548
rect 231728 293536 231734 293548
rect 245010 293536 245016 293548
rect 231728 293508 245016 293536
rect 231728 293496 231734 293508
rect 245010 293496 245016 293508
rect 245068 293496 245074 293548
rect 228358 293428 228364 293480
rect 228416 293468 228422 293480
rect 243538 293468 243544 293480
rect 228416 293440 243544 293468
rect 228416 293428 228422 293440
rect 243538 293428 243544 293440
rect 243596 293428 243602 293480
rect 236086 293360 236092 293412
rect 236144 293400 236150 293412
rect 278498 293400 278504 293412
rect 236144 293372 278504 293400
rect 236144 293360 236150 293372
rect 278498 293360 278504 293372
rect 278556 293360 278562 293412
rect 223942 293292 223948 293344
rect 224000 293332 224006 293344
rect 280706 293332 280712 293344
rect 224000 293304 280712 293332
rect 224000 293292 224006 293304
rect 280706 293292 280712 293304
rect 280764 293292 280770 293344
rect 3418 293224 3424 293276
rect 3476 293264 3482 293276
rect 258718 293264 258724 293276
rect 3476 293236 258724 293264
rect 3476 293224 3482 293236
rect 258718 293224 258724 293236
rect 258776 293224 258782 293276
rect 334710 293224 334716 293276
rect 334768 293264 334774 293276
rect 466454 293264 466460 293276
rect 334768 293236 466460 293264
rect 334768 293224 334774 293236
rect 466454 293224 466460 293236
rect 466512 293224 466518 293276
rect 223758 293020 223764 293072
rect 223816 293060 223822 293072
rect 224494 293060 224500 293072
rect 223816 293032 224500 293060
rect 223816 293020 223822 293032
rect 224494 293020 224500 293032
rect 224552 293020 224558 293072
rect 225046 293020 225052 293072
rect 225104 293060 225110 293072
rect 225966 293060 225972 293072
rect 225104 293032 225972 293060
rect 225104 293020 225110 293032
rect 225966 293020 225972 293032
rect 226024 293020 226030 293072
rect 226334 293020 226340 293072
rect 226392 293060 226398 293072
rect 227070 293060 227076 293072
rect 226392 293032 227076 293060
rect 226392 293020 226398 293032
rect 227070 293020 227076 293032
rect 227128 293020 227134 293072
rect 230474 293020 230480 293072
rect 230532 293060 230538 293072
rect 231118 293060 231124 293072
rect 230532 293032 231124 293060
rect 230532 293020 230538 293032
rect 231118 293020 231124 293032
rect 231176 293020 231182 293072
rect 235994 293020 236000 293072
rect 236052 293060 236058 293072
rect 237006 293060 237012 293072
rect 236052 293032 237012 293060
rect 236052 293020 236058 293032
rect 237006 293020 237012 293032
rect 237064 293020 237070 293072
rect 241514 293020 241520 293072
rect 241572 293060 241578 293072
rect 242158 293060 242164 293072
rect 241572 293032 242164 293060
rect 241572 293020 241578 293032
rect 242158 293020 242164 293032
rect 242216 293020 242222 293072
rect 242894 293020 242900 293072
rect 242952 293060 242958 293072
rect 243262 293060 243268 293072
rect 242952 293032 243268 293060
rect 242952 293020 242958 293032
rect 243262 293020 243268 293032
rect 243320 293020 243326 293072
rect 245746 293020 245752 293072
rect 245804 293060 245810 293072
rect 246574 293060 246580 293072
rect 245804 293032 246580 293060
rect 245804 293020 245810 293032
rect 246574 293020 246580 293032
rect 246632 293020 246638 293072
rect 247034 293020 247040 293072
rect 247092 293060 247098 293072
rect 247678 293060 247684 293072
rect 247092 293032 247684 293060
rect 247092 293020 247098 293032
rect 247678 293020 247684 293032
rect 247736 293020 247742 293072
rect 249794 293020 249800 293072
rect 249852 293060 249858 293072
rect 250254 293060 250260 293072
rect 249852 293032 250260 293060
rect 249852 293020 249858 293032
rect 250254 293020 250260 293032
rect 250312 293020 250318 293072
rect 251266 293020 251272 293072
rect 251324 293060 251330 293072
rect 252094 293060 252100 293072
rect 251324 293032 252100 293060
rect 251324 293020 251330 293032
rect 252094 293020 252100 293032
rect 252152 293020 252158 293072
rect 252646 293020 252652 293072
rect 252704 293060 252710 293072
rect 253198 293060 253204 293072
rect 252704 293032 253204 293060
rect 252704 293020 252710 293032
rect 253198 293020 253204 293032
rect 253256 293020 253262 293072
rect 242986 292952 242992 293004
rect 243044 292992 243050 293004
rect 243998 292992 244004 293004
rect 243044 292964 244004 292992
rect 243044 292952 243050 292964
rect 243998 292952 244004 292964
rect 244056 292952 244062 293004
rect 252554 292952 252560 293004
rect 252612 292992 252618 293004
rect 253566 292992 253572 293004
rect 252612 292964 253572 292992
rect 252612 292952 252618 292964
rect 253566 292952 253572 292964
rect 253624 292952 253630 293004
rect 220078 292544 220084 292596
rect 220136 292584 220142 292596
rect 223942 292584 223948 292596
rect 220136 292556 223948 292584
rect 220136 292544 220142 292556
rect 223942 292544 223948 292556
rect 224000 292544 224006 292596
rect 319438 292544 319444 292596
rect 319496 292584 319502 292596
rect 481634 292584 481640 292596
rect 319496 292556 481640 292584
rect 319496 292544 319502 292556
rect 481634 292544 481640 292556
rect 481692 292544 481698 292596
rect 238294 292476 238300 292528
rect 238352 292516 238358 292528
rect 239398 292516 239404 292528
rect 238352 292488 239404 292516
rect 238352 292476 238358 292488
rect 239398 292476 239404 292488
rect 239456 292476 239462 292528
rect 259638 292476 259644 292528
rect 259696 292516 259702 292528
rect 260190 292516 260196 292528
rect 259696 292488 260196 292516
rect 259696 292476 259702 292488
rect 260190 292476 260196 292488
rect 260248 292476 260254 292528
rect 262122 292476 262128 292528
rect 262180 292516 262186 292528
rect 262582 292516 262588 292528
rect 262180 292488 262588 292516
rect 262180 292476 262186 292488
rect 262582 292476 262588 292488
rect 262640 292476 262646 292528
rect 264238 292476 264244 292528
rect 264296 292516 264302 292528
rect 264790 292516 264796 292528
rect 264296 292488 264796 292516
rect 264296 292476 264302 292488
rect 264790 292476 264796 292488
rect 264848 292476 264854 292528
rect 234982 292136 234988 292188
rect 235040 292176 235046 292188
rect 236546 292176 236552 292188
rect 235040 292148 236552 292176
rect 235040 292136 235046 292148
rect 236546 292136 236552 292148
rect 236604 292136 236610 292188
rect 244918 292176 244924 292188
rect 236656 292148 244924 292176
rect 236362 292068 236368 292120
rect 236420 292108 236426 292120
rect 236656 292108 236684 292148
rect 244918 292136 244924 292148
rect 244976 292136 244982 292188
rect 253106 292108 253112 292120
rect 236420 292080 236684 292108
rect 236748 292080 253112 292108
rect 236420 292068 236426 292080
rect 234246 292000 234252 292052
rect 234304 292040 234310 292052
rect 236748 292040 236776 292080
rect 253106 292068 253112 292080
rect 253164 292068 253170 292120
rect 260282 292040 260288 292052
rect 234304 292012 236776 292040
rect 236840 292012 260288 292040
rect 234304 292000 234310 292012
rect 232038 291932 232044 291984
rect 232096 291972 232102 291984
rect 236840 291972 236868 292012
rect 260282 292000 260288 292012
rect 260340 292000 260346 292052
rect 263686 292000 263692 292052
rect 263744 292040 263750 292052
rect 275922 292040 275928 292052
rect 263744 292012 275928 292040
rect 263744 292000 263750 292012
rect 275922 292000 275928 292012
rect 275980 292000 275986 292052
rect 232096 291944 236868 291972
rect 232096 291932 232102 291944
rect 237558 291932 237564 291984
rect 237616 291972 237622 291984
rect 281074 291972 281080 291984
rect 237616 291944 281080 291972
rect 237616 291932 237622 291944
rect 281074 291932 281080 291944
rect 281132 291932 281138 291984
rect 235350 291864 235356 291916
rect 235408 291904 235414 291916
rect 281166 291904 281172 291916
rect 235408 291876 281172 291904
rect 235408 291864 235414 291876
rect 281166 291864 281172 291876
rect 281224 291864 281230 291916
rect 318242 291864 318248 291916
rect 318300 291904 318306 291916
rect 331674 291904 331680 291916
rect 318300 291876 331680 291904
rect 318300 291864 318306 291876
rect 331674 291864 331680 291876
rect 331732 291904 331738 291916
rect 331732 291876 335354 291904
rect 331732 291864 331738 291876
rect 217226 291796 217232 291848
rect 217284 291836 217290 291848
rect 262582 291836 262588 291848
rect 217284 291808 262588 291836
rect 217284 291796 217290 291808
rect 262582 291796 262588 291808
rect 262640 291796 262646 291848
rect 265894 291796 265900 291848
rect 265952 291836 265958 291848
rect 329006 291836 329012 291848
rect 265952 291808 329012 291836
rect 265952 291796 265958 291808
rect 329006 291796 329012 291808
rect 329064 291796 329070 291848
rect 335326 291836 335354 291876
rect 470594 291836 470600 291848
rect 335326 291808 470600 291836
rect 470594 291796 470600 291808
rect 470652 291796 470658 291848
rect 262306 291728 262312 291780
rect 262364 291768 262370 291780
rect 262766 291768 262772 291780
rect 262364 291740 262772 291768
rect 262364 291728 262370 291740
rect 262766 291728 262772 291740
rect 262824 291728 262830 291780
rect 197998 291660 198004 291712
rect 198056 291700 198062 291712
rect 263686 291700 263692 291712
rect 198056 291672 263692 291700
rect 198056 291660 198062 291672
rect 263686 291660 263692 291672
rect 263744 291660 263750 291712
rect 195238 291592 195244 291644
rect 195296 291632 195302 291644
rect 264790 291632 264796 291644
rect 195296 291604 264796 291632
rect 195296 291592 195302 291604
rect 264790 291592 264796 291604
rect 264848 291592 264854 291644
rect 225046 291524 225052 291576
rect 225104 291564 225110 291576
rect 226978 291564 226984 291576
rect 225104 291536 226984 291564
rect 225104 291524 225110 291536
rect 226978 291524 226984 291536
rect 227036 291524 227042 291576
rect 232222 291524 232228 291576
rect 232280 291564 232286 291576
rect 259638 291564 259644 291576
rect 232280 291536 259644 291564
rect 232280 291524 232286 291536
rect 259638 291524 259644 291536
rect 259696 291524 259702 291576
rect 226518 291456 226524 291508
rect 226576 291496 226582 291508
rect 256142 291496 256148 291508
rect 226576 291468 256148 291496
rect 226576 291456 226582 291468
rect 256142 291456 256148 291468
rect 256200 291456 256206 291508
rect 220906 291388 220912 291440
rect 220964 291428 220970 291440
rect 260098 291428 260104 291440
rect 220964 291400 260104 291428
rect 220964 291388 220970 291400
rect 260098 291388 260104 291400
rect 260156 291388 260162 291440
rect 219894 291320 219900 291372
rect 219952 291360 219958 291372
rect 261478 291360 261484 291372
rect 219952 291332 261484 291360
rect 219952 291320 219958 291332
rect 261478 291320 261484 291332
rect 261536 291320 261542 291372
rect 222010 291252 222016 291304
rect 222068 291292 222074 291304
rect 222068 291264 225460 291292
rect 222068 291252 222074 291264
rect 225432 291236 225460 291264
rect 222102 291184 222108 291236
rect 222160 291224 222166 291236
rect 224218 291224 224224 291236
rect 222160 291196 224224 291224
rect 222160 291184 222166 291196
rect 224218 291184 224224 291196
rect 224276 291184 224282 291236
rect 225414 291184 225420 291236
rect 225472 291224 225478 291236
rect 225598 291224 225604 291236
rect 225472 291196 225604 291224
rect 225472 291184 225478 291196
rect 225598 291184 225604 291196
rect 225656 291184 225662 291236
rect 230934 291184 230940 291236
rect 230992 291224 230998 291236
rect 230992 291196 246988 291224
rect 230992 291184 230998 291196
rect 246960 291156 246988 291196
rect 281350 291156 281356 291168
rect 246960 291128 281356 291156
rect 281350 291116 281356 291128
rect 281408 291116 281414 291168
rect 264882 290844 264888 290896
rect 264940 290884 264946 290896
rect 265526 290884 265532 290896
rect 264940 290856 265532 290884
rect 264940 290844 264946 290856
rect 265526 290844 265532 290856
rect 265584 290844 265590 290896
rect 239766 290640 239772 290692
rect 239824 290680 239830 290692
rect 255958 290680 255964 290692
rect 239824 290652 255964 290680
rect 239824 290640 239830 290652
rect 255958 290640 255964 290652
rect 256016 290640 256022 290692
rect 240870 290572 240876 290624
rect 240928 290612 240934 290624
rect 257338 290612 257344 290624
rect 240928 290584 257344 290612
rect 240928 290572 240934 290584
rect 257338 290572 257344 290584
rect 257396 290572 257402 290624
rect 116578 290504 116584 290556
rect 116636 290544 116642 290556
rect 264882 290544 264888 290556
rect 116636 290516 264888 290544
rect 116636 290504 116642 290516
rect 264882 290504 264888 290516
rect 264940 290504 264946 290556
rect 3510 290436 3516 290488
rect 3568 290476 3574 290488
rect 232222 290476 232228 290488
rect 3568 290448 232228 290476
rect 3568 290436 3574 290448
rect 232222 290436 232228 290448
rect 232280 290436 232286 290488
rect 243814 290436 243820 290488
rect 243872 290476 243878 290488
rect 275738 290476 275744 290488
rect 243872 290448 275744 290476
rect 243872 290436 243878 290448
rect 275738 290436 275744 290448
rect 275796 290436 275802 290488
rect 281350 290436 281356 290488
rect 281408 290476 281414 290488
rect 580718 290476 580724 290488
rect 281408 290448 580724 290476
rect 281408 290436 281414 290448
rect 580718 290436 580724 290448
rect 580776 290436 580782 290488
rect 219986 290096 219992 290148
rect 220044 290136 220050 290148
rect 259822 290136 259828 290148
rect 220044 290108 259828 290136
rect 220044 290096 220050 290108
rect 259822 290096 259828 290108
rect 259880 290096 259886 290148
rect 262490 290096 262496 290148
rect 262548 290136 262554 290148
rect 263318 290136 263324 290148
rect 262548 290108 263324 290136
rect 262548 290096 262554 290108
rect 263318 290096 263324 290108
rect 263376 290096 263382 290148
rect 229278 290028 229284 290080
rect 229336 290068 229342 290080
rect 229738 290068 229744 290080
rect 229336 290040 229744 290068
rect 229336 290028 229342 290040
rect 229738 290028 229744 290040
rect 229796 290068 229802 290080
rect 269942 290068 269948 290080
rect 229796 290040 269948 290068
rect 229796 290028 229802 290040
rect 269942 290028 269948 290040
rect 270000 290028 270006 290080
rect 213454 289960 213460 290012
rect 213512 290000 213518 290012
rect 260926 290000 260932 290012
rect 213512 289972 260932 290000
rect 213512 289960 213518 289972
rect 260926 289960 260932 289972
rect 260984 289960 260990 290012
rect 203518 289892 203524 289944
rect 203576 289932 203582 289944
rect 262122 289932 262128 289944
rect 203576 289904 262128 289932
rect 203576 289892 203582 289904
rect 262122 289892 262128 289904
rect 262180 289892 262186 289944
rect 192478 289824 192484 289876
rect 192536 289864 192542 289876
rect 262490 289864 262496 289876
rect 192536 289836 262496 289864
rect 192536 289824 192542 289836
rect 262490 289824 262496 289836
rect 262548 289824 262554 289876
rect 256142 289756 256148 289808
rect 256200 289796 256206 289808
rect 256510 289796 256516 289808
rect 256200 289768 256516 289796
rect 256200 289756 256206 289768
rect 256510 289756 256516 289768
rect 256568 289756 256574 289808
rect 259546 289756 259552 289808
rect 259604 289796 259610 289808
rect 260558 289796 260564 289808
rect 259604 289768 260564 289796
rect 259604 289756 259610 289768
rect 260558 289756 260564 289768
rect 260616 289756 260622 289808
rect 261294 289756 261300 289808
rect 261352 289796 261358 289808
rect 261662 289796 261668 289808
rect 261352 289768 261668 289796
rect 261352 289756 261358 289768
rect 261662 289756 261668 289768
rect 261720 289756 261726 289808
rect 249242 289620 249248 289672
rect 249300 289660 249306 289672
rect 249300 289632 258074 289660
rect 249300 289620 249306 289632
rect 227686 289564 249380 289592
rect 211798 289212 211804 289264
rect 211856 289252 211862 289264
rect 227686 289252 227714 289564
rect 249242 289484 249248 289536
rect 249300 289484 249306 289536
rect 249260 289388 249288 289484
rect 211856 289224 227714 289252
rect 241486 289360 245654 289388
rect 211856 289212 211862 289224
rect 199378 289144 199384 289196
rect 199436 289184 199442 289196
rect 222470 289184 222476 289196
rect 199436 289156 222476 289184
rect 199436 289144 199442 289156
rect 222470 289144 222476 289156
rect 222528 289144 222534 289196
rect 227180 289156 240134 289184
rect 91738 289076 91744 289128
rect 91796 289116 91802 289128
rect 91796 289088 219434 289116
rect 91796 289076 91802 289088
rect 219406 289048 219434 289088
rect 227180 289048 227208 289156
rect 240106 289116 240134 289156
rect 241486 289116 241514 289360
rect 245626 289252 245654 289360
rect 248386 289360 249288 289388
rect 248386 289252 248414 289360
rect 249352 289320 249380 289564
rect 258046 289524 258074 289632
rect 262766 289592 262772 289604
rect 261128 289564 262772 289592
rect 259546 289524 259552 289536
rect 258046 289496 259552 289524
rect 259546 289484 259552 289496
rect 259604 289484 259610 289536
rect 249352 289292 258074 289320
rect 245626 289224 248414 289252
rect 258046 289252 258074 289292
rect 261128 289252 261156 289564
rect 262766 289552 262772 289564
rect 262824 289552 262830 289604
rect 261294 289484 261300 289536
rect 261352 289484 261358 289536
rect 258046 289224 261156 289252
rect 261312 289184 261340 289484
rect 240106 289088 241514 289116
rect 249628 289156 261340 289184
rect 219406 289020 227208 289048
rect 249628 288980 249656 289156
rect 248386 288952 249656 288980
rect 248386 288912 248414 288952
rect 245626 288884 248414 288912
rect 222470 288804 222476 288856
rect 222528 288844 222534 288856
rect 245626 288844 245654 288884
rect 222528 288816 245654 288844
rect 222528 288804 222534 288816
rect 3418 286288 3424 286340
rect 3476 286328 3482 286340
rect 220906 286328 220912 286340
rect 3476 286300 220912 286328
rect 3476 286288 3482 286300
rect 220906 286288 220912 286300
rect 220964 286288 220970 286340
rect 270218 284928 270224 284980
rect 270276 284968 270282 284980
rect 290918 284968 290924 284980
rect 270276 284940 290924 284968
rect 270276 284928 270282 284940
rect 290918 284928 290924 284940
rect 290976 284928 290982 284980
rect 271782 283568 271788 283620
rect 271840 283608 271846 283620
rect 284570 283608 284576 283620
rect 271840 283580 284576 283608
rect 271840 283568 271846 283580
rect 284570 283568 284576 283580
rect 284628 283568 284634 283620
rect 271046 282140 271052 282192
rect 271104 282180 271110 282192
rect 286042 282180 286048 282192
rect 271104 282152 286048 282180
rect 271104 282140 271110 282152
rect 286042 282140 286048 282152
rect 286100 282140 286106 282192
rect 270310 275272 270316 275324
rect 270368 275312 270374 275324
rect 290734 275312 290740 275324
rect 270368 275284 290740 275312
rect 270368 275272 270374 275284
rect 290734 275272 290740 275284
rect 290792 275272 290798 275324
rect 270954 273912 270960 273964
rect 271012 273952 271018 273964
rect 283466 273952 283472 273964
rect 271012 273924 283472 273952
rect 271012 273912 271018 273924
rect 283466 273912 283472 273924
rect 283524 273912 283530 273964
rect 330478 273164 330484 273216
rect 330536 273204 330542 273216
rect 580166 273204 580172 273216
rect 330536 273176 580172 273204
rect 330536 273164 330542 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 320542 271804 320548 271856
rect 320600 271844 320606 271856
rect 321094 271844 321100 271856
rect 320600 271816 321100 271844
rect 320600 271804 320606 271816
rect 321094 271804 321100 271816
rect 321152 271804 321158 271856
rect 321094 270512 321100 270564
rect 321152 270552 321158 270564
rect 498194 270552 498200 270564
rect 321152 270524 498200 270552
rect 321152 270512 321158 270524
rect 498194 270512 498200 270524
rect 498252 270512 498258 270564
rect 313458 269016 313464 269068
rect 313516 269056 313522 269068
rect 314194 269056 314200 269068
rect 313516 269028 314200 269056
rect 313516 269016 313522 269028
rect 314194 269016 314200 269028
rect 314252 269016 314258 269068
rect 314194 267724 314200 267776
rect 314252 267764 314258 267776
rect 407206 267764 407212 267776
rect 314252 267736 407212 267764
rect 314252 267724 314258 267736
rect 407206 267724 407212 267736
rect 407264 267724 407270 267776
rect 319070 265820 319076 265872
rect 319128 265860 319134 265872
rect 319622 265860 319628 265872
rect 319128 265832 319628 265860
rect 319128 265820 319134 265832
rect 319622 265820 319628 265832
rect 319680 265820 319686 265872
rect 319622 264936 319628 264988
rect 319680 264976 319686 264988
rect 467834 264976 467840 264988
rect 319680 264948 467840 264976
rect 319680 264936 319686 264948
rect 467834 264936 467840 264948
rect 467892 264936 467898 264988
rect 270402 264188 270408 264240
rect 270460 264228 270466 264240
rect 291562 264228 291568 264240
rect 270460 264200 291568 264228
rect 270460 264188 270466 264200
rect 291562 264188 291568 264200
rect 291620 264188 291626 264240
rect 312078 263576 312084 263628
rect 312136 263616 312142 263628
rect 313458 263616 313464 263628
rect 312136 263588 313464 263616
rect 312136 263576 312142 263588
rect 313458 263576 313464 263588
rect 313516 263616 313522 263628
rect 386414 263616 386420 263628
rect 313516 263588 386420 263616
rect 313516 263576 313522 263588
rect 386414 263576 386420 263588
rect 386472 263576 386478 263628
rect 316310 262624 316316 262676
rect 316368 262664 316374 262676
rect 316770 262664 316776 262676
rect 316368 262636 316776 262664
rect 316368 262624 316374 262636
rect 316770 262624 316776 262636
rect 316828 262624 316834 262676
rect 316770 262216 316776 262268
rect 316828 262256 316834 262268
rect 438854 262256 438860 262268
rect 316828 262228 438860 262256
rect 316828 262216 316834 262228
rect 438854 262216 438860 262228
rect 438912 262216 438918 262268
rect 269666 260108 269672 260160
rect 269724 260148 269730 260160
rect 290826 260148 290832 260160
rect 269724 260120 290832 260148
rect 269724 260108 269730 260120
rect 290826 260108 290832 260120
rect 290884 260108 290890 260160
rect 306834 260108 306840 260160
rect 306892 260148 306898 260160
rect 320542 260148 320548 260160
rect 306892 260120 320548 260148
rect 306892 260108 306898 260120
rect 320542 260108 320548 260120
rect 320600 260108 320606 260160
rect 349154 259468 349160 259480
rect 309520 259440 349160 259468
rect 309520 259412 309548 259440
rect 349154 259428 349160 259440
rect 349212 259428 349218 259480
rect 308950 259360 308956 259412
rect 309008 259400 309014 259412
rect 309502 259400 309508 259412
rect 309008 259372 309508 259400
rect 309008 259360 309014 259372
rect 309502 259360 309508 259372
rect 309560 259360 309566 259412
rect 313366 259360 313372 259412
rect 313424 259400 313430 259412
rect 314378 259400 314384 259412
rect 313424 259372 314384 259400
rect 313424 259360 313430 259372
rect 314378 259360 314384 259372
rect 314436 259360 314442 259412
rect 320450 259360 320456 259412
rect 320508 259400 320514 259412
rect 321002 259400 321008 259412
rect 320508 259372 321008 259400
rect 320508 259360 320514 259372
rect 321002 259360 321008 259372
rect 321060 259360 321066 259412
rect 363598 259360 363604 259412
rect 363656 259400 363662 259412
rect 579798 259400 579804 259412
rect 363656 259372 579804 259400
rect 363656 259360 363662 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 314378 258136 314384 258188
rect 314436 258176 314442 258188
rect 402974 258176 402980 258188
rect 314436 258148 402980 258176
rect 314436 258136 314442 258148
rect 402974 258136 402980 258148
rect 403032 258136 403038 258188
rect 321002 258068 321008 258120
rect 321060 258108 321066 258120
rect 496814 258108 496820 258120
rect 321060 258080 496820 258108
rect 321060 258068 321066 258080
rect 496814 258068 496820 258080
rect 496872 258068 496878 258120
rect 319530 255280 319536 255332
rect 319588 255320 319594 255332
rect 320082 255320 320088 255332
rect 319588 255292 320088 255320
rect 319588 255280 319594 255292
rect 320082 255280 320088 255292
rect 320140 255320 320146 255332
rect 481726 255320 481732 255332
rect 320140 255292 481732 255320
rect 320140 255280 320146 255292
rect 481726 255280 481732 255292
rect 481784 255280 481790 255332
rect 314562 253920 314568 253972
rect 314620 253960 314626 253972
rect 314838 253960 314844 253972
rect 314620 253932 314844 253960
rect 314620 253920 314626 253932
rect 314838 253920 314844 253932
rect 314896 253960 314902 253972
rect 420914 253960 420920 253972
rect 314896 253932 420920 253960
rect 314896 253920 314902 253932
rect 420914 253920 420920 253932
rect 420972 253920 420978 253972
rect 3510 253172 3516 253224
rect 3568 253212 3574 253224
rect 219894 253212 219900 253224
rect 3568 253184 219900 253212
rect 3568 253172 3574 253184
rect 219894 253172 219900 253184
rect 219952 253172 219958 253224
rect 321922 252560 321928 252612
rect 321980 252600 321986 252612
rect 322290 252600 322296 252612
rect 321980 252572 322296 252600
rect 321980 252560 321986 252572
rect 322290 252560 322296 252572
rect 322348 252600 322354 252612
rect 510614 252600 510620 252612
rect 322348 252572 510620 252600
rect 322348 252560 322354 252572
rect 510614 252560 510620 252572
rect 510672 252560 510678 252612
rect 321830 252492 321836 252544
rect 321888 252532 321894 252544
rect 322566 252532 322572 252544
rect 321888 252504 322572 252532
rect 321888 252492 321894 252504
rect 322566 252492 322572 252504
rect 322624 252492 322630 252544
rect 269574 251812 269580 251864
rect 269632 251852 269638 251864
rect 291470 251852 291476 251864
rect 269632 251824 291476 251852
rect 269632 251812 269638 251824
rect 291470 251812 291476 251824
rect 291528 251812 291534 251864
rect 322566 251200 322572 251252
rect 322624 251240 322630 251252
rect 506474 251240 506480 251252
rect 322624 251212 506480 251240
rect 322624 251200 322630 251212
rect 506474 251200 506480 251212
rect 506532 251200 506538 251252
rect 312906 250452 312912 250504
rect 312964 250492 312970 250504
rect 326430 250492 326436 250504
rect 312964 250464 326436 250492
rect 312964 250452 312970 250464
rect 326430 250452 326436 250464
rect 326488 250492 326494 250504
rect 385034 250492 385040 250504
rect 326488 250464 385040 250492
rect 326488 250452 326494 250464
rect 385034 250452 385040 250464
rect 385092 250452 385098 250504
rect 314286 249024 314292 249076
rect 314344 249064 314350 249076
rect 322382 249064 322388 249076
rect 314344 249036 322388 249064
rect 314344 249024 314350 249036
rect 322382 249024 322388 249036
rect 322440 249064 322446 249076
rect 398834 249064 398840 249076
rect 322440 249036 398840 249064
rect 322440 249024 322446 249036
rect 398834 249024 398840 249036
rect 398892 249024 398898 249076
rect 312814 248412 312820 248464
rect 312872 248452 312878 248464
rect 389174 248452 389180 248464
rect 312872 248424 389180 248452
rect 312872 248412 312878 248424
rect 389174 248412 389180 248424
rect 389232 248412 389238 248464
rect 321738 247868 321744 247920
rect 321796 247908 321802 247920
rect 322382 247908 322388 247920
rect 321796 247880 322388 247908
rect 321796 247868 321802 247880
rect 322382 247868 322388 247880
rect 322440 247868 322446 247920
rect 316218 247120 316224 247172
rect 316276 247160 316282 247172
rect 442994 247160 443000 247172
rect 316276 247132 443000 247160
rect 316276 247120 316282 247132
rect 442994 247120 443000 247132
rect 443052 247120 443058 247172
rect 322382 247052 322388 247104
rect 322440 247092 322446 247104
rect 506566 247092 506572 247104
rect 322440 247064 506572 247092
rect 322440 247052 322446 247064
rect 506566 247052 506572 247064
rect 506624 247052 506630 247104
rect 269114 246304 269120 246356
rect 269172 246344 269178 246356
rect 324130 246344 324136 246356
rect 269172 246316 324136 246344
rect 269172 246304 269178 246316
rect 324130 246304 324136 246316
rect 324188 246304 324194 246356
rect 309042 245760 309048 245812
rect 309100 245800 309106 245812
rect 346394 245800 346400 245812
rect 309100 245772 346400 245800
rect 309100 245760 309106 245772
rect 346394 245760 346400 245772
rect 346452 245760 346458 245812
rect 320358 245692 320364 245744
rect 320416 245732 320422 245744
rect 321278 245732 321284 245744
rect 320416 245704 321284 245732
rect 320416 245692 320422 245704
rect 321278 245692 321284 245704
rect 321336 245732 321342 245744
rect 491294 245732 491300 245744
rect 321336 245704 491300 245732
rect 321336 245692 321342 245704
rect 491294 245692 491300 245704
rect 491352 245692 491358 245744
rect 321186 245624 321192 245676
rect 321244 245664 321250 245676
rect 321462 245664 321468 245676
rect 321244 245636 321468 245664
rect 321244 245624 321250 245636
rect 321462 245624 321468 245636
rect 321520 245664 321526 245676
rect 499574 245664 499580 245676
rect 321520 245636 499580 245664
rect 321520 245624 321526 245636
rect 499574 245624 499580 245636
rect 499632 245624 499638 245676
rect 310790 245148 310796 245200
rect 310848 245188 310854 245200
rect 311250 245188 311256 245200
rect 310848 245160 311256 245188
rect 310848 245148 310854 245160
rect 311250 245148 311256 245160
rect 311308 245148 311314 245200
rect 268930 244944 268936 244996
rect 268988 244984 268994 244996
rect 284478 244984 284484 244996
rect 268988 244956 284484 244984
rect 268988 244944 268994 244956
rect 284478 244944 284484 244956
rect 284536 244944 284542 244996
rect 269206 244876 269212 244928
rect 269264 244916 269270 244928
rect 323670 244916 323676 244928
rect 269264 244888 323676 244916
rect 269264 244876 269270 244888
rect 323670 244876 323676 244888
rect 323728 244876 323734 244928
rect 311250 244332 311256 244384
rect 311308 244372 311314 244384
rect 371234 244372 371240 244384
rect 311308 244344 371240 244372
rect 311308 244332 311314 244344
rect 371234 244332 371240 244344
rect 371292 244332 371298 244384
rect 322474 244264 322480 244316
rect 322532 244304 322538 244316
rect 503714 244304 503720 244316
rect 322532 244276 503720 244304
rect 322532 244264 322538 244276
rect 503714 244264 503720 244276
rect 503772 244264 503778 244316
rect 269022 243516 269028 243568
rect 269080 243556 269086 243568
rect 325694 243556 325700 243568
rect 269080 243528 325700 243556
rect 269080 243516 269086 243528
rect 325694 243516 325700 243528
rect 325752 243516 325758 243568
rect 321370 242904 321376 242956
rect 321428 242944 321434 242956
rect 492674 242944 492680 242956
rect 321428 242916 492680 242944
rect 321428 242904 321434 242916
rect 492674 242904 492680 242916
rect 492732 242904 492738 242956
rect 242866 241556 248828 241584
rect 215754 241476 215760 241528
rect 215812 241516 215818 241528
rect 220998 241516 221004 241528
rect 215812 241488 221004 241516
rect 215812 241476 215818 241488
rect 220998 241476 221004 241488
rect 221056 241476 221062 241528
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 219986 241448 219992 241460
rect 3476 241420 219992 241448
rect 3476 241408 3482 241420
rect 219986 241408 219992 241420
rect 220044 241408 220050 241460
rect 223546 241148 235994 241176
rect 220354 241000 220360 241052
rect 220412 241040 220418 241052
rect 223546 241040 223574 241148
rect 220412 241012 223574 241040
rect 220412 241000 220418 241012
rect 218790 240932 218796 240984
rect 218848 240972 218854 240984
rect 218848 240944 222194 240972
rect 218848 240932 218854 240944
rect 202874 240864 202880 240916
rect 202932 240904 202938 240916
rect 220354 240904 220360 240916
rect 202932 240876 220360 240904
rect 202932 240864 202938 240876
rect 220354 240864 220360 240876
rect 220412 240864 220418 240916
rect 193214 240796 193220 240848
rect 193272 240836 193278 240848
rect 220170 240836 220176 240848
rect 193272 240808 220176 240836
rect 193272 240796 193278 240808
rect 220170 240796 220176 240808
rect 220228 240836 220234 240848
rect 222166 240836 222194 240944
rect 222286 240864 222292 240916
rect 222344 240904 222350 240916
rect 222344 240876 234614 240904
rect 222344 240864 222350 240876
rect 220228 240808 221320 240836
rect 222166 240808 230842 240836
rect 220228 240796 220234 240808
rect 161474 240728 161480 240780
rect 161532 240768 161538 240780
rect 218790 240768 218796 240780
rect 161532 240740 218796 240768
rect 161532 240728 161538 240740
rect 218790 240728 218796 240740
rect 218848 240728 218854 240780
rect 219250 240592 219256 240644
rect 219308 240632 219314 240644
rect 220814 240632 220820 240644
rect 219308 240604 220820 240632
rect 219308 240592 219314 240604
rect 220814 240592 220820 240604
rect 220872 240592 220878 240644
rect 221292 240632 221320 240808
rect 221366 240728 221372 240780
rect 221424 240768 221430 240780
rect 221826 240768 221832 240780
rect 221424 240740 221832 240768
rect 221424 240728 221430 240740
rect 221826 240728 221832 240740
rect 221884 240728 221890 240780
rect 221734 240660 221740 240712
rect 221792 240700 221798 240712
rect 221792 240672 228404 240700
rect 221792 240660 221798 240672
rect 222286 240632 222292 240644
rect 221292 240604 222292 240632
rect 222286 240592 222292 240604
rect 222344 240592 222350 240644
rect 228376 240632 228404 240672
rect 228376 240604 230750 240632
rect 214374 240456 214380 240508
rect 214432 240496 214438 240508
rect 218698 240496 218704 240508
rect 214432 240468 218704 240496
rect 214432 240456 214438 240468
rect 218698 240456 218704 240468
rect 218756 240456 218762 240508
rect 219158 240456 219164 240508
rect 219216 240496 219222 240508
rect 221182 240496 221188 240508
rect 219216 240468 221188 240496
rect 219216 240456 219222 240468
rect 221182 240456 221188 240468
rect 221240 240456 221246 240508
rect 223546 240468 227990 240496
rect 214466 240388 214472 240440
rect 214524 240428 214530 240440
rect 223546 240428 223574 240468
rect 214524 240400 223574 240428
rect 214524 240388 214530 240400
rect 215570 240320 215576 240372
rect 215628 240360 215634 240372
rect 227962 240360 227990 240468
rect 215628 240332 227070 240360
rect 227962 240332 230658 240360
rect 215628 240320 215634 240332
rect 217686 240252 217692 240304
rect 217744 240292 217750 240304
rect 221090 240292 221096 240304
rect 217744 240264 221096 240292
rect 217744 240252 217750 240264
rect 221090 240252 221096 240264
rect 221148 240252 221154 240304
rect 222286 240252 222292 240304
rect 222344 240292 222350 240304
rect 222344 240264 223114 240292
rect 222344 240252 222350 240264
rect 216214 240184 216220 240236
rect 216272 240224 216278 240236
rect 221734 240224 221740 240236
rect 216272 240196 221740 240224
rect 216272 240184 216278 240196
rect 221734 240184 221740 240196
rect 221792 240184 221798 240236
rect 223086 240224 223114 240264
rect 227042 240224 227070 240332
rect 223086 240196 224862 240224
rect 227042 240196 230566 240224
rect 210418 240048 210424 240100
rect 210476 240088 210482 240100
rect 219342 240088 219348 240100
rect 210476 240060 219348 240088
rect 210476 240048 210482 240060
rect 219342 240048 219348 240060
rect 219400 240048 219406 240100
rect 222194 240048 222200 240100
rect 222252 240088 222258 240100
rect 222252 240060 223574 240088
rect 222252 240048 222258 240060
rect 222286 239980 222292 240032
rect 222344 240020 222350 240032
rect 222344 239992 222930 240020
rect 222344 239980 222350 239992
rect 222902 239964 222930 239992
rect 207014 239912 207020 239964
rect 207072 239952 207078 239964
rect 213362 239952 213368 239964
rect 207072 239924 213368 239952
rect 207072 239912 207078 239924
rect 213362 239912 213368 239924
rect 213420 239952 213426 239964
rect 213420 239924 220814 239952
rect 213420 239912 213426 239924
rect 216306 239844 216312 239896
rect 216364 239884 216370 239896
rect 216582 239884 216588 239896
rect 216364 239856 216588 239884
rect 216364 239844 216370 239856
rect 216582 239844 216588 239856
rect 216640 239844 216646 239896
rect 219158 239844 219164 239896
rect 219216 239884 219222 239896
rect 219342 239884 219348 239896
rect 219216 239856 219348 239884
rect 219216 239844 219222 239856
rect 219342 239844 219348 239856
rect 219400 239844 219406 239896
rect 197354 239776 197360 239828
rect 197412 239816 197418 239828
rect 220262 239816 220268 239828
rect 197412 239788 220268 239816
rect 197412 239776 197418 239788
rect 220262 239776 220268 239788
rect 220320 239776 220326 239828
rect 220786 239816 220814 239924
rect 221918 239912 221924 239964
rect 221976 239952 221982 239964
rect 222378 239952 222384 239964
rect 221976 239924 222384 239952
rect 221976 239912 221982 239924
rect 222378 239912 222384 239924
rect 222436 239912 222442 239964
rect 222884 239912 222890 239964
rect 222942 239912 222948 239964
rect 223344 239912 223350 239964
rect 223402 239912 223408 239964
rect 223436 239912 223442 239964
rect 223494 239912 223500 239964
rect 220998 239844 221004 239896
rect 221056 239884 221062 239896
rect 221056 239856 222608 239884
rect 221056 239844 221062 239856
rect 221274 239816 221280 239828
rect 220786 239788 221280 239816
rect 221274 239776 221280 239788
rect 221332 239776 221338 239828
rect 222580 239816 222608 239856
rect 222700 239844 222706 239896
rect 222758 239844 222764 239896
rect 222792 239844 222798 239896
rect 222850 239844 222856 239896
rect 223160 239884 223166 239896
rect 223132 239844 223166 239884
rect 223218 239844 223224 239896
rect 223362 239884 223390 239912
rect 223316 239856 223390 239884
rect 222718 239816 222746 239844
rect 222580 239788 222746 239816
rect 222810 239760 222838 239844
rect 182174 239708 182180 239760
rect 182232 239748 182238 239760
rect 219158 239748 219164 239760
rect 182232 239720 219164 239748
rect 182232 239708 182238 239720
rect 219158 239708 219164 239720
rect 219216 239708 219222 239760
rect 219250 239708 219256 239760
rect 219308 239748 219314 239760
rect 222194 239748 222200 239760
rect 219308 239720 222200 239748
rect 219308 239708 219314 239720
rect 222194 239708 222200 239720
rect 222252 239708 222258 239760
rect 222746 239708 222752 239760
rect 222804 239720 222838 239760
rect 222804 239708 222810 239720
rect 223132 239692 223160 239844
rect 175274 239640 175280 239692
rect 175332 239680 175338 239692
rect 218974 239680 218980 239692
rect 175332 239652 218980 239680
rect 175332 239640 175338 239652
rect 218974 239640 218980 239652
rect 219032 239680 219038 239692
rect 219342 239680 219348 239692
rect 219032 239652 219348 239680
rect 219032 239640 219038 239652
rect 219342 239640 219348 239652
rect 219400 239640 219406 239692
rect 223114 239640 223120 239692
rect 223172 239640 223178 239692
rect 139394 239572 139400 239624
rect 139452 239612 139458 239624
rect 139452 239584 215892 239612
rect 139452 239572 139458 239584
rect 125594 239504 125600 239556
rect 125652 239544 125658 239556
rect 214374 239544 214380 239556
rect 125652 239516 214380 239544
rect 125652 239504 125658 239516
rect 214374 239504 214380 239516
rect 214432 239504 214438 239556
rect 103514 239436 103520 239488
rect 103572 239476 103578 239488
rect 214558 239476 214564 239488
rect 103572 239448 214564 239476
rect 103572 239436 103578 239448
rect 214558 239436 214564 239448
rect 214616 239476 214622 239488
rect 215570 239476 215576 239488
rect 214616 239448 215576 239476
rect 214616 239436 214622 239448
rect 215570 239436 215576 239448
rect 215628 239436 215634 239488
rect 215864 239476 215892 239584
rect 217962 239572 217968 239624
rect 218020 239612 218026 239624
rect 222286 239612 222292 239624
rect 218020 239584 222292 239612
rect 218020 239572 218026 239584
rect 222286 239572 222292 239584
rect 222344 239612 222350 239624
rect 223316 239612 223344 239856
rect 223454 239692 223482 239912
rect 223546 239828 223574 240060
rect 224834 239964 224862 240196
rect 226214 239992 227162 240020
rect 226214 239964 226242 239992
rect 223712 239912 223718 239964
rect 223770 239952 223776 239964
rect 224540 239952 224546 239964
rect 223770 239912 223804 239952
rect 223528 239776 223534 239828
rect 223586 239776 223592 239828
rect 223390 239640 223396 239692
rect 223448 239652 223482 239692
rect 223448 239640 223454 239652
rect 223574 239640 223580 239692
rect 223632 239680 223638 239692
rect 223776 239680 223804 239912
rect 224190 239924 224546 239952
rect 223896 239844 223902 239896
rect 223954 239844 223960 239896
rect 223988 239844 223994 239896
rect 224046 239844 224052 239896
rect 223914 239816 223942 239844
rect 223868 239788 223942 239816
rect 223868 239692 223896 239788
rect 223632 239652 223804 239680
rect 223632 239640 223638 239652
rect 223850 239640 223856 239692
rect 223908 239640 223914 239692
rect 222344 239584 223344 239612
rect 222344 239572 222350 239584
rect 223482 239572 223488 239624
rect 223540 239612 223546 239624
rect 224006 239612 224034 239844
rect 223540 239584 224034 239612
rect 224190 239624 224218 239924
rect 224540 239912 224546 239924
rect 224598 239912 224604 239964
rect 224632 239912 224638 239964
rect 224690 239912 224696 239964
rect 224724 239912 224730 239964
rect 224782 239912 224788 239964
rect 224816 239912 224822 239964
rect 224874 239912 224880 239964
rect 225000 239912 225006 239964
rect 225058 239952 225064 239964
rect 225276 239952 225282 239964
rect 225058 239924 225184 239952
rect 225058 239912 225064 239924
rect 224264 239844 224270 239896
rect 224322 239844 224328 239896
rect 224356 239844 224362 239896
rect 224414 239844 224420 239896
rect 224282 239760 224310 239844
rect 224374 239816 224402 239844
rect 224650 239828 224678 239912
rect 224742 239828 224770 239912
rect 224374 239788 224540 239816
rect 224282 239720 224316 239760
rect 224310 239708 224316 239720
rect 224368 239708 224374 239760
rect 224512 239624 224540 239788
rect 224586 239776 224592 239828
rect 224644 239788 224678 239828
rect 224644 239776 224650 239788
rect 224724 239776 224730 239828
rect 224782 239776 224788 239828
rect 225156 239760 225184 239924
rect 225248 239912 225282 239952
rect 225334 239912 225340 239964
rect 225368 239912 225374 239964
rect 225426 239912 225432 239964
rect 225552 239952 225558 239964
rect 225524 239912 225558 239952
rect 225610 239912 225616 239964
rect 225644 239912 225650 239964
rect 225702 239912 225708 239964
rect 226196 239912 226202 239964
rect 226254 239912 226260 239964
rect 226932 239912 226938 239964
rect 226990 239912 226996 239964
rect 227024 239912 227030 239964
rect 227082 239912 227088 239964
rect 225138 239708 225144 239760
rect 225196 239708 225202 239760
rect 225248 239692 225276 239912
rect 225386 239884 225414 239912
rect 225340 239856 225414 239884
rect 225230 239640 225236 239692
rect 225288 239640 225294 239692
rect 225340 239624 225368 239856
rect 225524 239624 225552 239912
rect 225662 239828 225690 239912
rect 226104 239844 226110 239896
rect 226162 239844 226168 239896
rect 226564 239884 226570 239896
rect 226536 239844 226570 239884
rect 226622 239844 226628 239896
rect 226656 239844 226662 239896
rect 226714 239844 226720 239896
rect 226748 239844 226754 239896
rect 226806 239844 226812 239896
rect 225598 239776 225604 239828
rect 225656 239788 225690 239828
rect 225656 239776 225662 239788
rect 226122 239624 226150 239844
rect 224190 239584 224224 239624
rect 223540 239572 223546 239584
rect 224218 239572 224224 239584
rect 224276 239572 224282 239624
rect 224494 239572 224500 239624
rect 224552 239572 224558 239624
rect 224770 239572 224776 239624
rect 224828 239612 224834 239624
rect 225322 239612 225328 239624
rect 224828 239584 225328 239612
rect 224828 239572 224834 239584
rect 225322 239572 225328 239584
rect 225380 239572 225386 239624
rect 225506 239572 225512 239624
rect 225564 239572 225570 239624
rect 226058 239572 226064 239624
rect 226116 239584 226150 239624
rect 226536 239612 226564 239844
rect 226674 239692 226702 239844
rect 226610 239640 226616 239692
rect 226668 239652 226702 239692
rect 226766 239692 226794 239844
rect 226950 239760 226978 239912
rect 226886 239708 226892 239760
rect 226944 239720 226978 239760
rect 226944 239708 226950 239720
rect 226766 239652 226800 239692
rect 226668 239640 226674 239652
rect 226794 239640 226800 239652
rect 226852 239640 226858 239692
rect 226702 239612 226708 239624
rect 226536 239584 226708 239612
rect 226116 239572 226122 239584
rect 226702 239572 226708 239584
rect 226760 239572 226766 239624
rect 226886 239572 226892 239624
rect 226944 239612 226950 239624
rect 227042 239612 227070 239912
rect 227134 239760 227162 239992
rect 230538 239964 230566 240196
rect 227392 239952 227398 239964
rect 227318 239924 227398 239952
rect 227208 239844 227214 239896
rect 227266 239844 227272 239896
rect 227116 239708 227122 239760
rect 227174 239708 227180 239760
rect 227226 239612 227254 239844
rect 227318 239692 227346 239924
rect 227392 239912 227398 239924
rect 227450 239912 227456 239964
rect 227760 239912 227766 239964
rect 227818 239912 227824 239964
rect 228128 239912 228134 239964
rect 228186 239912 228192 239964
rect 228238 239924 228496 239952
rect 227484 239844 227490 239896
rect 227542 239844 227548 239896
rect 227576 239844 227582 239896
rect 227634 239884 227640 239896
rect 227634 239856 227714 239884
rect 227634 239844 227640 239856
rect 227502 239816 227530 239844
rect 227502 239788 227576 239816
rect 227548 239760 227576 239788
rect 227530 239708 227536 239760
rect 227588 239708 227594 239760
rect 227318 239652 227352 239692
rect 227346 239640 227352 239652
rect 227404 239640 227410 239692
rect 227686 239680 227714 239856
rect 227640 239652 227714 239680
rect 226944 239584 227070 239612
rect 227180 239584 227254 239612
rect 226944 239572 226950 239584
rect 227180 239556 227208 239584
rect 215938 239504 215944 239556
rect 215996 239544 216002 239556
rect 227070 239544 227076 239556
rect 215996 239516 227076 239544
rect 215996 239504 216002 239516
rect 227070 239504 227076 239516
rect 227128 239504 227134 239556
rect 227162 239504 227168 239556
rect 227220 239504 227226 239556
rect 227254 239504 227260 239556
rect 227312 239544 227318 239556
rect 227640 239544 227668 239652
rect 227778 239624 227806 239912
rect 228036 239844 228042 239896
rect 228094 239844 228100 239896
rect 227714 239572 227720 239624
rect 227772 239584 227806 239624
rect 227772 239572 227778 239584
rect 227312 239516 227668 239544
rect 228054 239544 228082 239844
rect 228146 239692 228174 239912
rect 228238 239896 228266 239924
rect 228220 239844 228226 239896
rect 228278 239844 228284 239896
rect 228146 239652 228180 239692
rect 228174 239640 228180 239652
rect 228232 239640 228238 239692
rect 228468 239612 228496 239924
rect 228680 239912 228686 239964
rect 228738 239912 228744 239964
rect 228864 239912 228870 239964
rect 228922 239912 228928 239964
rect 228956 239912 228962 239964
rect 229014 239912 229020 239964
rect 229968 239912 229974 239964
rect 230026 239912 230032 239964
rect 230244 239912 230250 239964
rect 230302 239912 230308 239964
rect 230520 239912 230526 239964
rect 230578 239912 230584 239964
rect 228588 239884 228594 239896
rect 228560 239844 228594 239884
rect 228646 239844 228652 239896
rect 228560 239760 228588 239844
rect 228542 239708 228548 239760
rect 228600 239708 228606 239760
rect 228698 239680 228726 239912
rect 228882 239760 228910 239912
rect 228818 239708 228824 239760
rect 228876 239720 228910 239760
rect 228974 239760 229002 239912
rect 229048 239844 229054 239896
rect 229106 239844 229112 239896
rect 229600 239844 229606 239896
rect 229658 239844 229664 239896
rect 229066 239816 229094 239844
rect 229066 239788 229140 239816
rect 228974 239720 229008 239760
rect 228876 239708 228882 239720
rect 229002 239708 229008 239720
rect 229060 239708 229066 239760
rect 228652 239652 228726 239680
rect 228652 239624 228680 239652
rect 228376 239584 228496 239612
rect 228376 239556 228404 239584
rect 228634 239572 228640 239624
rect 228692 239572 228698 239624
rect 228726 239572 228732 239624
rect 228784 239612 228790 239624
rect 229112 239612 229140 239788
rect 228784 239584 229140 239612
rect 228784 239572 228790 239584
rect 229186 239572 229192 239624
rect 229244 239612 229250 239624
rect 229618 239612 229646 239844
rect 229986 239760 230014 239912
rect 230060 239844 230066 239896
rect 230118 239884 230124 239896
rect 230118 239844 230152 239884
rect 230124 239760 230152 239844
rect 230262 239760 230290 239912
rect 230336 239844 230342 239896
rect 230394 239844 230400 239896
rect 230354 239816 230382 239844
rect 230354 239788 230428 239816
rect 230400 239760 230428 239788
rect 229986 239720 230020 239760
rect 230014 239708 230020 239720
rect 230072 239708 230078 239760
rect 230106 239708 230112 239760
rect 230164 239708 230170 239760
rect 230262 239720 230296 239760
rect 230290 239708 230296 239720
rect 230348 239708 230354 239760
rect 230382 239708 230388 239760
rect 230440 239708 230446 239760
rect 229244 239584 229646 239612
rect 229244 239572 229250 239584
rect 230382 239572 230388 239624
rect 230440 239612 230446 239624
rect 230630 239612 230658 240332
rect 230722 240020 230750 240604
rect 230814 240088 230842 240808
rect 234586 240428 234614 240876
rect 235966 240496 235994 241148
rect 235966 240468 237650 240496
rect 234586 240400 235994 240428
rect 235966 240224 235994 240400
rect 235966 240196 237558 240224
rect 230814 240060 235074 240088
rect 230722 239992 234660 240020
rect 230796 239912 230802 239964
rect 230854 239952 230860 239964
rect 230854 239924 231072 239952
rect 230854 239912 230860 239924
rect 230888 239844 230894 239896
rect 230946 239844 230952 239896
rect 230440 239584 230658 239612
rect 230440 239572 230446 239584
rect 230750 239572 230756 239624
rect 230808 239612 230814 239624
rect 230906 239612 230934 239844
rect 231044 239624 231072 239924
rect 231256 239912 231262 239964
rect 231314 239912 231320 239964
rect 231348 239912 231354 239964
rect 231406 239912 231412 239964
rect 231440 239912 231446 239964
rect 231498 239912 231504 239964
rect 231624 239912 231630 239964
rect 231682 239912 231688 239964
rect 232452 239912 232458 239964
rect 232510 239952 232516 239964
rect 232510 239924 232636 239952
rect 232510 239912 232516 239924
rect 231274 239624 231302 239912
rect 231366 239680 231394 239912
rect 231458 239760 231486 239912
rect 231642 239760 231670 239912
rect 231808 239844 231814 239896
rect 231866 239844 231872 239896
rect 231900 239844 231906 239896
rect 231958 239844 231964 239896
rect 232084 239844 232090 239896
rect 232142 239844 232148 239896
rect 231826 239760 231854 239844
rect 231458 239720 231492 239760
rect 231486 239708 231492 239720
rect 231544 239708 231550 239760
rect 231578 239708 231584 239760
rect 231636 239720 231670 239760
rect 231636 239708 231642 239720
rect 231762 239708 231768 239760
rect 231820 239720 231854 239760
rect 231820 239708 231826 239720
rect 231918 239680 231946 239844
rect 232102 239748 232130 239844
rect 232102 239720 232176 239748
rect 231366 239652 231854 239680
rect 231918 239652 232084 239680
rect 230808 239584 230934 239612
rect 230808 239572 230814 239584
rect 231026 239572 231032 239624
rect 231084 239572 231090 239624
rect 231274 239572 231308 239624
rect 231360 239572 231366 239624
rect 231826 239612 231854 239652
rect 231946 239612 231952 239624
rect 231826 239584 231952 239612
rect 231946 239572 231952 239584
rect 232004 239572 232010 239624
rect 228174 239544 228180 239556
rect 228054 239516 228180 239544
rect 227312 239504 227318 239516
rect 228174 239504 228180 239516
rect 228232 239504 228238 239556
rect 228358 239504 228364 239556
rect 228416 239504 228422 239556
rect 230566 239504 230572 239556
rect 230624 239544 230630 239556
rect 231274 239544 231302 239572
rect 230624 239516 231302 239544
rect 232056 239544 232084 239652
rect 232148 239624 232176 239720
rect 232608 239692 232636 239924
rect 232728 239912 232734 239964
rect 232786 239912 232792 239964
rect 232820 239912 232826 239964
rect 232878 239912 232884 239964
rect 233004 239952 233010 239964
rect 232976 239912 233010 239952
rect 233062 239912 233068 239964
rect 233188 239952 233194 239964
rect 233160 239912 233194 239952
rect 233246 239912 233252 239964
rect 233280 239912 233286 239964
rect 233338 239912 233344 239964
rect 233464 239912 233470 239964
rect 233522 239912 233528 239964
rect 233832 239912 233838 239964
rect 233890 239912 233896 239964
rect 234016 239912 234022 239964
rect 234074 239912 234080 239964
rect 234384 239912 234390 239964
rect 234442 239912 234448 239964
rect 232746 239884 232774 239912
rect 232700 239856 232774 239884
rect 232590 239640 232596 239692
rect 232648 239640 232654 239692
rect 232700 239624 232728 239856
rect 232838 239828 232866 239912
rect 232774 239776 232780 239828
rect 232832 239788 232866 239828
rect 232832 239776 232838 239788
rect 232976 239760 233004 239912
rect 232958 239708 232964 239760
rect 233016 239708 233022 239760
rect 233160 239692 233188 239912
rect 233142 239640 233148 239692
rect 233200 239640 233206 239692
rect 232130 239572 232136 239624
rect 232188 239572 232194 239624
rect 232682 239572 232688 239624
rect 232740 239572 232746 239624
rect 232222 239544 232228 239556
rect 232056 239516 232228 239544
rect 230624 239504 230630 239516
rect 232222 239504 232228 239516
rect 232280 239504 232286 239556
rect 220630 239476 220636 239488
rect 215864 239448 220636 239476
rect 220630 239436 220636 239448
rect 220688 239476 220694 239488
rect 233298 239476 233326 239912
rect 233482 239624 233510 239912
rect 233740 239844 233746 239896
rect 233798 239844 233804 239896
rect 233758 239760 233786 239844
rect 233850 239816 233878 239912
rect 233850 239788 233924 239816
rect 233694 239708 233700 239760
rect 233752 239720 233786 239760
rect 233752 239708 233758 239720
rect 233896 239680 233924 239788
rect 233712 239652 233924 239680
rect 233482 239584 233516 239624
rect 233510 239572 233516 239584
rect 233568 239572 233574 239624
rect 233712 239544 233740 239652
rect 233786 239572 233792 239624
rect 233844 239612 233850 239624
rect 234034 239612 234062 239912
rect 234402 239692 234430 239912
rect 234338 239640 234344 239692
rect 234396 239652 234430 239692
rect 234396 239640 234402 239652
rect 234632 239624 234660 239992
rect 235046 239964 235074 240060
rect 237530 239964 237558 240196
rect 237622 240088 237650 240468
rect 242866 240156 242894 241556
rect 240750 240128 242894 240156
rect 237622 240060 238294 240088
rect 238266 239964 238294 240060
rect 239278 239992 239858 240020
rect 234844 239912 234850 239964
rect 234902 239912 234908 239964
rect 235028 239912 235034 239964
rect 235086 239912 235092 239964
rect 235304 239912 235310 239964
rect 235362 239912 235368 239964
rect 235488 239912 235494 239964
rect 235546 239912 235552 239964
rect 235856 239912 235862 239964
rect 235914 239912 235920 239964
rect 236040 239912 236046 239964
rect 236098 239952 236104 239964
rect 236224 239952 236230 239964
rect 236098 239912 236132 239952
rect 234862 239760 234890 239912
rect 235212 239844 235218 239896
rect 235270 239844 235276 239896
rect 235230 239760 235258 239844
rect 234862 239720 234896 239760
rect 234890 239708 234896 239720
rect 234948 239708 234954 239760
rect 235166 239708 235172 239760
rect 235224 239720 235258 239760
rect 235224 239708 235230 239720
rect 235322 239692 235350 239912
rect 235258 239640 235264 239692
rect 235316 239652 235350 239692
rect 235316 239640 235322 239652
rect 233844 239584 234062 239612
rect 233844 239572 233850 239584
rect 234614 239572 234620 239624
rect 234672 239572 234678 239624
rect 235506 239556 235534 239912
rect 235764 239844 235770 239896
rect 235822 239844 235828 239896
rect 235782 239692 235810 239844
rect 235874 239760 235902 239912
rect 235874 239720 235908 239760
rect 235902 239708 235908 239720
rect 235960 239708 235966 239760
rect 235782 239652 235816 239692
rect 235810 239640 235816 239652
rect 235868 239640 235874 239692
rect 233970 239544 233976 239556
rect 233712 239516 233976 239544
rect 233970 239504 233976 239516
rect 234028 239504 234034 239556
rect 235442 239504 235448 239556
rect 235500 239516 235534 239556
rect 235500 239504 235506 239516
rect 220688 239448 233326 239476
rect 220688 239436 220694 239448
rect 3418 239368 3424 239420
rect 3476 239408 3482 239420
rect 217226 239408 217232 239420
rect 3476 239380 217232 239408
rect 3476 239368 3482 239380
rect 217226 239368 217232 239380
rect 217284 239368 217290 239420
rect 218698 239368 218704 239420
rect 218756 239408 218762 239420
rect 219066 239408 219072 239420
rect 218756 239380 219072 239408
rect 218756 239368 218762 239380
rect 219066 239368 219072 239380
rect 219124 239368 219130 239420
rect 219342 239368 219348 239420
rect 219400 239408 219406 239420
rect 236104 239408 236132 239912
rect 236196 239912 236230 239952
rect 236282 239912 236288 239964
rect 236316 239912 236322 239964
rect 236374 239912 236380 239964
rect 236684 239912 236690 239964
rect 236742 239912 236748 239964
rect 236776 239912 236782 239964
rect 236834 239912 236840 239964
rect 237236 239912 237242 239964
rect 237294 239912 237300 239964
rect 237512 239912 237518 239964
rect 237570 239912 237576 239964
rect 237788 239912 237794 239964
rect 237846 239952 237852 239964
rect 237846 239912 237880 239952
rect 237972 239912 237978 239964
rect 238030 239912 238036 239964
rect 238064 239912 238070 239964
rect 238122 239912 238128 239964
rect 238248 239912 238254 239964
rect 238306 239912 238312 239964
rect 239076 239912 239082 239964
rect 239134 239912 239140 239964
rect 236196 239556 236224 239912
rect 236178 239504 236184 239556
rect 236236 239504 236242 239556
rect 219400 239380 236132 239408
rect 219400 239368 219406 239380
rect 178034 239300 178040 239352
rect 178092 239340 178098 239352
rect 236334 239340 236362 239912
rect 236500 239844 236506 239896
rect 236558 239844 236564 239896
rect 236518 239760 236546 239844
rect 236518 239720 236552 239760
rect 236546 239708 236552 239720
rect 236604 239708 236610 239760
rect 236702 239680 236730 239912
rect 236472 239652 236730 239680
rect 236472 239544 236500 239652
rect 236546 239572 236552 239624
rect 236604 239612 236610 239624
rect 236794 239612 236822 239912
rect 237052 239844 237058 239896
rect 237110 239844 237116 239896
rect 237070 239760 237098 239844
rect 237006 239708 237012 239760
rect 237064 239720 237098 239760
rect 237064 239708 237070 239720
rect 236604 239584 236822 239612
rect 237254 239624 237282 239912
rect 237742 239816 237748 239828
rect 237668 239788 237748 239816
rect 237668 239692 237696 239788
rect 237742 239776 237748 239788
rect 237800 239776 237806 239828
rect 237650 239640 237656 239692
rect 237708 239640 237714 239692
rect 237742 239640 237748 239692
rect 237800 239680 237806 239692
rect 237852 239680 237880 239912
rect 237800 239652 237880 239680
rect 237800 239640 237806 239652
rect 237990 239624 238018 239912
rect 238082 239748 238110 239912
rect 238800 239844 238806 239896
rect 238858 239844 238864 239896
rect 238892 239844 238898 239896
rect 238950 239844 238956 239896
rect 239094 239884 239122 239912
rect 239048 239856 239122 239884
rect 238524 239776 238530 239828
rect 238582 239776 238588 239828
rect 238082 239720 238248 239748
rect 237254 239584 237288 239624
rect 236604 239572 236610 239584
rect 237282 239572 237288 239584
rect 237340 239572 237346 239624
rect 237990 239584 238024 239624
rect 238018 239572 238024 239584
rect 238076 239572 238082 239624
rect 236730 239544 236736 239556
rect 236472 239516 236736 239544
rect 236730 239504 236736 239516
rect 236788 239504 236794 239556
rect 238220 239544 238248 239720
rect 238542 239556 238570 239776
rect 238818 239624 238846 239844
rect 238910 239692 238938 239844
rect 238910 239652 238944 239692
rect 238938 239640 238944 239652
rect 238996 239640 239002 239692
rect 238754 239572 238760 239624
rect 238812 239584 238846 239624
rect 238812 239572 238818 239584
rect 238386 239544 238392 239556
rect 238220 239516 238392 239544
rect 238386 239504 238392 239516
rect 238444 239504 238450 239556
rect 238478 239504 238484 239556
rect 238536 239516 238570 239556
rect 238536 239504 238542 239516
rect 238846 239504 238852 239556
rect 238904 239544 238910 239556
rect 239048 239544 239076 239856
rect 239168 239844 239174 239896
rect 239226 239844 239232 239896
rect 239186 239816 239214 239844
rect 239140 239788 239214 239816
rect 239140 239760 239168 239788
rect 239278 239760 239306 239992
rect 239830 239964 239858 239992
rect 240750 239964 240778 240128
rect 241026 239992 242066 240020
rect 239444 239912 239450 239964
rect 239502 239912 239508 239964
rect 239536 239912 239542 239964
rect 239594 239952 239600 239964
rect 239594 239912 239628 239952
rect 239720 239912 239726 239964
rect 239778 239912 239784 239964
rect 239812 239912 239818 239964
rect 239870 239912 239876 239964
rect 239996 239952 240002 239964
rect 239968 239912 240002 239952
rect 240054 239912 240060 239964
rect 240180 239912 240186 239964
rect 240238 239912 240244 239964
rect 240732 239912 240738 239964
rect 240790 239912 240796 239964
rect 240916 239912 240922 239964
rect 240974 239912 240980 239964
rect 239352 239844 239358 239896
rect 239410 239844 239416 239896
rect 239122 239708 239128 239760
rect 239180 239708 239186 239760
rect 239214 239708 239220 239760
rect 239272 239720 239306 239760
rect 239272 239708 239278 239720
rect 239370 239612 239398 239844
rect 239462 239828 239490 239912
rect 239462 239788 239496 239828
rect 239490 239776 239496 239788
rect 239548 239776 239554 239828
rect 239600 239680 239628 239912
rect 239738 239828 239766 239912
rect 239738 239788 239772 239828
rect 239766 239776 239772 239788
rect 239824 239776 239830 239828
rect 239968 239760 239996 239912
rect 240088 239884 240094 239896
rect 240060 239844 240094 239884
rect 240146 239844 240152 239896
rect 239950 239708 239956 239760
rect 240008 239708 240014 239760
rect 240060 239692 240088 239844
rect 240198 239760 240226 239912
rect 240272 239844 240278 239896
rect 240330 239844 240336 239896
rect 240134 239708 240140 239760
rect 240192 239720 240226 239760
rect 240192 239708 240198 239720
rect 240290 239692 240318 239844
rect 240686 239708 240692 239760
rect 240744 239748 240750 239760
rect 240934 239748 240962 239912
rect 240744 239720 240962 239748
rect 240744 239708 240750 239720
rect 239508 239652 239628 239680
rect 239508 239624 239536 239652
rect 240042 239640 240048 239692
rect 240100 239640 240106 239692
rect 240226 239640 240232 239692
rect 240284 239652 240318 239692
rect 240284 239640 240290 239652
rect 239370 239584 239444 239612
rect 239416 239556 239444 239584
rect 239490 239572 239496 239624
rect 239548 239572 239554 239624
rect 238904 239516 239076 239544
rect 238904 239504 238910 239516
rect 239398 239504 239404 239556
rect 239456 239504 239462 239556
rect 236454 239436 236460 239488
rect 236512 239476 236518 239488
rect 241026 239476 241054 239992
rect 242038 239964 242066 239992
rect 241192 239912 241198 239964
rect 241250 239952 241256 239964
rect 241250 239924 241422 239952
rect 241250 239912 241256 239924
rect 241284 239844 241290 239896
rect 241342 239844 241348 239896
rect 241302 239760 241330 239844
rect 241238 239708 241244 239760
rect 241296 239720 241330 239760
rect 241296 239708 241302 239720
rect 241146 239572 241152 239624
rect 241204 239612 241210 239624
rect 241394 239612 241422 239924
rect 241468 239912 241474 239964
rect 241526 239912 241532 239964
rect 241928 239912 241934 239964
rect 241986 239912 241992 239964
rect 242020 239912 242026 239964
rect 242078 239912 242084 239964
rect 241204 239584 241422 239612
rect 241204 239572 241210 239584
rect 241330 239504 241336 239556
rect 241388 239544 241394 239556
rect 241486 239544 241514 239912
rect 241836 239844 241842 239896
rect 241894 239844 241900 239896
rect 241854 239816 241882 239844
rect 241624 239788 241882 239816
rect 241624 239556 241652 239788
rect 241946 239692 241974 239912
rect 241882 239640 241888 239692
rect 241940 239652 241974 239692
rect 241940 239640 241946 239652
rect 242176 239624 242204 240128
rect 245902 239992 246298 240020
rect 242296 239912 242302 239964
rect 242354 239912 242360 239964
rect 242388 239912 242394 239964
rect 242446 239912 242452 239964
rect 242572 239912 242578 239964
rect 242630 239912 242636 239964
rect 243400 239952 243406 239964
rect 243372 239912 243406 239952
rect 243458 239912 243464 239964
rect 243492 239912 243498 239964
rect 243550 239912 243556 239964
rect 243952 239912 243958 239964
rect 244010 239912 244016 239964
rect 244320 239912 244326 239964
rect 244378 239912 244384 239964
rect 244504 239912 244510 239964
rect 244562 239912 244568 239964
rect 244596 239912 244602 239964
rect 244654 239912 244660 239964
rect 245056 239912 245062 239964
rect 245114 239952 245120 239964
rect 245114 239924 245240 239952
rect 245114 239912 245120 239924
rect 242314 239680 242342 239912
rect 242406 239760 242434 239912
rect 242590 239884 242618 239912
rect 242590 239856 242848 239884
rect 242406 239720 242440 239760
rect 242434 239708 242440 239720
rect 242492 239708 242498 239760
rect 242526 239680 242532 239692
rect 242314 239652 242532 239680
rect 242526 239640 242532 239652
rect 242584 239640 242590 239692
rect 242820 239624 242848 239856
rect 242940 239844 242946 239896
rect 242998 239844 243004 239896
rect 243216 239844 243222 239896
rect 243274 239844 243280 239896
rect 242958 239760 242986 239844
rect 242958 239720 242992 239760
rect 242986 239708 242992 239720
rect 243044 239708 243050 239760
rect 242158 239572 242164 239624
rect 242216 239572 242222 239624
rect 242802 239572 242808 239624
rect 242860 239572 242866 239624
rect 241388 239516 241514 239544
rect 241388 239504 241394 239516
rect 241606 239504 241612 239556
rect 241664 239504 241670 239556
rect 236512 239448 241054 239476
rect 236512 239436 236518 239448
rect 242526 239436 242532 239488
rect 242584 239476 242590 239488
rect 242710 239476 242716 239488
rect 242584 239448 242716 239476
rect 242584 239436 242590 239448
rect 242710 239436 242716 239448
rect 242768 239436 242774 239488
rect 242986 239436 242992 239488
rect 243044 239476 243050 239488
rect 243234 239476 243262 239844
rect 243372 239624 243400 239912
rect 243510 239828 243538 239912
rect 243446 239776 243452 239828
rect 243504 239788 243538 239828
rect 243504 239776 243510 239788
rect 243970 239680 243998 239912
rect 244136 239844 244142 239896
rect 244194 239844 244200 239896
rect 244154 239816 244182 239844
rect 244154 239788 244228 239816
rect 244200 239692 244228 239788
rect 244338 239760 244366 239912
rect 244338 239720 244372 239760
rect 244366 239708 244372 239720
rect 244424 239708 244430 239760
rect 244090 239680 244096 239692
rect 243970 239652 244096 239680
rect 244090 239640 244096 239652
rect 244148 239640 244154 239692
rect 244182 239640 244188 239692
rect 244240 239640 244246 239692
rect 243354 239572 243360 239624
rect 243412 239572 243418 239624
rect 243044 239448 243262 239476
rect 243044 239436 243050 239448
rect 244522 239408 244550 239912
rect 244614 239476 244642 239912
rect 244688 239844 244694 239896
rect 244746 239844 244752 239896
rect 244872 239844 244878 239896
rect 244930 239844 244936 239896
rect 244706 239624 244734 239844
rect 244890 239760 244918 239844
rect 244890 239720 244924 239760
rect 244918 239708 244924 239720
rect 244976 239708 244982 239760
rect 245212 239692 245240 239924
rect 245332 239912 245338 239964
rect 245390 239912 245396 239964
rect 245424 239912 245430 239964
rect 245482 239912 245488 239964
rect 245516 239912 245522 239964
rect 245574 239912 245580 239964
rect 245700 239912 245706 239964
rect 245758 239912 245764 239964
rect 245350 239884 245378 239912
rect 245304 239856 245378 239884
rect 245194 239640 245200 239692
rect 245252 239640 245258 239692
rect 244706 239584 244740 239624
rect 244734 239572 244740 239584
rect 244792 239572 244798 239624
rect 245304 239612 245332 239856
rect 245442 239828 245470 239912
rect 245378 239776 245384 239828
rect 245436 239788 245470 239828
rect 245436 239776 245442 239788
rect 245534 239692 245562 239912
rect 245718 239692 245746 239912
rect 245534 239652 245568 239692
rect 245562 239640 245568 239652
rect 245620 239640 245626 239692
rect 245654 239640 245660 239692
rect 245712 239652 245746 239692
rect 245712 239640 245718 239652
rect 245212 239584 245332 239612
rect 245902 239612 245930 239992
rect 246270 239964 246298 239992
rect 246160 239912 246166 239964
rect 246218 239912 246224 239964
rect 246252 239912 246258 239964
rect 246310 239912 246316 239964
rect 246344 239912 246350 239964
rect 246402 239912 246408 239964
rect 246528 239912 246534 239964
rect 246586 239912 246592 239964
rect 246804 239912 246810 239964
rect 246862 239912 246868 239964
rect 246896 239912 246902 239964
rect 246954 239912 246960 239964
rect 247172 239912 247178 239964
rect 247230 239912 247236 239964
rect 247356 239912 247362 239964
rect 247414 239912 247420 239964
rect 247540 239912 247546 239964
rect 247598 239912 247604 239964
rect 248000 239912 248006 239964
rect 248058 239912 248064 239964
rect 248092 239912 248098 239964
rect 248150 239912 248156 239964
rect 248460 239912 248466 239964
rect 248518 239912 248524 239964
rect 248644 239912 248650 239964
rect 248702 239912 248708 239964
rect 245976 239844 245982 239896
rect 246034 239884 246040 239896
rect 246178 239884 246206 239912
rect 246034 239844 246068 239884
rect 246178 239856 246252 239884
rect 246040 239692 246068 239844
rect 246224 239828 246252 239856
rect 246206 239776 246212 239828
rect 246264 239776 246270 239828
rect 246022 239640 246028 239692
rect 246080 239640 246086 239692
rect 246206 239612 246212 239624
rect 245902 239584 246212 239612
rect 245212 239556 245240 239584
rect 246206 239572 246212 239584
rect 246264 239572 246270 239624
rect 245194 239504 245200 239556
rect 245252 239504 245258 239556
rect 245930 239476 245936 239488
rect 244614 239448 245936 239476
rect 245930 239436 245936 239448
rect 245988 239436 245994 239488
rect 244642 239408 244648 239420
rect 244522 239380 244648 239408
rect 244642 239368 244648 239380
rect 244700 239368 244706 239420
rect 246362 239408 246390 239912
rect 246546 239624 246574 239912
rect 246482 239572 246488 239624
rect 246540 239584 246574 239624
rect 246540 239572 246546 239584
rect 246666 239572 246672 239624
rect 246724 239612 246730 239624
rect 246822 239612 246850 239912
rect 246724 239584 246850 239612
rect 246724 239572 246730 239584
rect 246914 239556 246942 239912
rect 247034 239640 247040 239692
rect 247092 239680 247098 239692
rect 247190 239680 247218 239912
rect 247092 239652 247218 239680
rect 247092 239640 247098 239652
rect 247374 239624 247402 239912
rect 247558 239748 247586 239912
rect 248018 239760 248046 239912
rect 247862 239748 247868 239760
rect 247558 239720 247868 239748
rect 247862 239708 247868 239720
rect 247920 239708 247926 239760
rect 247954 239708 247960 239760
rect 248012 239720 248046 239760
rect 248012 239708 248018 239720
rect 248110 239624 248138 239912
rect 247374 239584 247408 239624
rect 247402 239572 247408 239584
rect 247460 239572 247466 239624
rect 248046 239572 248052 239624
rect 248104 239584 248138 239624
rect 248104 239572 248110 239584
rect 246850 239504 246856 239556
rect 246908 239516 246942 239556
rect 246908 239504 246914 239516
rect 248322 239436 248328 239488
rect 248380 239476 248386 239488
rect 248478 239476 248506 239912
rect 248662 239760 248690 239912
rect 248598 239708 248604 239760
rect 248656 239720 248690 239760
rect 248656 239708 248662 239720
rect 248800 239544 248828 241556
rect 259426 241420 260834 241448
rect 259426 241380 259454 241420
rect 249398 241352 259454 241380
rect 260806 241380 260834 241420
rect 260806 241352 264974 241380
rect 249168 239992 249334 240020
rect 248920 239952 248926 239964
rect 248892 239912 248926 239952
rect 248978 239912 248984 239964
rect 249012 239912 249018 239964
rect 249070 239912 249076 239964
rect 248892 239624 248920 239912
rect 249030 239828 249058 239912
rect 248966 239776 248972 239828
rect 249024 239788 249058 239828
rect 249024 239776 249030 239788
rect 248874 239572 248880 239624
rect 248932 239572 248938 239624
rect 249168 239544 249196 239992
rect 249306 239964 249334 239992
rect 249398 239964 249426 241352
rect 264946 241312 264974 241352
rect 267458 241312 267464 241324
rect 259426 241284 260834 241312
rect 264946 241284 267464 241312
rect 259426 240564 259454 241284
rect 260806 241176 260834 241284
rect 267458 241272 267464 241284
rect 267516 241272 267522 241324
rect 268102 241312 268108 241324
rect 267568 241284 268108 241312
rect 267568 241244 267596 241284
rect 268102 241272 268108 241284
rect 268160 241272 268166 241324
rect 264946 241216 267596 241244
rect 264946 241176 264974 241216
rect 267642 241204 267648 241256
rect 267700 241244 267706 241256
rect 268194 241244 268200 241256
rect 267700 241216 268200 241244
rect 267700 241204 267706 241216
rect 268194 241204 268200 241216
rect 268252 241204 268258 241256
rect 267734 241176 267740 241188
rect 260806 241148 264974 241176
rect 267706 241136 267740 241176
rect 267792 241136 267798 241188
rect 267706 241120 267734 241136
rect 267550 241108 267556 241120
rect 250778 240536 259454 240564
rect 260024 241080 267556 241108
rect 249288 239912 249294 239964
rect 249346 239912 249352 239964
rect 249380 239912 249386 239964
rect 249438 239912 249444 239964
rect 250116 239912 250122 239964
rect 250174 239912 250180 239964
rect 250300 239912 250306 239964
rect 250358 239912 250364 239964
rect 250392 239912 250398 239964
rect 250450 239952 250456 239964
rect 250450 239912 250484 239952
rect 250576 239912 250582 239964
rect 250634 239912 250640 239964
rect 250668 239912 250674 239964
rect 250726 239912 250732 239964
rect 249656 239844 249662 239896
rect 249714 239844 249720 239896
rect 249242 239544 249248 239556
rect 248800 239516 248920 239544
rect 249168 239516 249248 239544
rect 248892 239488 248920 239516
rect 249242 239504 249248 239516
rect 249300 239504 249306 239556
rect 249674 239544 249702 239844
rect 249794 239572 249800 239624
rect 249852 239612 249858 239624
rect 250134 239612 250162 239912
rect 250318 239884 250346 239912
rect 250318 239856 250392 239884
rect 250364 239692 250392 239856
rect 250346 239640 250352 239692
rect 250404 239640 250410 239692
rect 249852 239584 250162 239612
rect 249852 239572 249858 239584
rect 250254 239572 250260 239624
rect 250312 239612 250318 239624
rect 250456 239612 250484 239912
rect 250594 239884 250622 239912
rect 250548 239856 250622 239884
rect 250548 239624 250576 239856
rect 250686 239828 250714 239912
rect 250622 239776 250628 239828
rect 250680 239788 250714 239828
rect 250680 239776 250686 239788
rect 250778 239624 250806 240536
rect 260024 240496 260052 241080
rect 267550 241068 267556 241080
rect 267608 241068 267614 241120
rect 267642 241068 267648 241120
rect 267700 241080 267734 241120
rect 267700 241068 267706 241080
rect 313918 241040 313924 241052
rect 255286 240468 260052 240496
rect 260116 241012 313924 241040
rect 255286 240428 255314 240468
rect 252618 240400 255314 240428
rect 252250 239992 252462 240020
rect 252250 239964 252278 239992
rect 251128 239912 251134 239964
rect 251186 239912 251192 239964
rect 251220 239912 251226 239964
rect 251278 239912 251284 239964
rect 251772 239912 251778 239964
rect 251830 239912 251836 239964
rect 252232 239912 252238 239964
rect 252290 239912 252296 239964
rect 252324 239912 252330 239964
rect 252382 239912 252388 239964
rect 250944 239844 250950 239896
rect 251002 239844 251008 239896
rect 250962 239760 250990 239844
rect 251146 239816 251174 239912
rect 250898 239708 250904 239760
rect 250956 239720 250990 239760
rect 251100 239788 251174 239816
rect 250956 239708 250962 239720
rect 251100 239624 251128 239788
rect 251238 239760 251266 239912
rect 251312 239844 251318 239896
rect 251370 239844 251376 239896
rect 251588 239844 251594 239896
rect 251646 239844 251652 239896
rect 251680 239844 251686 239896
rect 251738 239844 251744 239896
rect 251174 239708 251180 239760
rect 251232 239720 251266 239760
rect 251232 239708 251238 239720
rect 251330 239624 251358 239844
rect 251606 239748 251634 239844
rect 251560 239720 251634 239748
rect 251560 239680 251588 239720
rect 251698 239692 251726 239844
rect 251790 239816 251818 239912
rect 252048 239884 252054 239896
rect 252020 239844 252054 239884
rect 252106 239844 252112 239896
rect 252140 239844 252146 239896
rect 252198 239844 252204 239896
rect 251790 239788 251956 239816
rect 251514 239652 251588 239680
rect 250312 239584 250484 239612
rect 250312 239572 250318 239584
rect 250530 239572 250536 239624
rect 250588 239572 250594 239624
rect 250714 239572 250720 239624
rect 250772 239584 250806 239624
rect 250772 239572 250778 239584
rect 251082 239572 251088 239624
rect 251140 239572 251146 239624
rect 251330 239584 251364 239624
rect 251358 239572 251364 239584
rect 251416 239572 251422 239624
rect 251514 239556 251542 239652
rect 251634 239640 251640 239692
rect 251692 239652 251726 239692
rect 251692 239640 251698 239652
rect 251928 239556 251956 239788
rect 252020 239760 252048 239844
rect 252002 239708 252008 239760
rect 252060 239708 252066 239760
rect 252158 239624 252186 239844
rect 252342 239748 252370 239912
rect 252434 239884 252462 239992
rect 252618 239964 252646 240400
rect 260116 240292 260144 241012
rect 313918 241000 313924 241012
rect 313976 241000 313982 241052
rect 267734 240932 267740 240984
rect 267792 240972 267798 240984
rect 309042 240972 309048 240984
rect 267792 240944 309048 240972
rect 267792 240932 267798 240944
rect 309042 240932 309048 240944
rect 309100 240932 309106 240984
rect 268102 240864 268108 240916
rect 268160 240904 268166 240916
rect 300394 240904 300400 240916
rect 268160 240876 300400 240904
rect 268160 240864 268166 240876
rect 300394 240864 300400 240876
rect 300452 240864 300458 240916
rect 267734 240796 267740 240848
rect 267792 240836 267798 240848
rect 316218 240836 316224 240848
rect 267792 240808 316224 240836
rect 267792 240796 267798 240808
rect 316218 240796 316224 240808
rect 316276 240796 316282 240848
rect 329098 240768 329104 240780
rect 255240 240264 260144 240292
rect 260484 240740 329104 240768
rect 255240 240020 255268 240264
rect 260484 240224 260512 240740
rect 329098 240728 329104 240740
rect 329156 240728 329162 240780
rect 267550 240660 267556 240712
rect 267608 240700 267614 240712
rect 267608 240672 273254 240700
rect 267608 240660 267614 240672
rect 267734 240632 267740 240644
rect 264394 240604 267740 240632
rect 264394 240360 264422 240604
rect 267734 240592 267740 240604
rect 267792 240592 267798 240644
rect 268286 240564 268292 240576
rect 256850 240196 260512 240224
rect 261082 240332 264422 240360
rect 264532 240536 268292 240564
rect 253400 239992 253658 240020
rect 252600 239912 252606 239964
rect 252658 239912 252664 239964
rect 252692 239912 252698 239964
rect 252750 239912 252756 239964
rect 253244 239912 253250 239964
rect 253302 239912 253308 239964
rect 252434 239856 252600 239884
rect 252416 239776 252422 239828
rect 252474 239776 252480 239828
rect 252296 239720 252370 239748
rect 252296 239692 252324 239720
rect 252434 239692 252462 239776
rect 252278 239640 252284 239692
rect 252336 239640 252342 239692
rect 252370 239640 252376 239692
rect 252428 239652 252462 239692
rect 252572 239680 252600 239856
rect 252710 239760 252738 239912
rect 252784 239844 252790 239896
rect 252842 239884 252848 239896
rect 253060 239884 253066 239896
rect 252842 239856 252968 239884
rect 252842 239844 252848 239856
rect 252710 239720 252744 239760
rect 252738 239708 252744 239720
rect 252796 239708 252802 239760
rect 252646 239680 252652 239692
rect 252572 239652 252652 239680
rect 252428 239640 252434 239652
rect 252646 239640 252652 239652
rect 252704 239640 252710 239692
rect 252158 239584 252192 239624
rect 252186 239572 252192 239584
rect 252244 239572 252250 239624
rect 252940 239612 252968 239856
rect 253032 239844 253066 239884
rect 253118 239844 253124 239896
rect 253032 239680 253060 239844
rect 253106 239708 253112 239760
rect 253164 239748 253170 239760
rect 253262 239748 253290 239912
rect 253164 239720 253290 239748
rect 253164 239708 253170 239720
rect 253400 239692 253428 239992
rect 253630 239964 253658 239992
rect 253814 239992 254256 240020
rect 253814 239964 253842 239992
rect 253520 239912 253526 239964
rect 253578 239912 253584 239964
rect 253612 239912 253618 239964
rect 253670 239912 253676 239964
rect 253796 239912 253802 239964
rect 253854 239912 253860 239964
rect 253888 239912 253894 239964
rect 253946 239912 253952 239964
rect 253032 239652 253244 239680
rect 253106 239612 253112 239624
rect 252940 239584 253112 239612
rect 253106 239572 253112 239584
rect 253164 239572 253170 239624
rect 253216 239612 253244 239652
rect 253382 239640 253388 239692
rect 253440 239640 253446 239692
rect 253538 239680 253566 239912
rect 253658 239680 253664 239692
rect 253538 239652 253664 239680
rect 253658 239640 253664 239652
rect 253716 239640 253722 239692
rect 253750 239640 253756 239692
rect 253808 239680 253814 239692
rect 253906 239680 253934 239912
rect 254072 239844 254078 239896
rect 254130 239844 254136 239896
rect 253808 239652 253934 239680
rect 254090 239692 254118 239844
rect 254228 239692 254256 239992
rect 254918 239992 255268 240020
rect 255470 240128 256786 240156
rect 254918 239964 254946 239992
rect 255470 239964 255498 240128
rect 256022 239992 256510 240020
rect 256022 239964 256050 239992
rect 254348 239912 254354 239964
rect 254406 239912 254412 239964
rect 254808 239912 254814 239964
rect 254866 239912 254872 239964
rect 254900 239912 254906 239964
rect 254958 239912 254964 239964
rect 255268 239912 255274 239964
rect 255326 239912 255332 239964
rect 255452 239912 255458 239964
rect 255510 239912 255516 239964
rect 255820 239952 255826 239964
rect 255654 239924 255826 239952
rect 254090 239652 254124 239692
rect 253808 239640 253814 239652
rect 254118 239640 254124 239652
rect 254176 239640 254182 239692
rect 254210 239640 254216 239692
rect 254268 239640 254274 239692
rect 253474 239612 253480 239624
rect 253216 239584 253480 239612
rect 253474 239572 253480 239584
rect 253532 239572 253538 239624
rect 254366 239612 254394 239912
rect 254440 239844 254446 239896
rect 254498 239844 254504 239896
rect 254624 239844 254630 239896
rect 254682 239844 254688 239896
rect 254458 239692 254486 239844
rect 254642 239748 254670 239844
rect 254826 239828 254854 239912
rect 254826 239788 254860 239828
rect 254854 239776 254860 239788
rect 254912 239776 254918 239828
rect 254642 239720 254992 239748
rect 254458 239652 254492 239692
rect 254486 239640 254492 239652
rect 254544 239640 254550 239692
rect 254762 239612 254768 239624
rect 254366 239584 254768 239612
rect 254762 239572 254768 239584
rect 254820 239572 254826 239624
rect 251266 239544 251272 239556
rect 249674 239516 251272 239544
rect 251266 239504 251272 239516
rect 251324 239504 251330 239556
rect 251514 239516 251548 239556
rect 251542 239504 251548 239516
rect 251600 239504 251606 239556
rect 251910 239504 251916 239556
rect 251968 239504 251974 239556
rect 254964 239544 254992 239720
rect 255038 239572 255044 239624
rect 255096 239612 255102 239624
rect 255286 239612 255314 239912
rect 255360 239844 255366 239896
rect 255418 239884 255424 239896
rect 255418 239844 255452 239884
rect 255544 239844 255550 239896
rect 255602 239844 255608 239896
rect 255096 239584 255314 239612
rect 255096 239572 255102 239584
rect 255314 239544 255320 239556
rect 254964 239516 255320 239544
rect 255314 239504 255320 239516
rect 255372 239504 255378 239556
rect 248380 239448 248506 239476
rect 248380 239436 248386 239448
rect 248874 239436 248880 239488
rect 248932 239436 248938 239488
rect 249058 239436 249064 239488
rect 249116 239476 249122 239488
rect 253198 239476 253204 239488
rect 249116 239448 253204 239476
rect 249116 239436 249122 239448
rect 253198 239436 253204 239448
rect 253256 239436 253262 239488
rect 255424 239476 255452 239844
rect 255562 239816 255590 239844
rect 255516 239788 255590 239816
rect 255516 239624 255544 239788
rect 255654 239624 255682 239924
rect 255820 239912 255826 239924
rect 255878 239912 255884 239964
rect 255912 239912 255918 239964
rect 255970 239912 255976 239964
rect 256004 239912 256010 239964
rect 256062 239912 256068 239964
rect 256096 239912 256102 239964
rect 256154 239952 256160 239964
rect 256372 239952 256378 239964
rect 256154 239912 256188 239952
rect 255728 239844 255734 239896
rect 255786 239844 255792 239896
rect 255498 239572 255504 239624
rect 255556 239572 255562 239624
rect 255590 239572 255596 239624
rect 255648 239584 255682 239624
rect 255746 239612 255774 239844
rect 255930 239692 255958 239912
rect 255930 239652 255964 239692
rect 255958 239640 255964 239652
rect 256016 239640 256022 239692
rect 256050 239612 256056 239624
rect 255746 239584 256056 239612
rect 255648 239572 255654 239584
rect 256050 239572 256056 239584
rect 256108 239572 256114 239624
rect 256160 239544 256188 239912
rect 256344 239912 256378 239952
rect 256430 239912 256436 239964
rect 256344 239624 256372 239912
rect 256326 239572 256332 239624
rect 256384 239572 256390 239624
rect 256482 239612 256510 239992
rect 256556 239844 256562 239896
rect 256614 239884 256620 239896
rect 256614 239844 256648 239884
rect 256620 239748 256648 239844
rect 256758 239816 256786 240128
rect 256850 239884 256878 240196
rect 261082 240156 261110 240332
rect 264532 240224 264560 240536
rect 268286 240524 268292 240536
rect 268344 240524 268350 240576
rect 273226 240496 273254 240672
rect 273226 240468 274634 240496
rect 268746 240428 268752 240440
rect 267476 240400 268752 240428
rect 267476 240360 267504 240400
rect 268746 240388 268752 240400
rect 268804 240388 268810 240440
rect 263152 240196 264560 240224
rect 265314 240332 267504 240360
rect 263152 240156 263180 240196
rect 265314 240156 265342 240332
rect 267734 240320 267740 240372
rect 267792 240360 267798 240372
rect 269298 240360 269304 240372
rect 267792 240332 269304 240360
rect 267792 240320 267798 240332
rect 269298 240320 269304 240332
rect 269356 240320 269362 240372
rect 269206 240292 269212 240304
rect 256942 240128 261110 240156
rect 261174 240128 263180 240156
rect 263244 240128 265342 240156
rect 265406 240264 269212 240292
rect 256942 239964 256970 240128
rect 257034 239992 257338 240020
rect 257034 239964 257062 239992
rect 256924 239912 256930 239964
rect 256982 239912 256988 239964
rect 257016 239912 257022 239964
rect 257074 239912 257080 239964
rect 257108 239884 257114 239896
rect 256850 239856 257114 239884
rect 257108 239844 257114 239856
rect 257166 239844 257172 239896
rect 256970 239816 256976 239828
rect 256758 239788 256976 239816
rect 256970 239776 256976 239788
rect 257028 239776 257034 239828
rect 257062 239748 257068 239760
rect 256620 239720 257068 239748
rect 257062 239708 257068 239720
rect 257120 239708 257126 239760
rect 256482 239584 256924 239612
rect 256510 239544 256516 239556
rect 256160 239516 256516 239544
rect 256510 239504 256516 239516
rect 256568 239504 256574 239556
rect 256694 239476 256700 239488
rect 255424 239448 256700 239476
rect 256694 239436 256700 239448
rect 256752 239436 256758 239488
rect 256896 239476 256924 239584
rect 256970 239572 256976 239624
rect 257028 239612 257034 239624
rect 257310 239612 257338 239992
rect 259702 239992 260190 240020
rect 259702 239964 259730 239992
rect 257752 239952 257758 239964
rect 257724 239912 257758 239952
rect 257810 239912 257816 239964
rect 257844 239912 257850 239964
rect 257902 239912 257908 239964
rect 258672 239952 258678 239964
rect 258230 239924 258678 239952
rect 257384 239844 257390 239896
rect 257442 239844 257448 239896
rect 257028 239584 257338 239612
rect 257402 239624 257430 239844
rect 257724 239680 257752 239912
rect 257862 239760 257890 239912
rect 258028 239844 258034 239896
rect 258086 239844 258092 239896
rect 258120 239844 258126 239896
rect 258178 239844 258184 239896
rect 257798 239708 257804 239760
rect 257856 239720 257890 239760
rect 257856 239708 257862 239720
rect 258046 239692 258074 239844
rect 257890 239680 257896 239692
rect 257724 239652 257896 239680
rect 257890 239640 257896 239652
rect 257948 239640 257954 239692
rect 257982 239640 257988 239692
rect 258040 239652 258074 239692
rect 258040 239640 258046 239652
rect 257402 239584 257436 239624
rect 257028 239572 257034 239584
rect 257430 239572 257436 239584
rect 257488 239572 257494 239624
rect 258138 239612 258166 239844
rect 258230 239680 258258 239924
rect 258672 239912 258678 239924
rect 258730 239912 258736 239964
rect 258856 239912 258862 239964
rect 258914 239952 258920 239964
rect 259408 239952 259414 239964
rect 258914 239924 259132 239952
rect 258914 239912 258920 239924
rect 258304 239844 258310 239896
rect 258362 239844 258368 239896
rect 258396 239844 258402 239896
rect 258454 239884 258460 239896
rect 258454 239856 258856 239884
rect 258454 239844 258460 239856
rect 258322 239760 258350 239844
rect 258322 239720 258356 239760
rect 258350 239708 258356 239720
rect 258408 239708 258414 239760
rect 258626 239680 258632 239692
rect 258230 239652 258632 239680
rect 258626 239640 258632 239652
rect 258684 239640 258690 239692
rect 258534 239612 258540 239624
rect 258138 239584 258540 239612
rect 258534 239572 258540 239584
rect 258592 239572 258598 239624
rect 258442 239504 258448 239556
rect 258500 239544 258506 239556
rect 258828 239544 258856 239856
rect 259104 239624 259132 239924
rect 259196 239924 259414 239952
rect 259196 239624 259224 239924
rect 259408 239912 259414 239924
rect 259466 239912 259472 239964
rect 259684 239912 259690 239964
rect 259742 239912 259748 239964
rect 259868 239912 259874 239964
rect 259926 239912 259932 239964
rect 259776 239844 259782 239896
rect 259834 239844 259840 239896
rect 259794 239692 259822 239844
rect 259362 239640 259368 239692
rect 259420 239640 259426 239692
rect 259730 239640 259736 239692
rect 259788 239652 259822 239692
rect 259788 239640 259794 239652
rect 259086 239572 259092 239624
rect 259144 239572 259150 239624
rect 259178 239572 259184 239624
rect 259236 239572 259242 239624
rect 259380 239612 259408 239640
rect 259886 239624 259914 239912
rect 259960 239844 259966 239896
rect 260018 239844 260024 239896
rect 259380 239584 259500 239612
rect 259472 239556 259500 239584
rect 259822 239572 259828 239624
rect 259880 239584 259914 239624
rect 259880 239572 259886 239584
rect 259978 239556 260006 239844
rect 260162 239612 260190 239992
rect 261174 239964 261202 240128
rect 263244 239964 263272 240128
rect 265406 240088 265434 240264
rect 269206 240252 269212 240264
rect 269264 240252 269270 240304
rect 268010 240224 268016 240236
rect 264302 240060 265434 240088
rect 265498 240196 268016 240224
rect 264302 239964 264330 240060
rect 265498 240020 265526 240196
rect 268010 240184 268016 240196
rect 268068 240184 268074 240236
rect 274606 240224 274634 240468
rect 309778 240224 309784 240236
rect 274606 240196 309784 240224
rect 309778 240184 309784 240196
rect 309836 240184 309842 240236
rect 265130 239992 265526 240020
rect 265774 240128 268056 240156
rect 265130 239964 265158 239992
rect 265774 239964 265802 240128
rect 267918 240088 267924 240100
rect 266004 240060 267924 240088
rect 260236 239912 260242 239964
rect 260294 239952 260300 239964
rect 260294 239924 260512 239952
rect 260294 239912 260300 239924
rect 260328 239844 260334 239896
rect 260386 239844 260392 239896
rect 260346 239692 260374 239844
rect 260282 239640 260288 239692
rect 260340 239652 260374 239692
rect 260340 239640 260346 239652
rect 260374 239612 260380 239624
rect 260162 239584 260380 239612
rect 260374 239572 260380 239584
rect 260432 239572 260438 239624
rect 258500 239516 258856 239544
rect 258500 239504 258506 239516
rect 259454 239504 259460 239556
rect 259512 239504 259518 239556
rect 259914 239504 259920 239556
rect 259972 239516 260006 239556
rect 259972 239504 259978 239516
rect 260098 239504 260104 239556
rect 260156 239544 260162 239556
rect 260484 239544 260512 239924
rect 260604 239912 260610 239964
rect 260662 239912 260668 239964
rect 260788 239952 260794 239964
rect 260760 239912 260794 239952
rect 260846 239912 260852 239964
rect 261064 239912 261070 239964
rect 261122 239912 261128 239964
rect 261156 239912 261162 239964
rect 261214 239912 261220 239964
rect 261248 239912 261254 239964
rect 261306 239912 261312 239964
rect 261340 239912 261346 239964
rect 261398 239912 261404 239964
rect 261432 239912 261438 239964
rect 261490 239912 261496 239964
rect 261616 239912 261622 239964
rect 261674 239912 261680 239964
rect 261708 239912 261714 239964
rect 261766 239912 261772 239964
rect 261984 239952 261990 239964
rect 261956 239912 261990 239952
rect 262042 239912 262048 239964
rect 262352 239912 262358 239964
rect 262410 239912 262416 239964
rect 262536 239912 262542 239964
rect 262594 239912 262600 239964
rect 262628 239912 262634 239964
rect 262686 239912 262692 239964
rect 263088 239912 263094 239964
rect 263146 239912 263152 239964
rect 263180 239912 263186 239964
rect 263238 239924 263272 239964
rect 263238 239912 263244 239924
rect 263456 239912 263462 239964
rect 263514 239952 263520 239964
rect 263514 239924 263870 239952
rect 263514 239912 263520 239924
rect 260622 239760 260650 239912
rect 260622 239720 260656 239760
rect 260650 239708 260656 239720
rect 260708 239708 260714 239760
rect 260760 239680 260788 239912
rect 260880 239884 260886 239896
rect 260852 239844 260886 239884
rect 260938 239844 260944 239896
rect 260972 239844 260978 239896
rect 261030 239844 261036 239896
rect 260852 239760 260880 239844
rect 260990 239760 261018 239844
rect 261082 239828 261110 239912
rect 261082 239788 261116 239828
rect 261110 239776 261116 239788
rect 261168 239776 261174 239828
rect 260834 239708 260840 239760
rect 260892 239708 260898 239760
rect 260990 239720 261024 239760
rect 261018 239708 261024 239720
rect 261076 239708 261082 239760
rect 260926 239680 260932 239692
rect 260760 239652 260932 239680
rect 260926 239640 260932 239652
rect 260984 239640 260990 239692
rect 260156 239516 260512 239544
rect 260156 239504 260162 239516
rect 257614 239476 257620 239488
rect 256896 239448 257620 239476
rect 257614 239436 257620 239448
rect 257672 239436 257678 239488
rect 258810 239436 258816 239488
rect 258868 239476 258874 239488
rect 260558 239476 260564 239488
rect 258868 239448 260564 239476
rect 258868 239436 258874 239448
rect 260558 239436 260564 239448
rect 260616 239436 260622 239488
rect 261266 239476 261294 239912
rect 261358 239760 261386 239912
rect 261340 239708 261346 239760
rect 261398 239708 261404 239760
rect 261450 239556 261478 239912
rect 261634 239556 261662 239912
rect 261386 239504 261392 239556
rect 261444 239516 261478 239556
rect 261444 239504 261450 239516
rect 261570 239504 261576 239556
rect 261628 239516 261662 239556
rect 261726 239544 261754 239912
rect 261800 239844 261806 239896
rect 261858 239884 261864 239896
rect 261858 239844 261892 239884
rect 261864 239692 261892 239844
rect 261956 239692 261984 239912
rect 262260 239844 262266 239896
rect 262318 239844 262324 239896
rect 262278 239692 262306 239844
rect 262370 239760 262398 239912
rect 262554 239828 262582 239912
rect 262646 239884 262674 239912
rect 262646 239856 262720 239884
rect 262554 239788 262588 239828
rect 262582 239776 262588 239788
rect 262640 239776 262646 239828
rect 262370 239720 262404 239760
rect 262398 239708 262404 239720
rect 262456 239708 262462 239760
rect 261846 239640 261852 239692
rect 261904 239640 261910 239692
rect 261938 239640 261944 239692
rect 261996 239640 262002 239692
rect 262278 239652 262312 239692
rect 262306 239640 262312 239652
rect 262364 239640 262370 239692
rect 262692 239624 262720 239856
rect 262904 239844 262910 239896
rect 262962 239844 262968 239896
rect 262996 239844 263002 239896
rect 263054 239844 263060 239896
rect 262490 239612 262496 239624
rect 262186 239584 262496 239612
rect 262186 239544 262214 239584
rect 262490 239572 262496 239584
rect 262548 239572 262554 239624
rect 262674 239572 262680 239624
rect 262732 239572 262738 239624
rect 261726 239516 262214 239544
rect 261628 239504 261634 239516
rect 262766 239504 262772 239556
rect 262824 239544 262830 239556
rect 262922 239544 262950 239844
rect 262824 239516 262950 239544
rect 263014 239544 263042 239844
rect 263106 239828 263134 239912
rect 263548 239844 263554 239896
rect 263606 239844 263612 239896
rect 263106 239788 263140 239828
rect 263134 239776 263140 239788
rect 263192 239776 263198 239828
rect 263226 239776 263232 239828
rect 263284 239776 263290 239828
rect 263244 239612 263272 239776
rect 263566 239748 263594 239844
rect 263520 239720 263594 239748
rect 263520 239692 263548 239720
rect 263502 239640 263508 239692
rect 263560 239640 263566 239692
rect 263842 239680 263870 239924
rect 263916 239912 263922 239964
rect 263974 239952 263980 239964
rect 263974 239912 264008 239952
rect 264100 239912 264106 239964
rect 264158 239912 264164 239964
rect 264192 239912 264198 239964
rect 264250 239912 264256 239964
rect 264284 239912 264290 239964
rect 264342 239912 264348 239964
rect 264652 239952 264658 239964
rect 264394 239924 264658 239952
rect 263980 239760 264008 239912
rect 264118 239816 264146 239912
rect 264072 239788 264146 239816
rect 264072 239760 264100 239788
rect 264210 239760 264238 239912
rect 263962 239708 263968 239760
rect 264020 239708 264026 239760
rect 264054 239708 264060 239760
rect 264112 239708 264118 239760
rect 264146 239708 264152 239760
rect 264204 239720 264238 239760
rect 264204 239708 264210 239720
rect 263842 239652 264330 239680
rect 263870 239612 263876 239624
rect 263244 239584 263876 239612
rect 263870 239572 263876 239584
rect 263928 239572 263934 239624
rect 263318 239544 263324 239556
rect 263014 239516 263324 239544
rect 262824 239504 262830 239516
rect 263318 239504 263324 239516
rect 263376 239504 263382 239556
rect 264302 239544 264330 239652
rect 264394 239612 264422 239924
rect 264652 239912 264658 239924
rect 264710 239912 264716 239964
rect 264744 239912 264750 239964
rect 264802 239912 264808 239964
rect 265020 239912 265026 239964
rect 265078 239912 265084 239964
rect 265112 239912 265118 239964
rect 265170 239912 265176 239964
rect 265296 239912 265302 239964
rect 265354 239912 265360 239964
rect 265388 239912 265394 239964
rect 265446 239912 265452 239964
rect 265664 239912 265670 239964
rect 265722 239912 265728 239964
rect 265756 239912 265762 239964
rect 265814 239912 265820 239964
rect 264762 239828 264790 239912
rect 265038 239884 265066 239912
rect 265038 239856 265112 239884
rect 265084 239828 265112 239856
rect 264560 239776 264566 239828
rect 264618 239776 264624 239828
rect 264698 239776 264704 239828
rect 264756 239788 264790 239828
rect 264756 239776 264762 239788
rect 265066 239776 265072 239828
rect 265124 239776 265130 239828
rect 264578 239748 264606 239776
rect 265314 239760 265342 239912
rect 264974 239748 264980 239760
rect 264578 239720 264980 239748
rect 264974 239708 264980 239720
rect 265032 239708 265038 239760
rect 265250 239708 265256 239760
rect 265308 239720 265342 239760
rect 265308 239708 265314 239720
rect 265406 239692 265434 239912
rect 265682 239828 265710 239912
rect 265682 239788 265716 239828
rect 265710 239776 265716 239788
rect 265768 239776 265774 239828
rect 265342 239640 265348 239692
rect 265400 239652 265434 239692
rect 265400 239640 265406 239652
rect 264790 239612 264796 239624
rect 264394 239584 264796 239612
rect 264790 239572 264796 239584
rect 264848 239612 264854 239624
rect 266004 239612 266032 240060
rect 267918 240048 267924 240060
rect 267976 240048 267982 240100
rect 268028 240088 268056 240128
rect 268286 240116 268292 240168
rect 268344 240156 268350 240168
rect 331582 240156 331588 240168
rect 268344 240128 331588 240156
rect 268344 240116 268350 240128
rect 331582 240116 331588 240128
rect 331640 240116 331646 240168
rect 269022 240088 269028 240100
rect 268028 240060 269028 240088
rect 269022 240048 269028 240060
rect 269080 240048 269086 240100
rect 306742 240048 306748 240100
rect 306800 240088 306806 240100
rect 314930 240088 314936 240100
rect 306800 240060 314936 240088
rect 306800 240048 306806 240060
rect 314930 240048 314936 240060
rect 314988 240048 314994 240100
rect 330386 240048 330392 240100
rect 330444 240088 330450 240100
rect 331122 240088 331128 240100
rect 330444 240060 331128 240088
rect 330444 240048 330450 240060
rect 331122 240048 331128 240060
rect 331180 240048 331186 240100
rect 267550 240020 267556 240032
rect 266326 239992 266722 240020
rect 266124 239952 266130 239964
rect 266096 239912 266130 239952
rect 266182 239912 266188 239964
rect 266216 239912 266222 239964
rect 266274 239912 266280 239964
rect 266096 239624 266124 239912
rect 266234 239748 266262 239912
rect 266326 239896 266354 239992
rect 266400 239912 266406 239964
rect 266458 239912 266464 239964
rect 266492 239912 266498 239964
rect 266550 239952 266556 239964
rect 266550 239924 266630 239952
rect 266550 239912 266556 239924
rect 266308 239844 266314 239896
rect 266366 239844 266372 239896
rect 266188 239720 266262 239748
rect 266418 239760 266446 239912
rect 266418 239720 266452 239760
rect 264848 239584 266032 239612
rect 264848 239572 264854 239584
rect 266078 239572 266084 239624
rect 266136 239572 266142 239624
rect 266188 239612 266216 239720
rect 266446 239708 266452 239720
rect 266504 239708 266510 239760
rect 266602 239624 266630 239924
rect 266694 239680 266722 239992
rect 266878 239992 267556 240020
rect 266878 239964 266906 239992
rect 267550 239980 267556 239992
rect 267608 239980 267614 240032
rect 292942 240020 292948 240032
rect 277366 239992 292948 240020
rect 266860 239912 266866 239964
rect 266918 239912 266924 239964
rect 267044 239912 267050 239964
rect 267102 239912 267108 239964
rect 267136 239912 267142 239964
rect 267194 239912 267200 239964
rect 267458 239912 267464 239964
rect 267516 239952 267522 239964
rect 267826 239952 267832 239964
rect 267516 239924 267832 239952
rect 267516 239912 267522 239924
rect 267826 239912 267832 239924
rect 267884 239912 267890 239964
rect 266768 239844 266774 239896
rect 266826 239844 266832 239896
rect 266786 239760 266814 239844
rect 267062 239760 267090 239912
rect 266786 239720 266820 239760
rect 266814 239708 266820 239720
rect 266872 239708 266878 239760
rect 266998 239708 267004 239760
rect 267056 239720 267090 239760
rect 267154 239748 267182 239912
rect 277366 239884 277394 239992
rect 292942 239980 292948 239992
rect 293000 239980 293006 240032
rect 271846 239856 277394 239884
rect 267550 239776 267556 239828
rect 267608 239816 267614 239828
rect 271846 239816 271874 239856
rect 291746 239816 291752 239828
rect 267608 239788 271874 239816
rect 274606 239788 291752 239816
rect 267608 239776 267614 239788
rect 267642 239748 267648 239760
rect 267154 239720 267648 239748
rect 267056 239708 267062 239720
rect 267642 239708 267648 239720
rect 267700 239708 267706 239760
rect 269390 239680 269396 239692
rect 266694 239652 269396 239680
rect 269390 239640 269396 239652
rect 269448 239640 269454 239692
rect 266354 239612 266360 239624
rect 266188 239584 266360 239612
rect 266354 239572 266360 239584
rect 266412 239572 266418 239624
rect 266602 239584 266636 239624
rect 266630 239572 266636 239584
rect 266688 239572 266694 239624
rect 274606 239612 274634 239788
rect 291746 239776 291752 239788
rect 291804 239776 291810 239828
rect 266832 239584 274634 239612
rect 264974 239544 264980 239556
rect 264302 239516 264980 239544
rect 264974 239504 264980 239516
rect 265032 239504 265038 239556
rect 265342 239504 265348 239556
rect 265400 239544 265406 239556
rect 266832 239544 266860 239584
rect 265400 239516 266860 239544
rect 265400 239504 265406 239516
rect 267366 239504 267372 239556
rect 267424 239544 267430 239556
rect 268194 239544 268200 239556
rect 267424 239516 268200 239544
rect 267424 239504 267430 239516
rect 268194 239504 268200 239516
rect 268252 239504 268258 239556
rect 269482 239504 269488 239556
rect 269540 239544 269546 239556
rect 286778 239544 286784 239556
rect 269540 239516 286784 239544
rect 269540 239504 269546 239516
rect 286778 239504 286784 239516
rect 286836 239504 286842 239556
rect 321094 239476 321100 239488
rect 261266 239448 321100 239476
rect 321094 239436 321100 239448
rect 321152 239436 321158 239488
rect 249610 239408 249616 239420
rect 246362 239380 249616 239408
rect 249610 239368 249616 239380
rect 249668 239368 249674 239420
rect 251634 239368 251640 239420
rect 251692 239408 251698 239420
rect 251692 239380 253704 239408
rect 251692 239368 251698 239380
rect 238110 239340 238116 239352
rect 178092 239312 238116 239340
rect 178092 239300 178098 239312
rect 238110 239300 238116 239312
rect 238168 239300 238174 239352
rect 247954 239300 247960 239352
rect 248012 239340 248018 239352
rect 249150 239340 249156 239352
rect 248012 239312 249156 239340
rect 248012 239300 248018 239312
rect 249150 239300 249156 239312
rect 249208 239300 249214 239352
rect 252554 239300 252560 239352
rect 252612 239340 252618 239352
rect 253382 239340 253388 239352
rect 252612 239312 253388 239340
rect 252612 239300 252618 239312
rect 253382 239300 253388 239312
rect 253440 239300 253446 239352
rect 253676 239340 253704 239380
rect 257338 239368 257344 239420
rect 257396 239408 257402 239420
rect 263502 239408 263508 239420
rect 257396 239380 263508 239408
rect 257396 239368 257402 239380
rect 263502 239368 263508 239380
rect 263560 239368 263566 239420
rect 266262 239368 266268 239420
rect 266320 239408 266326 239420
rect 297174 239408 297180 239420
rect 266320 239380 297180 239408
rect 266320 239368 266326 239380
rect 297174 239368 297180 239380
rect 297232 239368 297238 239420
rect 265342 239340 265348 239352
rect 253676 239312 265348 239340
rect 265342 239300 265348 239312
rect 265400 239300 265406 239352
rect 266538 239300 266544 239352
rect 266596 239340 266602 239352
rect 267366 239340 267372 239352
rect 266596 239312 267372 239340
rect 266596 239300 266602 239312
rect 267366 239300 267372 239312
rect 267424 239300 267430 239352
rect 268194 239300 268200 239352
rect 268252 239340 268258 239352
rect 274450 239340 274456 239352
rect 268252 239312 274456 239340
rect 268252 239300 268258 239312
rect 274450 239300 274456 239312
rect 274508 239300 274514 239352
rect 200114 239232 200120 239284
rect 200172 239272 200178 239284
rect 216030 239272 216036 239284
rect 200172 239244 216036 239272
rect 200172 239232 200178 239244
rect 216030 239232 216036 239244
rect 216088 239272 216094 239284
rect 216582 239272 216588 239284
rect 216088 239244 216588 239272
rect 216088 239232 216094 239244
rect 216582 239232 216588 239244
rect 216640 239232 216646 239284
rect 220262 239232 220268 239284
rect 220320 239272 220326 239284
rect 232038 239272 232044 239284
rect 220320 239244 232044 239272
rect 220320 239232 220326 239244
rect 232038 239232 232044 239244
rect 232096 239232 232102 239284
rect 232130 239232 232136 239284
rect 232188 239272 232194 239284
rect 232774 239272 232780 239284
rect 232188 239244 232780 239272
rect 232188 239232 232194 239244
rect 232774 239232 232780 239244
rect 232832 239232 232838 239284
rect 233418 239232 233424 239284
rect 233476 239272 233482 239284
rect 233476 239244 238340 239272
rect 233476 239232 233482 239244
rect 195974 239164 195980 239216
rect 196032 239204 196038 239216
rect 196032 239176 200114 239204
rect 196032 239164 196038 239176
rect 200086 239136 200114 239176
rect 219066 239164 219072 239216
rect 219124 239204 219130 239216
rect 234982 239204 234988 239216
rect 219124 239176 234988 239204
rect 219124 239164 219130 239176
rect 234982 239164 234988 239176
rect 235040 239164 235046 239216
rect 238312 239204 238340 239244
rect 247310 239232 247316 239284
rect 247368 239272 247374 239284
rect 248138 239272 248144 239284
rect 247368 239244 248144 239272
rect 247368 239232 247374 239244
rect 248138 239232 248144 239244
rect 248196 239232 248202 239284
rect 248230 239232 248236 239284
rect 248288 239272 248294 239284
rect 249334 239272 249340 239284
rect 248288 239244 249340 239272
rect 248288 239232 248294 239244
rect 249334 239232 249340 239244
rect 249392 239232 249398 239284
rect 250438 239232 250444 239284
rect 250496 239272 250502 239284
rect 252094 239272 252100 239284
rect 250496 239244 252100 239272
rect 250496 239232 250502 239244
rect 252094 239232 252100 239244
rect 252152 239232 252158 239284
rect 255038 239232 255044 239284
rect 255096 239272 255102 239284
rect 314194 239272 314200 239284
rect 255096 239244 314200 239272
rect 255096 239232 255102 239244
rect 314194 239232 314200 239244
rect 314252 239232 314258 239284
rect 252554 239204 252560 239216
rect 238312 239176 252560 239204
rect 252554 239164 252560 239176
rect 252612 239164 252618 239216
rect 256418 239164 256424 239216
rect 256476 239204 256482 239216
rect 294230 239204 294236 239216
rect 256476 239176 294236 239204
rect 256476 239164 256482 239176
rect 294230 239164 294236 239176
rect 294288 239164 294294 239216
rect 306650 239164 306656 239216
rect 306708 239204 306714 239216
rect 321554 239204 321560 239216
rect 306708 239176 321560 239204
rect 306708 239164 306714 239176
rect 321554 239164 321560 239176
rect 321612 239164 321618 239216
rect 216122 239136 216128 239148
rect 200086 239108 216128 239136
rect 216122 239096 216128 239108
rect 216180 239136 216186 239148
rect 216180 239108 229094 239136
rect 216180 239096 216186 239108
rect 215570 239028 215576 239080
rect 215628 239068 215634 239080
rect 228358 239068 228364 239080
rect 215628 239040 228364 239068
rect 215628 239028 215634 239040
rect 228358 239028 228364 239040
rect 228416 239028 228422 239080
rect 229066 239068 229094 239108
rect 229738 239096 229744 239148
rect 229796 239136 229802 239148
rect 231854 239136 231860 239148
rect 229796 239108 231860 239136
rect 229796 239096 229802 239108
rect 231854 239096 231860 239108
rect 231912 239096 231918 239148
rect 232038 239096 232044 239148
rect 232096 239136 232102 239148
rect 237742 239136 237748 239148
rect 232096 239108 237748 239136
rect 232096 239096 232102 239108
rect 237742 239096 237748 239108
rect 237800 239096 237806 239148
rect 237926 239096 237932 239148
rect 237984 239136 237990 239148
rect 238386 239136 238392 239148
rect 237984 239108 238392 239136
rect 237984 239096 237990 239108
rect 238386 239096 238392 239108
rect 238444 239136 238450 239148
rect 253934 239136 253940 239148
rect 238444 239108 253940 239136
rect 238444 239096 238450 239108
rect 253934 239096 253940 239108
rect 253992 239096 253998 239148
rect 256528 239108 260834 239136
rect 237650 239068 237656 239080
rect 229066 239040 237656 239068
rect 237650 239028 237656 239040
rect 237708 239028 237714 239080
rect 248874 239028 248880 239080
rect 248932 239068 248938 239080
rect 250714 239068 250720 239080
rect 248932 239040 250720 239068
rect 248932 239028 248938 239040
rect 250714 239028 250720 239040
rect 250772 239028 250778 239080
rect 254210 239028 254216 239080
rect 254268 239068 254274 239080
rect 254268 239040 255636 239068
rect 254268 239028 254274 239040
rect 216582 238960 216588 239012
rect 216640 239000 216646 239012
rect 238018 239000 238024 239012
rect 216640 238972 226334 239000
rect 216640 238960 216646 238972
rect 221642 238892 221648 238944
rect 221700 238932 221706 238944
rect 225598 238932 225604 238944
rect 221700 238904 225604 238932
rect 221700 238892 221706 238904
rect 225598 238892 225604 238904
rect 225656 238892 225662 238944
rect 226306 238932 226334 238972
rect 227502 238972 238024 239000
rect 227502 238932 227530 238972
rect 238018 238960 238024 238972
rect 238076 238960 238082 239012
rect 250162 238960 250168 239012
rect 250220 239000 250226 239012
rect 250438 239000 250444 239012
rect 250220 238972 250444 239000
rect 250220 238960 250226 238972
rect 250438 238960 250444 238972
rect 250496 238960 250502 239012
rect 255608 239000 255636 239040
rect 256528 239000 256556 239108
rect 257706 239028 257712 239080
rect 257764 239068 257770 239080
rect 260466 239068 260472 239080
rect 257764 239040 260472 239068
rect 257764 239028 257770 239040
rect 260466 239028 260472 239040
rect 260524 239028 260530 239080
rect 260806 239068 260834 239108
rect 261846 239096 261852 239148
rect 261904 239136 261910 239148
rect 322566 239136 322572 239148
rect 261904 239108 322572 239136
rect 261904 239096 261910 239108
rect 322566 239096 322572 239108
rect 322624 239096 322630 239148
rect 314378 239068 314384 239080
rect 260806 239040 314384 239068
rect 314378 239028 314384 239040
rect 314436 239028 314442 239080
rect 313458 239000 313464 239012
rect 255608 238972 256556 239000
rect 256666 238972 313464 239000
rect 226306 238904 227530 238932
rect 232130 238892 232136 238944
rect 232188 238932 232194 238944
rect 239582 238932 239588 238944
rect 232188 238904 239588 238932
rect 232188 238892 232194 238904
rect 239582 238892 239588 238904
rect 239640 238892 239646 238944
rect 256418 238932 256424 238944
rect 239968 238904 256424 238932
rect 217778 238824 217784 238876
rect 217836 238864 217842 238876
rect 226334 238864 226340 238876
rect 217836 238836 226340 238864
rect 217836 238824 217842 238836
rect 226334 238824 226340 238836
rect 226392 238864 226398 238876
rect 227162 238864 227168 238876
rect 226392 238836 227168 238864
rect 226392 238824 226398 238836
rect 227162 238824 227168 238836
rect 227220 238824 227226 238876
rect 233694 238824 233700 238876
rect 233752 238864 233758 238876
rect 234614 238864 234620 238876
rect 233752 238836 234620 238864
rect 233752 238824 233758 238836
rect 234614 238824 234620 238836
rect 234672 238864 234678 238876
rect 239968 238864 239996 238904
rect 256418 238892 256424 238904
rect 256476 238892 256482 238944
rect 256666 238932 256694 238972
rect 313458 238960 313464 238972
rect 313516 238960 313522 239012
rect 267550 238932 267556 238944
rect 256574 238904 256694 238932
rect 260300 238904 267556 238932
rect 234672 238836 239996 238864
rect 234672 238824 234678 238836
rect 247402 238824 247408 238876
rect 247460 238864 247466 238876
rect 248046 238864 248052 238876
rect 247460 238836 248052 238864
rect 247460 238824 247466 238836
rect 248046 238824 248052 238836
rect 248104 238824 248110 238876
rect 251634 238864 251640 238876
rect 248386 238836 251640 238864
rect 220354 238756 220360 238808
rect 220412 238796 220418 238808
rect 235166 238796 235172 238808
rect 220412 238768 235172 238796
rect 220412 238756 220418 238768
rect 235166 238756 235172 238768
rect 235224 238756 235230 238808
rect 236454 238756 236460 238808
rect 236512 238796 236518 238808
rect 236638 238796 236644 238808
rect 236512 238768 236644 238796
rect 236512 238756 236518 238768
rect 236638 238756 236644 238768
rect 236696 238756 236702 238808
rect 237926 238756 237932 238808
rect 237984 238796 237990 238808
rect 238662 238796 238668 238808
rect 237984 238768 238668 238796
rect 237984 238756 237990 238768
rect 238662 238756 238668 238768
rect 238720 238756 238726 238808
rect 239582 238756 239588 238808
rect 239640 238796 239646 238808
rect 248386 238796 248414 238836
rect 251634 238824 251640 238836
rect 251692 238824 251698 238876
rect 253382 238824 253388 238876
rect 253440 238864 253446 238876
rect 256574 238864 256602 238904
rect 253440 238836 256602 238864
rect 253440 238824 253446 238836
rect 258810 238824 258816 238876
rect 258868 238864 258874 238876
rect 260300 238864 260328 238904
rect 267550 238892 267556 238904
rect 267608 238892 267614 238944
rect 267918 238892 267924 238944
rect 267976 238932 267982 238944
rect 331122 238932 331128 238944
rect 267976 238904 331128 238932
rect 267976 238892 267982 238904
rect 331122 238892 331128 238904
rect 331180 238892 331186 238944
rect 258868 238836 260328 238864
rect 258868 238824 258874 238836
rect 260466 238824 260472 238876
rect 260524 238864 260530 238876
rect 268194 238864 268200 238876
rect 260524 238836 268200 238864
rect 260524 238824 260530 238836
rect 268194 238824 268200 238836
rect 268252 238824 268258 238876
rect 332962 238864 332968 238876
rect 273226 238836 332968 238864
rect 239640 238768 248414 238796
rect 239640 238756 239646 238768
rect 250346 238756 250352 238808
rect 250404 238796 250410 238808
rect 250898 238796 250904 238808
rect 250404 238768 250904 238796
rect 250404 238756 250410 238768
rect 250898 238756 250904 238768
rect 250956 238756 250962 238808
rect 251266 238756 251272 238808
rect 251324 238796 251330 238808
rect 254486 238796 254492 238808
rect 251324 238768 254492 238796
rect 251324 238756 251330 238768
rect 254486 238756 254492 238768
rect 254544 238756 254550 238808
rect 259178 238796 259184 238808
rect 256574 238768 259184 238796
rect 206370 238688 206376 238740
rect 206428 238728 206434 238740
rect 212074 238728 212080 238740
rect 206428 238700 212080 238728
rect 206428 238688 206434 238700
rect 212074 238688 212080 238700
rect 212132 238728 212138 238740
rect 225690 238728 225696 238740
rect 212132 238700 225696 238728
rect 212132 238688 212138 238700
rect 225690 238688 225696 238700
rect 225748 238688 225754 238740
rect 225966 238688 225972 238740
rect 226024 238728 226030 238740
rect 233142 238728 233148 238740
rect 226024 238700 233148 238728
rect 226024 238688 226030 238700
rect 233142 238688 233148 238700
rect 233200 238688 233206 238740
rect 234246 238688 234252 238740
rect 234304 238728 234310 238740
rect 239214 238728 239220 238740
rect 234304 238700 239220 238728
rect 234304 238688 234310 238700
rect 239214 238688 239220 238700
rect 239272 238688 239278 238740
rect 240870 238688 240876 238740
rect 240928 238728 240934 238740
rect 241422 238728 241428 238740
rect 240928 238700 241428 238728
rect 240928 238688 240934 238700
rect 241422 238688 241428 238700
rect 241480 238688 241486 238740
rect 241974 238688 241980 238740
rect 242032 238728 242038 238740
rect 242250 238728 242256 238740
rect 242032 238700 242256 238728
rect 242032 238688 242038 238700
rect 242250 238688 242256 238700
rect 242308 238688 242314 238740
rect 244550 238688 244556 238740
rect 244608 238728 244614 238740
rect 244734 238728 244740 238740
rect 244608 238700 244740 238728
rect 244608 238688 244614 238700
rect 244734 238688 244740 238700
rect 244792 238688 244798 238740
rect 245010 238688 245016 238740
rect 245068 238728 245074 238740
rect 245194 238728 245200 238740
rect 245068 238700 245200 238728
rect 245068 238688 245074 238700
rect 245194 238688 245200 238700
rect 245252 238688 245258 238740
rect 246022 238688 246028 238740
rect 246080 238728 246086 238740
rect 246482 238728 246488 238740
rect 246080 238700 246488 238728
rect 246080 238688 246086 238700
rect 246482 238688 246488 238700
rect 246540 238688 246546 238740
rect 246574 238688 246580 238740
rect 246632 238728 246638 238740
rect 246758 238728 246764 238740
rect 246632 238700 246764 238728
rect 246632 238688 246638 238700
rect 246758 238688 246764 238700
rect 246816 238688 246822 238740
rect 247402 238688 247408 238740
rect 247460 238728 247466 238740
rect 247586 238728 247592 238740
rect 247460 238700 247592 238728
rect 247460 238688 247466 238700
rect 247586 238688 247592 238700
rect 247644 238688 247650 238740
rect 250622 238688 250628 238740
rect 250680 238728 250686 238740
rect 250806 238728 250812 238740
rect 250680 238700 250812 238728
rect 250680 238688 250686 238700
rect 250806 238688 250812 238700
rect 250864 238688 250870 238740
rect 251726 238688 251732 238740
rect 251784 238728 251790 238740
rect 251910 238728 251916 238740
rect 251784 238700 251916 238728
rect 251784 238688 251790 238700
rect 251910 238688 251916 238700
rect 251968 238688 251974 238740
rect 256574 238728 256602 238768
rect 259178 238756 259184 238768
rect 259236 238756 259242 238808
rect 260282 238756 260288 238808
rect 260340 238796 260346 238808
rect 267918 238796 267924 238808
rect 260340 238768 267924 238796
rect 260340 238756 260346 238768
rect 267918 238756 267924 238768
rect 267976 238756 267982 238808
rect 256344 238700 256602 238728
rect 221550 238620 221556 238672
rect 221608 238660 221614 238672
rect 242986 238660 242992 238672
rect 221608 238632 242992 238660
rect 221608 238620 221614 238632
rect 242986 238620 242992 238632
rect 243044 238620 243050 238672
rect 250438 238620 250444 238672
rect 250496 238660 250502 238672
rect 250898 238660 250904 238672
rect 250496 238632 250904 238660
rect 250496 238620 250502 238632
rect 250898 238620 250904 238632
rect 250956 238620 250962 238672
rect 253198 238620 253204 238672
rect 253256 238660 253262 238672
rect 256344 238660 256372 238700
rect 263502 238688 263508 238740
rect 263560 238728 263566 238740
rect 266262 238728 266268 238740
rect 263560 238700 266268 238728
rect 263560 238688 263566 238700
rect 266262 238688 266268 238700
rect 266320 238688 266326 238740
rect 267274 238688 267280 238740
rect 267332 238728 267338 238740
rect 267734 238728 267740 238740
rect 267332 238700 267740 238728
rect 267332 238688 267338 238700
rect 267734 238688 267740 238700
rect 267792 238688 267798 238740
rect 253256 238632 256372 238660
rect 253256 238620 253262 238632
rect 260834 238620 260840 238672
rect 260892 238660 260898 238672
rect 273226 238660 273254 238836
rect 332962 238824 332968 238836
rect 333020 238824 333026 238876
rect 296622 238796 296628 238808
rect 260892 238632 273254 238660
rect 295352 238768 296628 238796
rect 260892 238620 260898 238632
rect 221366 238552 221372 238604
rect 221424 238592 221430 238604
rect 226610 238592 226616 238604
rect 221424 238564 226616 238592
rect 221424 238552 221430 238564
rect 226610 238552 226616 238564
rect 226668 238552 226674 238604
rect 229002 238552 229008 238604
rect 229060 238592 229066 238604
rect 239490 238592 239496 238604
rect 229060 238564 239496 238592
rect 229060 238552 229066 238564
rect 239490 238552 239496 238564
rect 239548 238552 239554 238604
rect 245746 238552 245752 238604
rect 245804 238592 245810 238604
rect 249058 238592 249064 238604
rect 245804 238564 249064 238592
rect 245804 238552 245810 238564
rect 249058 238552 249064 238564
rect 249116 238552 249122 238604
rect 249610 238552 249616 238604
rect 249668 238592 249674 238604
rect 253382 238592 253388 238604
rect 249668 238564 253388 238592
rect 249668 238552 249674 238564
rect 253382 238552 253388 238564
rect 253440 238552 253446 238604
rect 264238 238552 264244 238604
rect 264296 238592 264302 238604
rect 264514 238592 264520 238604
rect 264296 238564 264520 238592
rect 264296 238552 264302 238564
rect 264514 238552 264520 238564
rect 264572 238552 264578 238604
rect 212258 238484 212264 238536
rect 212316 238524 212322 238536
rect 225230 238524 225236 238536
rect 212316 238496 225236 238524
rect 212316 238484 212322 238496
rect 225230 238484 225236 238496
rect 225288 238524 225294 238536
rect 226242 238524 226248 238536
rect 225288 238496 226248 238524
rect 225288 238484 225294 238496
rect 226242 238484 226248 238496
rect 226300 238484 226306 238536
rect 227070 238484 227076 238536
rect 227128 238524 227134 238536
rect 231854 238524 231860 238536
rect 227128 238496 231860 238524
rect 227128 238484 227134 238496
rect 231854 238484 231860 238496
rect 231912 238484 231918 238536
rect 232038 238484 232044 238536
rect 232096 238524 232102 238536
rect 232866 238524 232872 238536
rect 232096 238496 232872 238524
rect 232096 238484 232102 238496
rect 232866 238484 232872 238496
rect 232924 238484 232930 238536
rect 233142 238484 233148 238536
rect 233200 238524 233206 238536
rect 238478 238524 238484 238536
rect 233200 238496 238484 238524
rect 233200 238484 233206 238496
rect 238478 238484 238484 238496
rect 238536 238484 238542 238536
rect 241514 238484 241520 238536
rect 241572 238524 241578 238536
rect 246390 238524 246396 238536
rect 241572 238496 246396 238524
rect 241572 238484 241578 238496
rect 246390 238484 246396 238496
rect 246448 238484 246454 238536
rect 248506 238484 248512 238536
rect 248564 238524 248570 238536
rect 250438 238524 250444 238536
rect 248564 238496 250444 238524
rect 248564 238484 248570 238496
rect 250438 238484 250444 238496
rect 250496 238484 250502 238536
rect 256234 238484 256240 238536
rect 256292 238524 256298 238536
rect 258994 238524 259000 238536
rect 256292 238496 259000 238524
rect 256292 238484 256298 238496
rect 258994 238484 259000 238496
rect 259052 238484 259058 238536
rect 261662 238484 261668 238536
rect 261720 238524 261726 238536
rect 295352 238524 295380 238768
rect 296622 238756 296628 238768
rect 296680 238796 296686 238808
rect 489914 238796 489920 238808
rect 296680 238768 489920 238796
rect 296680 238756 296686 238768
rect 489914 238756 489920 238768
rect 489972 238756 489978 238808
rect 261720 238496 295380 238524
rect 261720 238484 261726 238496
rect 221182 238416 221188 238468
rect 221240 238456 221246 238468
rect 224310 238456 224316 238468
rect 221240 238428 224316 238456
rect 221240 238416 221246 238428
rect 224310 238416 224316 238428
rect 224368 238416 224374 238468
rect 224586 238416 224592 238468
rect 224644 238456 224650 238468
rect 229462 238456 229468 238468
rect 224644 238428 229468 238456
rect 224644 238416 224650 238428
rect 229462 238416 229468 238428
rect 229520 238416 229526 238468
rect 229922 238416 229928 238468
rect 229980 238456 229986 238468
rect 270310 238456 270316 238468
rect 229980 238428 270316 238456
rect 229980 238416 229986 238428
rect 270310 238416 270316 238428
rect 270368 238416 270374 238468
rect 221734 238348 221740 238400
rect 221792 238388 221798 238400
rect 230382 238388 230388 238400
rect 221792 238360 230388 238388
rect 221792 238348 221798 238360
rect 230382 238348 230388 238360
rect 230440 238348 230446 238400
rect 230474 238348 230480 238400
rect 230532 238388 230538 238400
rect 270218 238388 270224 238400
rect 230532 238360 270224 238388
rect 230532 238348 230538 238360
rect 270218 238348 270224 238360
rect 270276 238348 270282 238400
rect 220262 238280 220268 238332
rect 220320 238320 220326 238332
rect 228910 238320 228916 238332
rect 220320 238292 228916 238320
rect 220320 238280 220326 238292
rect 228910 238280 228916 238292
rect 228968 238280 228974 238332
rect 231762 238280 231768 238332
rect 231820 238320 231826 238332
rect 270402 238320 270408 238332
rect 231820 238292 270408 238320
rect 231820 238280 231826 238292
rect 270402 238280 270408 238292
rect 270460 238280 270466 238332
rect 214558 238212 214564 238264
rect 214616 238252 214622 238264
rect 221182 238252 221188 238264
rect 214616 238224 221188 238252
rect 214616 238212 214622 238224
rect 221182 238212 221188 238224
rect 221240 238212 221246 238264
rect 221274 238212 221280 238264
rect 221332 238252 221338 238264
rect 225966 238252 225972 238264
rect 221332 238224 225972 238252
rect 221332 238212 221338 238224
rect 225966 238212 225972 238224
rect 226024 238212 226030 238264
rect 226610 238212 226616 238264
rect 226668 238252 226674 238264
rect 227530 238252 227536 238264
rect 226668 238224 227536 238252
rect 226668 238212 226674 238224
rect 227530 238212 227536 238224
rect 227588 238212 227594 238264
rect 230934 238212 230940 238264
rect 230992 238252 230998 238264
rect 269666 238252 269672 238264
rect 230992 238224 269672 238252
rect 230992 238212 230998 238224
rect 269666 238212 269672 238224
rect 269724 238212 269730 238264
rect 213362 238144 213368 238196
rect 213420 238184 213426 238196
rect 223942 238184 223948 238196
rect 213420 238156 223948 238184
rect 213420 238144 213426 238156
rect 223942 238144 223948 238156
rect 224000 238144 224006 238196
rect 227254 238144 227260 238196
rect 227312 238184 227318 238196
rect 232590 238184 232596 238196
rect 227312 238156 232596 238184
rect 227312 238144 227318 238156
rect 232590 238144 232596 238156
rect 232648 238144 232654 238196
rect 232774 238144 232780 238196
rect 232832 238184 232838 238196
rect 269574 238184 269580 238196
rect 232832 238156 269580 238184
rect 232832 238144 232838 238156
rect 269574 238144 269580 238156
rect 269632 238144 269638 238196
rect 194594 238076 194600 238128
rect 194652 238116 194658 238128
rect 194652 238088 215294 238116
rect 194652 238076 194658 238088
rect 85574 238008 85580 238060
rect 85632 238048 85638 238060
rect 214650 238048 214656 238060
rect 85632 238020 214656 238048
rect 85632 238008 85638 238020
rect 214650 238008 214656 238020
rect 214708 238008 214714 238060
rect 215266 237980 215294 238088
rect 221642 238076 221648 238128
rect 221700 238116 221706 238128
rect 227622 238116 227628 238128
rect 221700 238088 227628 238116
rect 221700 238076 221706 238088
rect 227622 238076 227628 238088
rect 227680 238076 227686 238128
rect 231854 238076 231860 238128
rect 231912 238116 231918 238128
rect 235810 238116 235816 238128
rect 231912 238088 235816 238116
rect 231912 238076 231918 238088
rect 235810 238076 235816 238088
rect 235868 238076 235874 238128
rect 238110 238076 238116 238128
rect 238168 238116 238174 238128
rect 239214 238116 239220 238128
rect 238168 238088 239220 238116
rect 238168 238076 238174 238088
rect 239214 238076 239220 238088
rect 239272 238076 239278 238128
rect 243814 238076 243820 238128
rect 243872 238116 243878 238128
rect 244826 238116 244832 238128
rect 243872 238088 244832 238116
rect 243872 238076 243878 238088
rect 244826 238076 244832 238088
rect 244884 238076 244890 238128
rect 245746 238076 245752 238128
rect 245804 238116 245810 238128
rect 246298 238116 246304 238128
rect 245804 238088 246304 238116
rect 245804 238076 245810 238088
rect 246298 238076 246304 238088
rect 246356 238076 246362 238128
rect 255222 238076 255228 238128
rect 255280 238116 255286 238128
rect 260466 238116 260472 238128
rect 255280 238088 260472 238116
rect 255280 238076 255286 238088
rect 260466 238076 260472 238088
rect 260524 238076 260530 238128
rect 262950 238076 262956 238128
rect 263008 238116 263014 238128
rect 264882 238116 264888 238128
rect 263008 238088 264888 238116
rect 263008 238076 263014 238088
rect 264882 238076 264888 238088
rect 264940 238076 264946 238128
rect 302694 238116 302700 238128
rect 268304 238088 302700 238116
rect 217410 238008 217416 238060
rect 217468 238048 217474 238060
rect 230198 238048 230204 238060
rect 217468 238020 230204 238048
rect 217468 238008 217474 238020
rect 230198 238008 230204 238020
rect 230256 238008 230262 238060
rect 230474 238008 230480 238060
rect 230532 238048 230538 238060
rect 231026 238048 231032 238060
rect 230532 238020 231032 238048
rect 230532 238008 230538 238020
rect 231026 238008 231032 238020
rect 231084 238008 231090 238060
rect 236178 238008 236184 238060
rect 236236 238048 236242 238060
rect 237190 238048 237196 238060
rect 236236 238020 237196 238048
rect 236236 238008 236242 238020
rect 237190 238008 237196 238020
rect 237248 238008 237254 238060
rect 240226 238008 240232 238060
rect 240284 238048 240290 238060
rect 240410 238048 240416 238060
rect 240284 238020 240416 238048
rect 240284 238008 240290 238020
rect 240410 238008 240416 238020
rect 240468 238008 240474 238060
rect 242802 238008 242808 238060
rect 242860 238048 242866 238060
rect 246942 238048 246948 238060
rect 242860 238020 246948 238048
rect 242860 238008 242866 238020
rect 246942 238008 246948 238020
rect 247000 238008 247006 238060
rect 249702 238008 249708 238060
rect 249760 238048 249766 238060
rect 250162 238048 250168 238060
rect 249760 238020 250168 238048
rect 249760 238008 249766 238020
rect 250162 238008 250168 238020
rect 250220 238008 250226 238060
rect 255958 238008 255964 238060
rect 256016 238048 256022 238060
rect 256418 238048 256424 238060
rect 256016 238020 256424 238048
rect 256016 238008 256022 238020
rect 256418 238008 256424 238020
rect 256476 238008 256482 238060
rect 256510 238008 256516 238060
rect 256568 238048 256574 238060
rect 257062 238048 257068 238060
rect 256568 238020 257068 238048
rect 256568 238008 256574 238020
rect 257062 238008 257068 238020
rect 257120 238008 257126 238060
rect 267826 238008 267832 238060
rect 267884 238048 267890 238060
rect 268304 238048 268332 238088
rect 302694 238076 302700 238088
rect 302752 238076 302758 238128
rect 267884 238020 268332 238048
rect 267884 238008 267890 238020
rect 268654 238008 268660 238060
rect 268712 238048 268718 238060
rect 308398 238048 308404 238060
rect 268712 238020 308404 238048
rect 268712 238008 268718 238020
rect 308398 238008 308404 238020
rect 308456 238008 308462 238060
rect 216398 237980 216404 237992
rect 215266 237952 216404 237980
rect 216398 237940 216404 237952
rect 216456 237980 216462 237992
rect 237558 237980 237564 237992
rect 216456 237952 237564 237980
rect 216456 237940 216462 237952
rect 237558 237940 237564 237952
rect 237616 237940 237622 237992
rect 253934 237940 253940 237992
rect 253992 237980 253998 237992
rect 257338 237980 257344 237992
rect 253992 237952 257344 237980
rect 253992 237940 253998 237952
rect 257338 237940 257344 237952
rect 257396 237940 257402 237992
rect 214650 237872 214656 237924
rect 214708 237912 214714 237924
rect 229094 237912 229100 237924
rect 214708 237884 229100 237912
rect 214708 237872 214714 237884
rect 229094 237872 229100 237884
rect 229152 237872 229158 237924
rect 231026 237872 231032 237924
rect 231084 237912 231090 237924
rect 231762 237912 231768 237924
rect 231084 237884 231768 237912
rect 231084 237872 231090 237884
rect 231762 237872 231768 237884
rect 231820 237872 231826 237924
rect 234706 237872 234712 237924
rect 234764 237912 234770 237924
rect 242158 237912 242164 237924
rect 234764 237884 242164 237912
rect 234764 237872 234770 237884
rect 242158 237872 242164 237884
rect 242216 237872 242222 237924
rect 245562 237872 245568 237924
rect 245620 237912 245626 237924
rect 257062 237912 257068 237924
rect 245620 237884 257068 237912
rect 245620 237872 245626 237884
rect 257062 237872 257068 237884
rect 257120 237872 257126 237924
rect 260558 237872 260564 237924
rect 260616 237912 260622 237924
rect 270126 237912 270132 237924
rect 260616 237884 270132 237912
rect 260616 237872 260622 237884
rect 270126 237872 270132 237884
rect 270184 237872 270190 237924
rect 221458 237804 221464 237856
rect 221516 237844 221522 237856
rect 242802 237844 242808 237856
rect 221516 237816 242808 237844
rect 221516 237804 221522 237816
rect 242802 237804 242808 237816
rect 242860 237804 242866 237856
rect 252554 237804 252560 237856
rect 252612 237844 252618 237856
rect 258718 237844 258724 237856
rect 252612 237816 258724 237844
rect 252612 237804 252618 237816
rect 258718 237804 258724 237816
rect 258776 237804 258782 237856
rect 315482 237844 315488 237856
rect 260806 237816 315488 237844
rect 221090 237736 221096 237788
rect 221148 237776 221154 237788
rect 222746 237776 222752 237788
rect 221148 237748 222752 237776
rect 221148 237736 221154 237748
rect 222746 237736 222752 237748
rect 222804 237736 222810 237788
rect 224402 237736 224408 237788
rect 224460 237776 224466 237788
rect 224862 237776 224868 237788
rect 224460 237748 224868 237776
rect 224460 237736 224466 237748
rect 224862 237736 224868 237748
rect 224920 237736 224926 237788
rect 226058 237736 226064 237788
rect 226116 237776 226122 237788
rect 226978 237776 226984 237788
rect 226116 237748 226984 237776
rect 226116 237736 226122 237748
rect 226978 237736 226984 237748
rect 227036 237736 227042 237788
rect 246114 237736 246120 237788
rect 246172 237776 246178 237788
rect 251910 237776 251916 237788
rect 246172 237748 251916 237776
rect 246172 237736 246178 237748
rect 251910 237736 251916 237748
rect 251968 237736 251974 237788
rect 256878 237736 256884 237788
rect 256936 237776 256942 237788
rect 260806 237776 260834 237816
rect 315482 237804 315488 237816
rect 315540 237804 315546 237856
rect 256936 237748 260834 237776
rect 256936 237736 256942 237748
rect 261478 237736 261484 237788
rect 261536 237776 261542 237788
rect 269114 237776 269120 237788
rect 261536 237748 269120 237776
rect 261536 237736 261542 237748
rect 269114 237736 269120 237748
rect 269172 237736 269178 237788
rect 220170 237668 220176 237720
rect 220228 237708 220234 237720
rect 228726 237708 228732 237720
rect 220228 237680 228732 237708
rect 220228 237668 220234 237680
rect 228726 237668 228732 237680
rect 228784 237668 228790 237720
rect 271046 237708 271052 237720
rect 235966 237680 271052 237708
rect 218974 237600 218980 237652
rect 219032 237640 219038 237652
rect 223298 237640 223304 237652
rect 219032 237612 223304 237640
rect 219032 237600 219038 237612
rect 223298 237600 223304 237612
rect 223356 237600 223362 237652
rect 224954 237600 224960 237652
rect 225012 237640 225018 237652
rect 225138 237640 225144 237652
rect 225012 237612 225144 237640
rect 225012 237600 225018 237612
rect 225138 237600 225144 237612
rect 225196 237600 225202 237652
rect 226150 237600 226156 237652
rect 226208 237640 226214 237652
rect 235966 237640 235994 237680
rect 271046 237668 271052 237680
rect 271104 237668 271110 237720
rect 226208 237612 235994 237640
rect 226208 237600 226214 237612
rect 243078 237600 243084 237652
rect 243136 237640 243142 237652
rect 249702 237640 249708 237652
rect 243136 237612 249708 237640
rect 243136 237600 243142 237612
rect 249702 237600 249708 237612
rect 249760 237600 249766 237652
rect 254762 237600 254768 237652
rect 254820 237640 254826 237652
rect 256878 237640 256884 237652
rect 254820 237612 256884 237640
rect 254820 237600 254826 237612
rect 256878 237600 256884 237612
rect 256936 237600 256942 237652
rect 220814 237532 220820 237584
rect 220872 237572 220878 237584
rect 224126 237572 224132 237584
rect 220872 237544 224132 237572
rect 220872 237532 220878 237544
rect 224126 237532 224132 237544
rect 224184 237532 224190 237584
rect 224862 237532 224868 237584
rect 224920 237572 224926 237584
rect 225414 237572 225420 237584
rect 224920 237544 225420 237572
rect 224920 237532 224926 237544
rect 225414 237532 225420 237544
rect 225472 237532 225478 237584
rect 231394 237532 231400 237584
rect 231452 237572 231458 237584
rect 290642 237572 290648 237584
rect 231452 237544 290648 237572
rect 231452 237532 231458 237544
rect 290642 237532 290648 237544
rect 290700 237532 290706 237584
rect 213178 237464 213184 237516
rect 213236 237504 213242 237516
rect 235718 237504 235724 237516
rect 213236 237476 235724 237504
rect 213236 237464 213242 237476
rect 235718 237464 235724 237476
rect 235776 237504 235782 237516
rect 236822 237504 236828 237516
rect 235776 237476 236828 237504
rect 235776 237464 235782 237476
rect 236822 237464 236828 237476
rect 236880 237464 236886 237516
rect 249058 237464 249064 237516
rect 249116 237504 249122 237516
rect 254762 237504 254768 237516
rect 249116 237476 254768 237504
rect 249116 237464 249122 237476
rect 254762 237464 254768 237476
rect 254820 237464 254826 237516
rect 256050 237464 256056 237516
rect 256108 237504 256114 237516
rect 315390 237504 315396 237516
rect 256108 237476 315396 237504
rect 256108 237464 256114 237476
rect 315390 237464 315396 237476
rect 315448 237464 315454 237516
rect 157334 237396 157340 237448
rect 157392 237436 157398 237448
rect 233694 237436 233700 237448
rect 157392 237408 233700 237436
rect 157392 237396 157398 237408
rect 233694 237396 233700 237408
rect 233752 237396 233758 237448
rect 267734 237396 267740 237448
rect 267792 237436 267798 237448
rect 335998 237436 336004 237448
rect 267792 237408 336004 237436
rect 267792 237396 267798 237408
rect 335998 237396 336004 237408
rect 336056 237396 336062 237448
rect 212350 237328 212356 237380
rect 212408 237368 212414 237380
rect 215294 237368 215300 237380
rect 212408 237340 215300 237368
rect 212408 237328 212414 237340
rect 215294 237328 215300 237340
rect 215352 237368 215358 237380
rect 216582 237368 216588 237380
rect 215352 237340 216588 237368
rect 215352 237328 215358 237340
rect 216582 237328 216588 237340
rect 216640 237328 216646 237380
rect 222562 237328 222568 237380
rect 222620 237368 222626 237380
rect 223114 237368 223120 237380
rect 222620 237340 223120 237368
rect 222620 237328 222626 237340
rect 223114 237328 223120 237340
rect 223172 237328 223178 237380
rect 234614 237328 234620 237380
rect 234672 237368 234678 237380
rect 239490 237368 239496 237380
rect 234672 237340 239496 237368
rect 234672 237328 234678 237340
rect 239490 237328 239496 237340
rect 239548 237328 239554 237380
rect 249978 237328 249984 237380
rect 250036 237368 250042 237380
rect 250714 237368 250720 237380
rect 250036 237340 250720 237368
rect 250036 237328 250042 237340
rect 250714 237328 250720 237340
rect 250772 237328 250778 237380
rect 265066 237328 265072 237380
rect 265124 237368 265130 237380
rect 333974 237368 333980 237380
rect 265124 237340 333980 237368
rect 265124 237328 265130 237340
rect 333974 237328 333980 237340
rect 334032 237368 334038 237380
rect 334434 237368 334440 237380
rect 334032 237340 334440 237368
rect 334032 237328 334038 237340
rect 334434 237328 334440 237340
rect 334492 237328 334498 237380
rect 220998 237260 221004 237312
rect 221056 237300 221062 237312
rect 223022 237300 223028 237312
rect 221056 237272 223028 237300
rect 221056 237260 221062 237272
rect 223022 237260 223028 237272
rect 223080 237260 223086 237312
rect 224770 237260 224776 237312
rect 224828 237300 224834 237312
rect 225138 237300 225144 237312
rect 224828 237272 225144 237300
rect 224828 237260 224834 237272
rect 225138 237260 225144 237272
rect 225196 237260 225202 237312
rect 226242 237260 226248 237312
rect 226300 237300 226306 237312
rect 232406 237300 232412 237312
rect 226300 237272 232412 237300
rect 226300 237260 226306 237272
rect 232406 237260 232412 237272
rect 232464 237260 232470 237312
rect 246942 237260 246948 237312
rect 247000 237300 247006 237312
rect 247000 237272 253934 237300
rect 247000 237260 247006 237272
rect 222654 237192 222660 237244
rect 222712 237232 222718 237244
rect 223390 237232 223396 237244
rect 222712 237204 223396 237232
rect 222712 237192 222718 237204
rect 223390 237192 223396 237204
rect 223448 237192 223454 237244
rect 253906 237232 253934 237272
rect 265618 237260 265624 237312
rect 265676 237300 265682 237312
rect 330202 237300 330208 237312
rect 265676 237272 330208 237300
rect 265676 237260 265682 237272
rect 330202 237260 330208 237272
rect 330260 237260 330266 237312
rect 260374 237232 260380 237244
rect 253906 237204 260380 237232
rect 260374 237192 260380 237204
rect 260432 237192 260438 237244
rect 260742 237192 260748 237244
rect 260800 237232 260806 237244
rect 321278 237232 321284 237244
rect 260800 237204 321284 237232
rect 260800 237192 260806 237204
rect 321278 237192 321284 237204
rect 321336 237192 321342 237244
rect 215110 237124 215116 237176
rect 215168 237164 215174 237176
rect 230014 237164 230020 237176
rect 215168 237136 230020 237164
rect 215168 237124 215174 237136
rect 230014 237124 230020 237136
rect 230072 237124 230078 237176
rect 237558 237124 237564 237176
rect 237616 237164 237622 237176
rect 240134 237164 240140 237176
rect 237616 237136 240140 237164
rect 237616 237124 237622 237136
rect 240134 237124 240140 237136
rect 240192 237164 240198 237176
rect 298094 237164 298100 237176
rect 240192 237136 298100 237164
rect 240192 237124 240198 237136
rect 298094 237124 298100 237136
rect 298152 237124 298158 237176
rect 214926 237056 214932 237108
rect 214984 237096 214990 237108
rect 225414 237096 225420 237108
rect 214984 237068 225420 237096
rect 214984 237056 214990 237068
rect 225414 237056 225420 237068
rect 225472 237056 225478 237108
rect 249334 237056 249340 237108
rect 249392 237096 249398 237108
rect 307570 237096 307576 237108
rect 249392 237068 307576 237096
rect 249392 237056 249398 237068
rect 307570 237056 307576 237068
rect 307628 237056 307634 237108
rect 215018 236988 215024 237040
rect 215076 237028 215082 237040
rect 224954 237028 224960 237040
rect 215076 237000 224960 237028
rect 215076 236988 215082 237000
rect 224954 236988 224960 237000
rect 225012 236988 225018 237040
rect 250990 236988 250996 237040
rect 251048 237028 251054 237040
rect 258994 237028 259000 237040
rect 251048 237000 259000 237028
rect 251048 236988 251054 237000
rect 258994 236988 259000 237000
rect 259052 236988 259058 237040
rect 259822 236988 259828 237040
rect 259880 237028 259886 237040
rect 319438 237028 319444 237040
rect 259880 237000 319444 237028
rect 259880 236988 259886 237000
rect 319438 236988 319444 237000
rect 319496 236988 319502 237040
rect 215846 236920 215852 236972
rect 215904 236960 215910 236972
rect 224586 236960 224592 236972
rect 215904 236932 224592 236960
rect 215904 236920 215910 236932
rect 224586 236920 224592 236932
rect 224644 236920 224650 236972
rect 232314 236920 232320 236972
rect 232372 236960 232378 236972
rect 281258 236960 281264 236972
rect 232372 236932 281264 236960
rect 232372 236920 232378 236932
rect 281258 236920 281264 236932
rect 281316 236920 281322 236972
rect 217870 236852 217876 236904
rect 217928 236892 217934 236904
rect 225966 236892 225972 236904
rect 217928 236864 225972 236892
rect 217928 236852 217934 236864
rect 225966 236852 225972 236864
rect 226024 236852 226030 236904
rect 228726 236852 228732 236904
rect 228784 236892 228790 236904
rect 231118 236892 231124 236904
rect 228784 236864 231124 236892
rect 228784 236852 228790 236864
rect 231118 236852 231124 236864
rect 231176 236852 231182 236904
rect 239214 236852 239220 236904
rect 239272 236892 239278 236904
rect 275646 236892 275652 236904
rect 239272 236864 275652 236892
rect 239272 236852 239278 236864
rect 275646 236852 275652 236864
rect 275704 236852 275710 236904
rect 331122 236852 331128 236904
rect 331180 236892 331186 236904
rect 487154 236892 487160 236904
rect 331180 236864 487160 236892
rect 331180 236852 331186 236864
rect 487154 236852 487160 236864
rect 487212 236852 487218 236904
rect 216306 236824 216312 236836
rect 215266 236796 216312 236824
rect 191834 236716 191840 236768
rect 191892 236756 191898 236768
rect 215266 236756 215294 236796
rect 216306 236784 216312 236796
rect 216364 236824 216370 236836
rect 235994 236824 236000 236836
rect 216364 236796 236000 236824
rect 216364 236784 216370 236796
rect 235994 236784 236000 236796
rect 236052 236784 236058 236836
rect 243078 236784 243084 236836
rect 243136 236824 243142 236836
rect 244182 236824 244188 236836
rect 243136 236796 244188 236824
rect 243136 236784 243142 236796
rect 244182 236784 244188 236796
rect 244240 236784 244246 236836
rect 244918 236784 244924 236836
rect 244976 236824 244982 236836
rect 279418 236824 279424 236836
rect 244976 236796 279424 236824
rect 244976 236784 244982 236796
rect 279418 236784 279424 236796
rect 279476 236784 279482 236836
rect 332962 236784 332968 236836
rect 333020 236824 333026 236836
rect 494054 236824 494060 236836
rect 333020 236796 494060 236824
rect 333020 236784 333026 236796
rect 494054 236784 494060 236796
rect 494112 236784 494118 236836
rect 191892 236728 215294 236756
rect 191892 236716 191898 236728
rect 231118 236716 231124 236768
rect 231176 236756 231182 236768
rect 231394 236756 231400 236768
rect 231176 236728 231400 236756
rect 231176 236716 231182 236728
rect 231394 236716 231400 236728
rect 231452 236716 231458 236768
rect 243446 236716 243452 236768
rect 243504 236756 243510 236768
rect 246942 236756 246948 236768
rect 243504 236728 246948 236756
rect 243504 236716 243510 236728
rect 246942 236716 246948 236728
rect 247000 236756 247006 236768
rect 278682 236756 278688 236768
rect 247000 236728 278688 236756
rect 247000 236716 247006 236728
rect 278682 236716 278688 236728
rect 278740 236716 278746 236768
rect 330202 236716 330208 236768
rect 330260 236756 330266 236768
rect 529198 236756 529204 236768
rect 330260 236728 529204 236756
rect 330260 236716 330266 236728
rect 529198 236716 529204 236728
rect 529256 236716 529262 236768
rect 126974 236648 126980 236700
rect 127032 236688 127038 236700
rect 220538 236688 220544 236700
rect 127032 236660 220544 236688
rect 127032 236648 127038 236660
rect 220538 236648 220544 236660
rect 220596 236688 220602 236700
rect 226242 236688 226248 236700
rect 220596 236660 226248 236688
rect 220596 236648 220602 236660
rect 226242 236648 226248 236660
rect 226300 236648 226306 236700
rect 231854 236648 231860 236700
rect 231912 236688 231918 236700
rect 232130 236688 232136 236700
rect 231912 236660 232136 236688
rect 231912 236648 231918 236660
rect 232130 236648 232136 236660
rect 232188 236648 232194 236700
rect 237466 236648 237472 236700
rect 237524 236688 237530 236700
rect 238110 236688 238116 236700
rect 237524 236660 238116 236688
rect 237524 236648 237530 236660
rect 238110 236648 238116 236660
rect 238168 236648 238174 236700
rect 241330 236648 241336 236700
rect 241388 236688 241394 236700
rect 244274 236688 244280 236700
rect 241388 236660 244280 236688
rect 241388 236648 241394 236660
rect 244274 236648 244280 236660
rect 244332 236648 244338 236700
rect 245930 236648 245936 236700
rect 245988 236688 245994 236700
rect 245988 236660 265756 236688
rect 245988 236648 245994 236660
rect 210970 236580 210976 236632
rect 211028 236620 211034 236632
rect 226886 236620 226892 236632
rect 211028 236592 226892 236620
rect 211028 236580 211034 236592
rect 226886 236580 226892 236592
rect 226944 236580 226950 236632
rect 256694 236580 256700 236632
rect 256752 236620 256758 236632
rect 265250 236620 265256 236632
rect 256752 236592 265256 236620
rect 256752 236580 256758 236592
rect 265250 236580 265256 236592
rect 265308 236580 265314 236632
rect 265728 236620 265756 236660
rect 266446 236648 266452 236700
rect 266504 236688 266510 236700
rect 267182 236688 267188 236700
rect 266504 236660 267188 236688
rect 266504 236648 266510 236660
rect 267182 236648 267188 236660
rect 267240 236648 267246 236700
rect 271138 236648 271144 236700
rect 271196 236688 271202 236700
rect 271690 236688 271696 236700
rect 271196 236660 271696 236688
rect 271196 236648 271202 236660
rect 271690 236648 271696 236660
rect 271748 236648 271754 236700
rect 307570 236648 307576 236700
rect 307628 236688 307634 236700
rect 332594 236688 332600 236700
rect 307628 236660 332600 236688
rect 307628 236648 307634 236660
rect 332594 236648 332600 236660
rect 332652 236648 332658 236700
rect 333974 236648 333980 236700
rect 334032 236688 334038 236700
rect 540238 236688 540244 236700
rect 334032 236660 540244 236688
rect 334032 236648 334038 236660
rect 540238 236648 540244 236660
rect 540296 236648 540302 236700
rect 271156 236620 271184 236648
rect 265728 236592 271184 236620
rect 214742 236512 214748 236564
rect 214800 236552 214806 236564
rect 220906 236552 220912 236564
rect 214800 236524 220912 236552
rect 214800 236512 214806 236524
rect 220906 236512 220912 236524
rect 220964 236552 220970 236564
rect 223666 236552 223672 236564
rect 220964 236524 223672 236552
rect 220964 236512 220970 236524
rect 223666 236512 223672 236524
rect 223724 236512 223730 236564
rect 246758 236512 246764 236564
rect 246816 236552 246822 236564
rect 255958 236552 255964 236564
rect 246816 236524 255964 236552
rect 246816 236512 246822 236524
rect 255958 236512 255964 236524
rect 256016 236512 256022 236564
rect 256786 236512 256792 236564
rect 256844 236552 256850 236564
rect 257982 236552 257988 236564
rect 256844 236524 257988 236552
rect 256844 236512 256850 236524
rect 257982 236512 257988 236524
rect 258040 236512 258046 236564
rect 213546 236444 213552 236496
rect 213604 236484 213610 236496
rect 229370 236484 229376 236496
rect 213604 236456 229376 236484
rect 213604 236444 213610 236456
rect 229370 236444 229376 236456
rect 229428 236444 229434 236496
rect 253658 236444 253664 236496
rect 253716 236484 253722 236496
rect 261662 236484 261668 236496
rect 253716 236456 261668 236484
rect 253716 236444 253722 236456
rect 261662 236444 261668 236456
rect 261720 236444 261726 236496
rect 253014 236376 253020 236428
rect 253072 236416 253078 236428
rect 256786 236416 256792 236428
rect 253072 236388 256792 236416
rect 253072 236376 253078 236388
rect 256786 236376 256792 236388
rect 256844 236376 256850 236428
rect 258718 236376 258724 236428
rect 258776 236416 258782 236428
rect 269758 236416 269764 236428
rect 258776 236388 269764 236416
rect 258776 236376 258782 236388
rect 269758 236376 269764 236388
rect 269816 236376 269822 236428
rect 213914 236308 213920 236360
rect 213972 236348 213978 236360
rect 214466 236348 214472 236360
rect 213972 236320 214472 236348
rect 213972 236308 213978 236320
rect 214466 236308 214472 236320
rect 214524 236308 214530 236360
rect 224218 236308 224224 236360
rect 224276 236348 224282 236360
rect 224494 236348 224500 236360
rect 224276 236320 224500 236348
rect 224276 236308 224282 236320
rect 224494 236308 224500 236320
rect 224552 236308 224558 236360
rect 235166 236308 235172 236360
rect 235224 236348 235230 236360
rect 282730 236348 282736 236360
rect 235224 236320 282736 236348
rect 235224 236308 235230 236320
rect 282730 236308 282736 236320
rect 282788 236308 282794 236360
rect 220722 236240 220728 236292
rect 220780 236280 220786 236292
rect 223574 236280 223580 236292
rect 220780 236252 223580 236280
rect 220780 236240 220786 236252
rect 223574 236240 223580 236252
rect 223632 236240 223638 236292
rect 228358 236240 228364 236292
rect 228416 236280 228422 236292
rect 235442 236280 235448 236292
rect 228416 236252 235448 236280
rect 228416 236240 228422 236252
rect 235442 236240 235448 236252
rect 235500 236280 235506 236292
rect 278130 236280 278136 236292
rect 235500 236252 278136 236280
rect 235500 236240 235506 236252
rect 278130 236240 278136 236252
rect 278188 236240 278194 236292
rect 244826 236172 244832 236224
rect 244884 236212 244890 236224
rect 258718 236212 258724 236224
rect 244884 236184 258724 236212
rect 244884 236172 244890 236184
rect 258718 236172 258724 236184
rect 258776 236172 258782 236224
rect 249886 236104 249892 236156
rect 249944 236144 249950 236156
rect 250346 236144 250352 236156
rect 249944 236116 250352 236144
rect 249944 236104 249950 236116
rect 250346 236104 250352 236116
rect 250404 236104 250410 236156
rect 252370 236104 252376 236156
rect 252428 236144 252434 236156
rect 260742 236144 260748 236156
rect 252428 236116 260748 236144
rect 252428 236104 252434 236116
rect 260742 236104 260748 236116
rect 260800 236104 260806 236156
rect 266170 236036 266176 236088
rect 266228 236076 266234 236088
rect 269022 236076 269028 236088
rect 266228 236048 269028 236076
rect 266228 236036 266234 236048
rect 269022 236036 269028 236048
rect 269080 236036 269086 236088
rect 214650 235968 214656 236020
rect 214708 236008 214714 236020
rect 215110 236008 215116 236020
rect 214708 235980 215116 236008
rect 214708 235968 214714 235980
rect 215110 235968 215116 235980
rect 215168 235968 215174 236020
rect 252922 235968 252928 236020
rect 252980 236008 252986 236020
rect 256142 236008 256148 236020
rect 252980 235980 256148 236008
rect 252980 235968 252986 235980
rect 256142 235968 256148 235980
rect 256200 235968 256206 236020
rect 263778 235968 263784 236020
rect 263836 236008 263842 236020
rect 264146 236008 264152 236020
rect 263836 235980 264152 236008
rect 263836 235968 263842 235980
rect 264146 235968 264152 235980
rect 264204 235968 264210 236020
rect 212442 235900 212448 235952
rect 212500 235940 212506 235952
rect 229186 235940 229192 235952
rect 212500 235912 229192 235940
rect 212500 235900 212506 235912
rect 229186 235900 229192 235912
rect 229244 235900 229250 235952
rect 251542 235900 251548 235952
rect 251600 235940 251606 235952
rect 253198 235940 253204 235952
rect 251600 235912 253204 235940
rect 251600 235900 251606 235912
rect 253198 235900 253204 235912
rect 253256 235900 253262 235952
rect 253934 235900 253940 235952
rect 253992 235940 253998 235952
rect 337010 235940 337016 235952
rect 253992 235912 337016 235940
rect 253992 235900 253998 235912
rect 337010 235900 337016 235912
rect 337068 235940 337074 235952
rect 338022 235940 338028 235952
rect 337068 235912 338028 235940
rect 337068 235900 337074 235912
rect 338022 235900 338028 235912
rect 338080 235900 338086 235952
rect 256510 235832 256516 235884
rect 256568 235872 256574 235884
rect 263134 235872 263140 235884
rect 256568 235844 263140 235872
rect 256568 235832 256574 235844
rect 263134 235832 263140 235844
rect 263192 235832 263198 235884
rect 265434 235832 265440 235884
rect 265492 235872 265498 235884
rect 331490 235872 331496 235884
rect 265492 235844 331496 235872
rect 265492 235832 265498 235844
rect 331490 235832 331496 235844
rect 331548 235832 331554 235884
rect 220814 235764 220820 235816
rect 220872 235804 220878 235816
rect 237650 235804 237656 235816
rect 220872 235776 237656 235804
rect 220872 235764 220878 235776
rect 237650 235764 237656 235776
rect 237708 235764 237714 235816
rect 250898 235764 250904 235816
rect 250956 235804 250962 235816
rect 267734 235804 267740 235816
rect 250956 235776 267740 235804
rect 250956 235764 250962 235776
rect 267734 235764 267740 235776
rect 267792 235764 267798 235816
rect 218606 235696 218612 235748
rect 218664 235736 218670 235748
rect 230474 235736 230480 235748
rect 218664 235708 230480 235736
rect 218664 235696 218670 235708
rect 230474 235696 230480 235708
rect 230532 235696 230538 235748
rect 294598 235736 294604 235748
rect 241486 235708 294604 235736
rect 209774 235628 209780 235680
rect 209832 235668 209838 235680
rect 238754 235668 238760 235680
rect 209832 235640 238760 235668
rect 209832 235628 209838 235640
rect 238754 235628 238760 235640
rect 238812 235668 238818 235680
rect 241486 235668 241514 235708
rect 294598 235696 294604 235708
rect 294656 235696 294662 235748
rect 238812 235640 241514 235668
rect 238812 235628 238818 235640
rect 246574 235628 246580 235680
rect 246632 235668 246638 235680
rect 298738 235668 298744 235680
rect 246632 235640 298744 235668
rect 246632 235628 246638 235640
rect 298738 235628 298744 235640
rect 298796 235628 298802 235680
rect 211154 235560 211160 235612
rect 211212 235600 211218 235612
rect 238938 235600 238944 235612
rect 211212 235572 238944 235600
rect 211212 235560 211218 235572
rect 238938 235560 238944 235572
rect 238996 235600 239002 235612
rect 286870 235600 286876 235612
rect 238996 235572 286876 235600
rect 238996 235560 239002 235572
rect 286870 235560 286876 235572
rect 286928 235560 286934 235612
rect 175918 235492 175924 235544
rect 175976 235532 175982 235544
rect 226150 235532 226156 235544
rect 175976 235504 226156 235532
rect 175976 235492 175982 235504
rect 226150 235492 226156 235504
rect 226208 235492 226214 235544
rect 235994 235492 236000 235544
rect 236052 235532 236058 235544
rect 236178 235532 236184 235544
rect 236052 235504 236184 235532
rect 236052 235492 236058 235504
rect 236178 235492 236184 235504
rect 236236 235532 236242 235544
rect 282638 235532 282644 235544
rect 236236 235504 282644 235532
rect 236236 235492 236242 235504
rect 282638 235492 282644 235504
rect 282696 235492 282702 235544
rect 115198 235424 115204 235476
rect 115256 235464 115262 235476
rect 230566 235464 230572 235476
rect 115256 235436 230572 235464
rect 115256 235424 115262 235436
rect 230566 235424 230572 235436
rect 230624 235424 230630 235476
rect 235718 235424 235724 235476
rect 235776 235464 235782 235476
rect 275278 235464 275284 235476
rect 235776 235436 275284 235464
rect 235776 235424 235782 235436
rect 275278 235424 275284 235436
rect 275336 235424 275342 235476
rect 95878 235356 95884 235408
rect 95936 235396 95942 235408
rect 212442 235396 212448 235408
rect 95936 235368 212448 235396
rect 95936 235356 95942 235368
rect 212442 235356 212448 235368
rect 212500 235356 212506 235408
rect 213270 235356 213276 235408
rect 213328 235396 213334 235408
rect 237374 235396 237380 235408
rect 213328 235368 237380 235396
rect 213328 235356 213334 235368
rect 237374 235356 237380 235368
rect 237432 235396 237438 235408
rect 237432 235368 238800 235396
rect 237432 235356 237438 235368
rect 106274 235288 106280 235340
rect 106332 235328 106338 235340
rect 230842 235328 230848 235340
rect 106332 235300 230848 235328
rect 106332 235288 106338 235300
rect 230842 235288 230848 235300
rect 230900 235288 230906 235340
rect 232498 235288 232504 235340
rect 232556 235328 232562 235340
rect 232866 235328 232872 235340
rect 232556 235300 232872 235328
rect 232556 235288 232562 235300
rect 232866 235288 232872 235300
rect 232924 235288 232930 235340
rect 60734 235220 60740 235272
rect 60792 235260 60798 235272
rect 226794 235260 226800 235272
rect 60792 235232 226800 235260
rect 60792 235220 60798 235232
rect 226794 235220 226800 235232
rect 226852 235220 226858 235272
rect 228726 235220 228732 235272
rect 228784 235260 228790 235272
rect 237558 235260 237564 235272
rect 228784 235232 237564 235260
rect 228784 235220 228790 235232
rect 237558 235220 237564 235232
rect 237616 235220 237622 235272
rect 224034 235152 224040 235204
rect 224092 235192 224098 235204
rect 224678 235192 224684 235204
rect 224092 235164 224684 235192
rect 224092 235152 224098 235164
rect 224678 235152 224684 235164
rect 224736 235152 224742 235204
rect 238772 235192 238800 235368
rect 244366 235356 244372 235408
rect 244424 235396 244430 235408
rect 281534 235396 281540 235408
rect 244424 235368 281540 235396
rect 244424 235356 244430 235368
rect 281534 235356 281540 235368
rect 281592 235396 281598 235408
rect 282822 235396 282828 235408
rect 281592 235368 282828 235396
rect 281592 235356 281598 235368
rect 282822 235356 282828 235368
rect 282880 235356 282886 235408
rect 338022 235356 338028 235408
rect 338080 235396 338086 235408
rect 369854 235396 369860 235408
rect 338080 235368 369860 235396
rect 338080 235356 338086 235368
rect 369854 235356 369860 235368
rect 369912 235356 369918 235408
rect 243262 235288 243268 235340
rect 243320 235328 243326 235340
rect 262950 235328 262956 235340
rect 243320 235300 262956 235328
rect 243320 235288 243326 235300
rect 262950 235288 262956 235300
rect 263008 235288 263014 235340
rect 263474 235300 270494 235328
rect 243998 235220 244004 235272
rect 244056 235260 244062 235272
rect 263474 235260 263502 235300
rect 244056 235232 263502 235260
rect 244056 235220 244062 235232
rect 266354 235220 266360 235272
rect 266412 235260 266418 235272
rect 266814 235260 266820 235272
rect 266412 235232 266820 235260
rect 266412 235220 266418 235232
rect 266814 235220 266820 235232
rect 266872 235220 266878 235272
rect 270466 235260 270494 235300
rect 331582 235288 331588 235340
rect 331640 235328 331646 235340
rect 498286 235328 498292 235340
rect 331640 235300 498292 235328
rect 331640 235288 331646 235300
rect 498286 235288 498292 235300
rect 498344 235288 498350 235340
rect 275922 235260 275928 235272
rect 270466 235232 275928 235260
rect 275922 235220 275928 235232
rect 275980 235260 275986 235272
rect 294690 235260 294696 235272
rect 275980 235232 294696 235260
rect 275980 235220 275986 235232
rect 294690 235220 294696 235232
rect 294748 235220 294754 235272
rect 331490 235220 331496 235272
rect 331548 235260 331554 235272
rect 550634 235260 550640 235272
rect 331548 235232 550640 235260
rect 331548 235220 331554 235232
rect 550634 235220 550640 235232
rect 550692 235220 550698 235272
rect 238772 235164 244274 235192
rect 244246 235124 244274 235164
rect 258166 235152 258172 235204
rect 258224 235192 258230 235204
rect 258442 235192 258448 235204
rect 258224 235164 258448 235192
rect 258224 235152 258230 235164
rect 258442 235152 258448 235164
rect 258500 235152 258506 235204
rect 262214 235152 262220 235204
rect 262272 235192 262278 235204
rect 262858 235192 262864 235204
rect 262272 235164 262864 235192
rect 262272 235152 262278 235164
rect 262858 235152 262864 235164
rect 262916 235152 262922 235204
rect 262950 235152 262956 235204
rect 263008 235192 263014 235204
rect 267826 235192 267832 235204
rect 263008 235164 267832 235192
rect 263008 235152 263014 235164
rect 267826 235152 267832 235164
rect 267884 235152 267890 235204
rect 272978 235124 272984 235136
rect 244246 235096 272984 235124
rect 272978 235084 272984 235096
rect 273036 235084 273042 235136
rect 237650 235016 237656 235068
rect 237708 235056 237714 235068
rect 239674 235056 239680 235068
rect 237708 235028 239680 235056
rect 237708 235016 237714 235028
rect 239674 235016 239680 235028
rect 239732 235056 239738 235068
rect 296254 235056 296260 235068
rect 239732 235028 296260 235056
rect 239732 235016 239738 235028
rect 296254 235016 296260 235028
rect 296312 235016 296318 235068
rect 235810 234948 235816 235000
rect 235868 234988 235874 235000
rect 279878 234988 279884 235000
rect 235868 234960 279884 234988
rect 235868 234948 235874 234960
rect 279878 234948 279884 234960
rect 279936 234948 279942 235000
rect 251174 234880 251180 234932
rect 251232 234920 251238 234932
rect 253934 234920 253940 234932
rect 251232 234892 253940 234920
rect 251232 234880 251238 234892
rect 253934 234880 253940 234892
rect 253992 234880 253998 234932
rect 257430 234880 257436 234932
rect 257488 234920 257494 234932
rect 260190 234920 260196 234932
rect 257488 234892 260196 234920
rect 257488 234880 257494 234892
rect 260190 234880 260196 234892
rect 260248 234880 260254 234932
rect 262306 234880 262312 234932
rect 262364 234920 262370 234932
rect 263410 234920 263416 234932
rect 262364 234892 263416 234920
rect 262364 234880 262370 234892
rect 263410 234880 263416 234892
rect 263468 234880 263474 234932
rect 236086 234608 236092 234660
rect 236144 234648 236150 234660
rect 236454 234648 236460 234660
rect 236144 234620 236460 234648
rect 236144 234608 236150 234620
rect 236454 234608 236460 234620
rect 236512 234608 236518 234660
rect 331490 234608 331496 234660
rect 331548 234648 331554 234660
rect 331950 234648 331956 234660
rect 331548 234620 331956 234648
rect 331548 234608 331554 234620
rect 331950 234608 331956 234620
rect 332008 234648 332014 234660
rect 512638 234648 512644 234660
rect 332008 234620 512644 234648
rect 332008 234608 332014 234620
rect 512638 234608 512644 234620
rect 512696 234608 512702 234660
rect 234246 234540 234252 234592
rect 234304 234580 234310 234592
rect 294138 234580 294144 234592
rect 234304 234552 294144 234580
rect 234304 234540 234310 234552
rect 294138 234540 294144 234552
rect 294196 234540 294202 234592
rect 234338 234472 234344 234524
rect 234396 234512 234402 234524
rect 292758 234512 292764 234524
rect 234396 234484 292764 234512
rect 234396 234472 234402 234484
rect 292758 234472 292764 234484
rect 292816 234472 292822 234524
rect 234798 234404 234804 234456
rect 234856 234444 234862 234456
rect 235350 234444 235356 234456
rect 234856 234416 235356 234444
rect 234856 234404 234862 234416
rect 235350 234404 235356 234416
rect 235408 234404 235414 234456
rect 236546 234404 236552 234456
rect 236604 234444 236610 234456
rect 239398 234444 239404 234456
rect 236604 234416 239404 234444
rect 236604 234404 236610 234416
rect 239398 234404 239404 234416
rect 239456 234444 239462 234456
rect 299198 234444 299204 234456
rect 239456 234416 299204 234444
rect 239456 234404 239462 234416
rect 299198 234404 299204 234416
rect 299256 234404 299262 234456
rect 247494 234336 247500 234388
rect 247552 234376 247558 234388
rect 306650 234376 306656 234388
rect 247552 234348 306656 234376
rect 247552 234336 247558 234348
rect 306650 234336 306656 234348
rect 306708 234336 306714 234388
rect 233970 234268 233976 234320
rect 234028 234308 234034 234320
rect 292850 234308 292856 234320
rect 234028 234280 292856 234308
rect 234028 234268 234034 234280
rect 292850 234268 292856 234280
rect 292908 234268 292914 234320
rect 231762 234200 231768 234252
rect 231820 234240 231826 234252
rect 240502 234240 240508 234252
rect 231820 234212 240508 234240
rect 231820 234200 231826 234212
rect 240502 234200 240508 234212
rect 240560 234240 240566 234252
rect 298830 234240 298836 234252
rect 240560 234212 298836 234240
rect 240560 234200 240566 234212
rect 298830 234200 298836 234212
rect 298888 234200 298894 234252
rect 254026 234132 254032 234184
rect 254084 234172 254090 234184
rect 311802 234172 311808 234184
rect 254084 234144 311808 234172
rect 254084 234132 254090 234144
rect 311802 234132 311808 234144
rect 311860 234172 311866 234184
rect 311860 234144 316034 234172
rect 311860 234132 311866 234144
rect 229554 234064 229560 234116
rect 229612 234104 229618 234116
rect 230198 234104 230204 234116
rect 229612 234076 230204 234104
rect 229612 234064 229618 234076
rect 230198 234064 230204 234076
rect 230256 234064 230262 234116
rect 235718 234064 235724 234116
rect 235776 234104 235782 234116
rect 236730 234104 236736 234116
rect 235776 234076 236736 234104
rect 235776 234064 235782 234076
rect 236730 234064 236736 234076
rect 236788 234104 236794 234116
rect 293218 234104 293224 234116
rect 236788 234076 293224 234104
rect 236788 234064 236794 234076
rect 293218 234064 293224 234076
rect 293276 234064 293282 234116
rect 218054 233996 218060 234048
rect 218112 234036 218118 234048
rect 236546 234036 236552 234048
rect 218112 234008 236552 234036
rect 218112 233996 218118 234008
rect 236546 233996 236552 234008
rect 236604 233996 236610 234048
rect 241514 233996 241520 234048
rect 241572 234036 241578 234048
rect 242250 234036 242256 234048
rect 241572 234008 242256 234036
rect 241572 233996 241578 234008
rect 242250 233996 242256 234008
rect 242308 233996 242314 234048
rect 243170 233996 243176 234048
rect 243228 234036 243234 234048
rect 244182 234036 244188 234048
rect 243228 234008 244188 234036
rect 243228 233996 243234 234008
rect 244182 233996 244188 234008
rect 244240 233996 244246 234048
rect 247126 233996 247132 234048
rect 247184 234036 247190 234048
rect 247184 234008 296714 234036
rect 247184 233996 247190 234008
rect 228266 233928 228272 233980
rect 228324 233968 228330 233980
rect 228818 233968 228824 233980
rect 228324 233940 228824 233968
rect 228324 233928 228330 233940
rect 228818 233928 228824 233940
rect 228876 233928 228882 233980
rect 232958 233928 232964 233980
rect 233016 233968 233022 233980
rect 282454 233968 282460 233980
rect 233016 233940 282460 233968
rect 233016 233928 233022 233940
rect 282454 233928 282460 233940
rect 282512 233928 282518 233980
rect 296686 233968 296714 234008
rect 300946 233968 300952 233980
rect 296686 233940 300952 233968
rect 300946 233928 300952 233940
rect 301004 233968 301010 233980
rect 313918 233968 313924 233980
rect 301004 233940 313924 233968
rect 301004 233928 301010 233940
rect 313918 233928 313924 233940
rect 313976 233928 313982 233980
rect 143534 233860 143540 233912
rect 143592 233900 143598 233912
rect 233602 233900 233608 233912
rect 143592 233872 233608 233900
rect 143592 233860 143598 233872
rect 233602 233860 233608 233872
rect 233660 233900 233666 233912
rect 234338 233900 234344 233912
rect 233660 233872 234344 233900
rect 233660 233860 233666 233872
rect 234338 233860 234344 233872
rect 234396 233860 234402 233912
rect 237558 233860 237564 233912
rect 237616 233900 237622 233912
rect 238386 233900 238392 233912
rect 237616 233872 238392 233900
rect 237616 233860 237622 233872
rect 238386 233860 238392 233872
rect 238444 233860 238450 233912
rect 241514 233860 241520 233912
rect 241572 233900 241578 233912
rect 241882 233900 241888 233912
rect 241572 233872 241888 233900
rect 241572 233860 241578 233872
rect 241882 233860 241888 233872
rect 241940 233860 241946 233912
rect 245378 233860 245384 233912
rect 245436 233900 245442 233912
rect 277210 233900 277216 233912
rect 245436 233872 277216 233900
rect 245436 233860 245442 233872
rect 277210 233860 277216 233872
rect 277268 233900 277274 233912
rect 278038 233900 278044 233912
rect 277268 233872 278044 233900
rect 277268 233860 277274 233872
rect 278038 233860 278044 233872
rect 278096 233860 278102 233912
rect 316006 233900 316034 234144
rect 405734 233900 405740 233912
rect 316006 233872 405740 233900
rect 405734 233860 405740 233872
rect 405792 233860 405798 233912
rect 227898 233792 227904 233844
rect 227956 233832 227962 233844
rect 228542 233832 228548 233844
rect 227956 233804 228548 233832
rect 227956 233792 227962 233804
rect 228542 233792 228548 233804
rect 228600 233792 228606 233844
rect 229738 233792 229744 233844
rect 229796 233832 229802 233844
rect 230382 233832 230388 233844
rect 229796 233804 230388 233832
rect 229796 233792 229802 233804
rect 230382 233792 230388 233804
rect 230440 233792 230446 233844
rect 245102 233792 245108 233844
rect 245160 233832 245166 233844
rect 274542 233832 274548 233844
rect 245160 233804 274548 233832
rect 245160 233792 245166 233804
rect 274542 233792 274548 233804
rect 274600 233832 274606 233844
rect 275278 233832 275284 233844
rect 274600 233804 275284 233832
rect 274600 233792 274606 233804
rect 275278 233792 275284 233804
rect 275336 233792 275342 233844
rect 271230 233764 271236 233776
rect 244246 233736 271236 233764
rect 243538 233656 243544 233708
rect 243596 233696 243602 233708
rect 244246 233696 244274 233736
rect 271230 233724 271236 233736
rect 271288 233724 271294 233776
rect 272610 233696 272616 233708
rect 243596 233668 244274 233696
rect 263566 233668 272616 233696
rect 243596 233656 243602 233668
rect 226610 233588 226616 233640
rect 226668 233628 226674 233640
rect 227346 233628 227352 233640
rect 226668 233600 227352 233628
rect 226668 233588 226674 233600
rect 227346 233588 227352 233600
rect 227404 233588 227410 233640
rect 227990 233588 227996 233640
rect 228048 233628 228054 233640
rect 228450 233628 228456 233640
rect 228048 233600 228456 233628
rect 228048 233588 228054 233600
rect 228450 233588 228456 233600
rect 228508 233588 228514 233640
rect 233602 233452 233608 233504
rect 233660 233492 233666 233504
rect 234154 233492 234160 233504
rect 233660 233464 234160 233492
rect 233660 233452 233666 233464
rect 234154 233452 234160 233464
rect 234212 233452 234218 233504
rect 227806 233384 227812 233436
rect 227864 233384 227870 233436
rect 249702 233384 249708 233436
rect 249760 233424 249766 233436
rect 263566 233424 263594 233668
rect 272610 233656 272616 233668
rect 272668 233656 272674 233708
rect 249760 233396 263594 233424
rect 249760 233384 249766 233396
rect 227824 233096 227852 233384
rect 256786 233316 256792 233368
rect 256844 233356 256850 233368
rect 257430 233356 257436 233368
rect 256844 233328 257436 233356
rect 256844 233316 256850 233328
rect 257430 233316 257436 233328
rect 257488 233316 257494 233368
rect 234062 233180 234068 233232
rect 234120 233220 234126 233232
rect 294506 233220 294512 233232
rect 234120 233192 294512 233220
rect 234120 233180 234126 233192
rect 294506 233180 294512 233192
rect 294564 233180 294570 233232
rect 345658 233180 345664 233232
rect 345716 233220 345722 233232
rect 579982 233220 579988 233232
rect 345716 233192 579988 233220
rect 345716 233180 345722 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 241974 233112 241980 233164
rect 242032 233152 242038 233164
rect 242710 233152 242716 233164
rect 242032 233124 242716 233152
rect 242032 233112 242038 233124
rect 242710 233112 242716 233124
rect 242768 233112 242774 233164
rect 249794 233112 249800 233164
rect 249852 233152 249858 233164
rect 310146 233152 310152 233164
rect 249852 233124 310152 233152
rect 249852 233112 249858 233124
rect 310146 233112 310152 233124
rect 310204 233152 310210 233164
rect 310422 233152 310428 233164
rect 310204 233124 310428 233152
rect 310204 233112 310210 233124
rect 310422 233112 310428 233124
rect 310480 233112 310486 233164
rect 227806 233044 227812 233096
rect 227864 233044 227870 233096
rect 247402 233044 247408 233096
rect 247460 233084 247466 233096
rect 303706 233084 303712 233096
rect 247460 233056 303712 233084
rect 247460 233044 247466 233056
rect 303706 233044 303712 233056
rect 303764 233044 303770 233096
rect 242158 232976 242164 233028
rect 242216 233016 242222 233028
rect 251174 233016 251180 233028
rect 242216 232988 251180 233016
rect 242216 232976 242222 232988
rect 251174 232976 251180 232988
rect 251232 232976 251238 233028
rect 254486 232976 254492 233028
rect 254544 233016 254550 233028
rect 309502 233016 309508 233028
rect 254544 232988 309508 233016
rect 254544 232976 254550 232988
rect 309502 232976 309508 232988
rect 309560 232976 309566 233028
rect 239582 232908 239588 232960
rect 239640 232948 239646 232960
rect 239858 232948 239864 232960
rect 239640 232920 239864 232948
rect 239640 232908 239646 232920
rect 239858 232908 239864 232920
rect 239916 232948 239922 232960
rect 292022 232948 292028 232960
rect 239916 232920 292028 232948
rect 239916 232908 239922 232920
rect 292022 232908 292028 232920
rect 292080 232908 292086 232960
rect 191098 232840 191104 232892
rect 191156 232880 191162 232892
rect 235994 232880 236000 232892
rect 191156 232852 236000 232880
rect 191156 232840 191162 232852
rect 235994 232840 236000 232852
rect 236052 232840 236058 232892
rect 245654 232840 245660 232892
rect 245712 232880 245718 232892
rect 295978 232880 295984 232892
rect 245712 232852 295984 232880
rect 245712 232840 245718 232852
rect 295978 232840 295984 232852
rect 296036 232840 296042 232892
rect 183554 232772 183560 232824
rect 183612 232812 183618 232824
rect 235718 232812 235724 232824
rect 183612 232784 235724 232812
rect 183612 232772 183618 232784
rect 235718 232772 235724 232784
rect 235776 232772 235782 232824
rect 238754 232772 238760 232824
rect 238812 232812 238818 232824
rect 240962 232812 240968 232824
rect 238812 232784 240968 232812
rect 238812 232772 238818 232784
rect 240962 232772 240968 232784
rect 241020 232812 241026 232824
rect 279602 232812 279608 232824
rect 241020 232784 279608 232812
rect 241020 232772 241026 232784
rect 279602 232772 279608 232784
rect 279660 232772 279666 232824
rect 132494 232704 132500 232756
rect 132552 232744 132558 232756
rect 220078 232744 220084 232756
rect 132552 232716 220084 232744
rect 132552 232704 132558 232716
rect 220078 232704 220084 232716
rect 220136 232704 220142 232756
rect 238478 232704 238484 232756
rect 238536 232744 238542 232756
rect 240686 232744 240692 232756
rect 238536 232716 240692 232744
rect 238536 232704 238542 232716
rect 240686 232704 240692 232716
rect 240744 232704 240750 232756
rect 241238 232704 241244 232756
rect 241296 232744 241302 232756
rect 241422 232744 241428 232756
rect 241296 232716 241428 232744
rect 241296 232704 241302 232716
rect 241422 232704 241428 232716
rect 241480 232744 241486 232756
rect 272794 232744 272800 232756
rect 241480 232716 272800 232744
rect 241480 232704 241486 232716
rect 272794 232704 272800 232716
rect 272852 232704 272858 232756
rect 111794 232636 111800 232688
rect 111852 232676 111858 232688
rect 231302 232676 231308 232688
rect 111852 232648 231308 232676
rect 111852 232636 111858 232648
rect 231302 232636 231308 232648
rect 231360 232636 231366 232688
rect 246390 232636 246396 232688
rect 246448 232676 246454 232688
rect 276934 232676 276940 232688
rect 246448 232648 276940 232676
rect 246448 232636 246454 232648
rect 276934 232636 276940 232648
rect 276992 232636 276998 232688
rect 89714 232568 89720 232620
rect 89772 232608 89778 232620
rect 213546 232608 213552 232620
rect 89772 232580 213552 232608
rect 89772 232568 89778 232580
rect 213546 232568 213552 232580
rect 213604 232568 213610 232620
rect 243906 232568 243912 232620
rect 243964 232608 243970 232620
rect 271874 232608 271880 232620
rect 243964 232580 271880 232608
rect 243964 232568 243970 232580
rect 271874 232568 271880 232580
rect 271932 232568 271938 232620
rect 62758 232500 62764 232552
rect 62816 232540 62822 232552
rect 210970 232540 210976 232552
rect 62816 232512 210976 232540
rect 62816 232500 62822 232512
rect 210970 232500 210976 232512
rect 211028 232500 211034 232552
rect 242526 232500 242532 232552
rect 242584 232540 242590 232552
rect 251082 232540 251088 232552
rect 242584 232512 251088 232540
rect 242584 232500 242590 232512
rect 251082 232500 251088 232512
rect 251140 232540 251146 232552
rect 300302 232540 300308 232552
rect 251140 232512 300308 232540
rect 251140 232500 251146 232512
rect 300302 232500 300308 232512
rect 300360 232500 300366 232552
rect 310422 232500 310428 232552
rect 310480 232540 310486 232552
rect 356054 232540 356060 232552
rect 310480 232512 356060 232540
rect 310480 232500 310486 232512
rect 356054 232500 356060 232512
rect 356112 232500 356118 232552
rect 251174 232432 251180 232484
rect 251232 232472 251238 232484
rect 252370 232472 252376 232484
rect 251232 232444 252376 232472
rect 251232 232432 251238 232444
rect 252370 232432 252376 232444
rect 252428 232472 252434 232484
rect 279786 232472 279792 232484
rect 252428 232444 279792 232472
rect 252428 232432 252434 232444
rect 279786 232432 279792 232444
rect 279844 232432 279850 232484
rect 242710 232364 242716 232416
rect 242768 232404 242774 232416
rect 268378 232404 268384 232416
rect 242768 232376 268384 232404
rect 242768 232364 242774 232376
rect 268378 232364 268384 232376
rect 268436 232364 268442 232416
rect 242250 232296 242256 232348
rect 242308 232336 242314 232348
rect 248322 232336 248328 232348
rect 242308 232308 248328 232336
rect 242308 232296 242314 232308
rect 248322 232296 248328 232308
rect 248380 232336 248386 232348
rect 272886 232336 272892 232348
rect 248380 232308 272892 232336
rect 248380 232296 248386 232308
rect 272886 232296 272892 232308
rect 272944 232296 272950 232348
rect 266078 232228 266084 232280
rect 266136 232268 266142 232280
rect 269390 232268 269396 232280
rect 266136 232240 269396 232268
rect 266136 232228 266142 232240
rect 269390 232228 269396 232240
rect 269448 232228 269454 232280
rect 227714 232160 227720 232212
rect 227772 232200 227778 232212
rect 228726 232200 228732 232212
rect 227772 232172 228732 232200
rect 227772 232160 227778 232172
rect 228726 232160 228732 232172
rect 228784 232160 228790 232212
rect 252186 232160 252192 232212
rect 252244 232200 252250 232212
rect 255314 232200 255320 232212
rect 252244 232172 255320 232200
rect 252244 232160 252250 232172
rect 255314 232160 255320 232172
rect 255372 232160 255378 232212
rect 271874 232160 271880 232212
rect 271932 232200 271938 232212
rect 273162 232200 273168 232212
rect 271932 232172 273168 232200
rect 271932 232160 271938 232172
rect 273162 232160 273168 232172
rect 273220 232200 273226 232212
rect 273898 232200 273904 232212
rect 273220 232172 273904 232200
rect 273220 232160 273226 232172
rect 273898 232160 273904 232172
rect 273956 232160 273962 232212
rect 240318 231888 240324 231940
rect 240376 231928 240382 231940
rect 240870 231928 240876 231940
rect 240376 231900 240876 231928
rect 240376 231888 240382 231900
rect 240870 231888 240876 231900
rect 240928 231888 240934 231940
rect 245654 231820 245660 231872
rect 245712 231860 245718 231872
rect 246390 231860 246396 231872
rect 245712 231832 246396 231860
rect 245712 231820 245718 231832
rect 246390 231820 246396 231832
rect 246448 231820 246454 231872
rect 303706 231820 303712 231872
rect 303764 231860 303770 231872
rect 324590 231860 324596 231872
rect 303764 231832 324596 231860
rect 303764 231820 303770 231832
rect 324590 231820 324596 231832
rect 324648 231820 324654 231872
rect 241790 231752 241796 231804
rect 241848 231792 241854 231804
rect 243630 231792 243636 231804
rect 241848 231764 243636 231792
rect 241848 231752 241854 231764
rect 243630 231752 243636 231764
rect 243688 231752 243694 231804
rect 250162 231752 250168 231804
rect 250220 231792 250226 231804
rect 335814 231792 335820 231804
rect 250220 231764 335820 231792
rect 250220 231752 250226 231764
rect 335814 231752 335820 231764
rect 335872 231792 335878 231804
rect 336642 231792 336648 231804
rect 335872 231764 336648 231792
rect 335872 231752 335878 231764
rect 336642 231752 336648 231764
rect 336700 231752 336706 231804
rect 248874 231684 248880 231736
rect 248932 231724 248938 231736
rect 328822 231724 328828 231736
rect 248932 231696 328828 231724
rect 248932 231684 248938 231696
rect 328822 231684 328828 231696
rect 328880 231724 328886 231736
rect 329190 231724 329196 231736
rect 328880 231696 329196 231724
rect 328880 231684 328886 231696
rect 329190 231684 329196 231696
rect 329248 231684 329254 231736
rect 251358 231616 251364 231668
rect 251416 231656 251422 231668
rect 311250 231656 311256 231668
rect 251416 231628 311256 231656
rect 251416 231616 251422 231628
rect 311250 231616 311256 231628
rect 311308 231616 311314 231668
rect 248046 231548 248052 231600
rect 248104 231588 248110 231600
rect 306558 231588 306564 231600
rect 248104 231560 306564 231588
rect 248104 231548 248110 231560
rect 306558 231548 306564 231560
rect 306616 231588 306622 231600
rect 307570 231588 307576 231600
rect 306616 231560 307576 231588
rect 306616 231548 306622 231560
rect 307570 231548 307576 231560
rect 307628 231548 307634 231600
rect 225230 231480 225236 231532
rect 225288 231520 225294 231532
rect 226058 231520 226064 231532
rect 225288 231492 226064 231520
rect 225288 231480 225294 231492
rect 226058 231480 226064 231492
rect 226116 231480 226122 231532
rect 236546 231480 236552 231532
rect 236604 231520 236610 231532
rect 239306 231520 239312 231532
rect 236604 231492 239312 231520
rect 236604 231480 236610 231492
rect 239306 231480 239312 231492
rect 239364 231520 239370 231532
rect 299014 231520 299020 231532
rect 239364 231492 299020 231520
rect 239364 231480 239370 231492
rect 299014 231480 299020 231492
rect 299072 231480 299078 231532
rect 240410 231412 240416 231464
rect 240468 231452 240474 231464
rect 240778 231452 240784 231464
rect 240468 231424 240784 231452
rect 240468 231412 240474 231424
rect 240778 231412 240784 231424
rect 240836 231452 240842 231464
rect 299842 231452 299848 231464
rect 240836 231424 299848 231452
rect 240836 231412 240842 231424
rect 299842 231412 299848 231424
rect 299900 231412 299906 231464
rect 265250 231344 265256 231396
rect 265308 231384 265314 231396
rect 265308 231356 306374 231384
rect 265308 231344 265314 231356
rect 233234 231276 233240 231328
rect 233292 231316 233298 231328
rect 240594 231316 240600 231328
rect 233292 231288 240600 231316
rect 233292 231276 233298 231288
rect 240594 231276 240600 231288
rect 240652 231316 240658 231328
rect 282546 231316 282552 231328
rect 240652 231288 282552 231316
rect 240652 231276 240658 231288
rect 282546 231276 282552 231288
rect 282604 231276 282610 231328
rect 244826 231208 244832 231260
rect 244884 231248 244890 231260
rect 284202 231248 284208 231260
rect 244884 231220 284208 231248
rect 244884 231208 244890 231220
rect 284202 231208 284208 231220
rect 284260 231208 284266 231260
rect 235994 231140 236000 231192
rect 236052 231180 236058 231192
rect 240870 231180 240876 231192
rect 236052 231152 240876 231180
rect 236052 231140 236058 231152
rect 240870 231140 240876 231152
rect 240928 231180 240934 231192
rect 279694 231180 279700 231192
rect 240928 231152 279700 231180
rect 240928 231140 240934 231152
rect 279694 231140 279700 231152
rect 279752 231140 279758 231192
rect 74534 231072 74540 231124
rect 74592 231112 74598 231124
rect 228910 231112 228916 231124
rect 74592 231084 228916 231112
rect 74592 231072 74598 231084
rect 228910 231072 228916 231084
rect 228968 231072 228974 231124
rect 257062 231072 257068 231124
rect 257120 231112 257126 231124
rect 296714 231112 296720 231124
rect 257120 231084 296720 231112
rect 257120 231072 257126 231084
rect 296714 231072 296720 231084
rect 296772 231112 296778 231124
rect 298002 231112 298008 231124
rect 296772 231084 298008 231112
rect 296772 231072 296778 231084
rect 298002 231072 298008 231084
rect 298060 231072 298066 231124
rect 306346 231112 306374 231356
rect 307570 231140 307576 231192
rect 307628 231180 307634 231192
rect 320174 231180 320180 231192
rect 307628 231152 320180 231180
rect 307628 231140 307634 231152
rect 320174 231140 320180 231152
rect 320232 231140 320238 231192
rect 336642 231140 336648 231192
rect 336700 231180 336706 231192
rect 351178 231180 351184 231192
rect 336700 231152 351184 231180
rect 336700 231140 336706 231152
rect 351178 231140 351184 231152
rect 351236 231140 351242 231192
rect 315758 231112 315764 231124
rect 306346 231084 315764 231112
rect 315758 231072 315764 231084
rect 315816 231112 315822 231124
rect 421558 231112 421564 231124
rect 315816 231084 421564 231112
rect 315816 231072 315822 231084
rect 421558 231072 421564 231084
rect 421616 231072 421622 231124
rect 275554 231044 275560 231056
rect 238312 231016 275560 231044
rect 238312 230988 238340 231016
rect 275554 231004 275560 231016
rect 275612 231004 275618 231056
rect 233878 230936 233884 230988
rect 233936 230976 233942 230988
rect 234062 230976 234068 230988
rect 233936 230948 234068 230976
rect 233936 230936 233942 230948
rect 234062 230936 234068 230948
rect 234120 230936 234126 230988
rect 237650 230936 237656 230988
rect 237708 230976 237714 230988
rect 238294 230976 238300 230988
rect 237708 230948 238300 230976
rect 237708 230936 237714 230948
rect 238294 230936 238300 230948
rect 238352 230936 238358 230988
rect 239950 230936 239956 230988
rect 240008 230976 240014 230988
rect 274358 230976 274364 230988
rect 240008 230948 274364 230976
rect 240008 230936 240014 230948
rect 274358 230936 274364 230948
rect 274416 230936 274422 230988
rect 239398 230868 239404 230920
rect 239456 230908 239462 230920
rect 271598 230908 271604 230920
rect 239456 230880 271604 230908
rect 239456 230868 239462 230880
rect 271598 230868 271604 230880
rect 271656 230868 271662 230920
rect 233694 230732 233700 230784
rect 233752 230772 233758 230784
rect 234522 230772 234528 230784
rect 233752 230744 234528 230772
rect 233752 230732 233758 230744
rect 234522 230732 234528 230744
rect 234580 230732 234586 230784
rect 264054 230732 264060 230784
rect 264112 230772 264118 230784
rect 264882 230772 264888 230784
rect 264112 230744 264888 230772
rect 264112 230732 264118 230744
rect 264882 230732 264888 230744
rect 264940 230732 264946 230784
rect 226426 230596 226432 230648
rect 226484 230636 226490 230648
rect 227254 230636 227260 230648
rect 226484 230608 227260 230636
rect 226484 230596 226490 230608
rect 227254 230596 227260 230608
rect 227312 230596 227318 230648
rect 239490 230460 239496 230512
rect 239548 230500 239554 230512
rect 239950 230500 239956 230512
rect 239548 230472 239956 230500
rect 239548 230460 239554 230472
rect 239950 230460 239956 230472
rect 240008 230460 240014 230512
rect 254302 230460 254308 230512
rect 254360 230500 254366 230512
rect 254762 230500 254768 230512
rect 254360 230472 254768 230500
rect 254360 230460 254366 230472
rect 254762 230460 254768 230472
rect 254820 230460 254826 230512
rect 236730 230392 236736 230444
rect 236788 230432 236794 230444
rect 237282 230432 237288 230444
rect 236788 230404 237288 230432
rect 236788 230392 236794 230404
rect 237282 230392 237288 230404
rect 237340 230392 237346 230444
rect 298002 230392 298008 230444
rect 298060 230432 298066 230444
rect 305362 230432 305368 230444
rect 298060 230404 305368 230432
rect 298060 230392 298066 230404
rect 305362 230392 305368 230404
rect 305420 230392 305426 230444
rect 232682 230324 232688 230376
rect 232740 230364 232746 230376
rect 292666 230364 292672 230376
rect 232740 230336 292672 230364
rect 232740 230324 232746 230336
rect 292666 230324 292672 230336
rect 292724 230324 292730 230376
rect 251450 230256 251456 230308
rect 251508 230296 251514 230308
rect 311250 230296 311256 230308
rect 251508 230268 311256 230296
rect 251508 230256 251514 230268
rect 311250 230256 311256 230268
rect 311308 230296 311314 230308
rect 311618 230296 311624 230308
rect 311308 230268 311624 230296
rect 311308 230256 311314 230268
rect 311618 230256 311624 230268
rect 311676 230256 311682 230308
rect 232866 230188 232872 230240
rect 232924 230228 232930 230240
rect 291654 230228 291660 230240
rect 232924 230200 291660 230228
rect 232924 230188 232930 230200
rect 291654 230188 291660 230200
rect 291712 230188 291718 230240
rect 248414 230120 248420 230172
rect 248472 230160 248478 230172
rect 306098 230160 306104 230172
rect 248472 230132 306104 230160
rect 248472 230120 248478 230132
rect 306098 230120 306104 230132
rect 306156 230120 306162 230172
rect 237282 230052 237288 230104
rect 237340 230092 237346 230104
rect 289262 230092 289268 230104
rect 237340 230064 289268 230092
rect 237340 230052 237346 230064
rect 289262 230052 289268 230064
rect 289320 230052 289326 230104
rect 218146 229984 218152 230036
rect 218204 230024 218210 230036
rect 236546 230024 236552 230036
rect 218204 229996 236552 230024
rect 218204 229984 218210 229996
rect 236546 229984 236552 229996
rect 236604 229984 236610 230036
rect 244458 229984 244464 230036
rect 244516 230024 244522 230036
rect 245194 230024 245200 230036
rect 244516 229996 245200 230024
rect 244516 229984 244522 229996
rect 245194 229984 245200 229996
rect 245252 229984 245258 230036
rect 246114 229984 246120 230036
rect 246172 230024 246178 230036
rect 291838 230024 291844 230036
rect 246172 229996 291844 230024
rect 246172 229984 246178 229996
rect 291838 229984 291844 229996
rect 291896 229984 291902 230036
rect 235534 229916 235540 229968
rect 235592 229956 235598 229968
rect 278314 229956 278320 229968
rect 235592 229928 278320 229956
rect 235592 229916 235598 229928
rect 278314 229916 278320 229928
rect 278372 229916 278378 229968
rect 234982 229848 234988 229900
rect 235040 229888 235046 229900
rect 276842 229888 276848 229900
rect 235040 229860 276848 229888
rect 235040 229848 235046 229860
rect 276842 229848 276848 229860
rect 276900 229848 276906 229900
rect 179414 229780 179420 229832
rect 179472 229820 179478 229832
rect 236362 229820 236368 229832
rect 179472 229792 236368 229820
rect 179472 229780 179478 229792
rect 236362 229780 236368 229792
rect 236420 229820 236426 229832
rect 274174 229820 274180 229832
rect 236420 229792 274180 229820
rect 236420 229780 236426 229792
rect 274174 229780 274180 229792
rect 274232 229780 274238 229832
rect 10318 229712 10324 229764
rect 10376 229752 10382 229764
rect 221918 229752 221924 229764
rect 10376 229724 221924 229752
rect 10376 229712 10382 229724
rect 221918 229712 221924 229724
rect 221976 229712 221982 229764
rect 232590 229712 232596 229764
rect 232648 229752 232654 229764
rect 232958 229752 232964 229764
rect 232648 229724 232964 229752
rect 232648 229712 232654 229724
rect 232958 229712 232964 229724
rect 233016 229712 233022 229764
rect 236638 229712 236644 229764
rect 236696 229752 236702 229764
rect 274266 229752 274272 229764
rect 236696 229724 274272 229752
rect 236696 229712 236702 229724
rect 274266 229712 274272 229724
rect 274324 229712 274330 229764
rect 311250 229712 311256 229764
rect 311308 229752 311314 229764
rect 374086 229752 374092 229764
rect 311308 229724 374092 229752
rect 311308 229712 311314 229724
rect 374086 229712 374092 229724
rect 374144 229712 374150 229764
rect 243078 229644 243084 229696
rect 243136 229684 243142 229696
rect 278774 229684 278780 229696
rect 243136 229656 278780 229684
rect 243136 229644 243142 229656
rect 278774 229644 278780 229656
rect 278832 229644 278838 229696
rect 235902 229576 235908 229628
rect 235960 229616 235966 229628
rect 235960 229588 264376 229616
rect 235960 229576 235966 229588
rect 239122 229508 239128 229560
rect 239180 229548 239186 229560
rect 239180 229520 263732 229548
rect 239180 229508 239186 229520
rect 236270 229440 236276 229492
rect 236328 229480 236334 229492
rect 236328 229452 253934 229480
rect 236328 229440 236334 229452
rect 244366 229372 244372 229424
rect 244424 229412 244430 229424
rect 245286 229412 245292 229424
rect 244424 229384 245292 229412
rect 244424 229372 244430 229384
rect 245286 229372 245292 229384
rect 245344 229372 245350 229424
rect 238018 229304 238024 229356
rect 238076 229344 238082 229356
rect 239122 229344 239128 229356
rect 238076 229316 239128 229344
rect 238076 229304 238082 229316
rect 239122 229304 239128 229316
rect 239180 229304 239186 229356
rect 253906 229276 253934 229452
rect 254118 229440 254124 229492
rect 254176 229480 254182 229492
rect 254578 229480 254584 229492
rect 254176 229452 254584 229480
rect 254176 229440 254182 229452
rect 254578 229440 254584 229452
rect 254636 229440 254642 229492
rect 255774 229440 255780 229492
rect 255832 229480 255838 229492
rect 256510 229480 256516 229492
rect 255832 229452 256516 229480
rect 255832 229440 255838 229452
rect 256510 229440 256516 229452
rect 256568 229440 256574 229492
rect 256694 229440 256700 229492
rect 256752 229480 256758 229492
rect 257706 229480 257712 229492
rect 256752 229452 257712 229480
rect 256752 229440 256758 229452
rect 257706 229440 257712 229452
rect 257764 229440 257770 229492
rect 258258 229440 258264 229492
rect 258316 229480 258322 229492
rect 258902 229480 258908 229492
rect 258316 229452 258908 229480
rect 258316 229440 258322 229452
rect 258902 229440 258908 229452
rect 258960 229440 258966 229492
rect 260834 229440 260840 229492
rect 260892 229480 260898 229492
rect 261386 229480 261392 229492
rect 260892 229452 261392 229480
rect 260892 229440 260898 229452
rect 261386 229440 261392 229452
rect 261444 229440 261450 229492
rect 254026 229372 254032 229424
rect 254084 229412 254090 229424
rect 254854 229412 254860 229424
rect 254084 229384 254860 229412
rect 254084 229372 254090 229384
rect 254854 229372 254860 229384
rect 254912 229372 254918 229424
rect 258074 229372 258080 229424
rect 258132 229412 258138 229424
rect 258626 229412 258632 229424
rect 258132 229384 258632 229412
rect 258132 229372 258138 229384
rect 258626 229372 258632 229384
rect 258684 229372 258690 229424
rect 260926 229372 260932 229424
rect 260984 229412 260990 229424
rect 261570 229412 261576 229424
rect 260984 229384 261576 229412
rect 260984 229372 260990 229384
rect 261570 229372 261576 229384
rect 261628 229372 261634 229424
rect 263704 229412 263732 229520
rect 264348 229480 264376 229588
rect 264422 229576 264428 229628
rect 264480 229616 264486 229628
rect 264698 229616 264704 229628
rect 264480 229588 264704 229616
rect 264480 229576 264486 229588
rect 264698 229576 264704 229588
rect 264756 229576 264762 229628
rect 265526 229576 265532 229628
rect 265584 229616 265590 229628
rect 265986 229616 265992 229628
rect 265584 229588 265992 229616
rect 265584 229576 265590 229588
rect 265986 229576 265992 229588
rect 266044 229576 266050 229628
rect 271414 229480 271420 229492
rect 264348 229452 271420 229480
rect 271414 229440 271420 229452
rect 271472 229440 271478 229492
rect 297082 229480 297088 229492
rect 273226 229452 297088 229480
rect 272702 229412 272708 229424
rect 263704 229384 272708 229412
rect 272702 229372 272708 229384
rect 272760 229372 272766 229424
rect 258166 229304 258172 229356
rect 258224 229344 258230 229356
rect 259270 229344 259276 229356
rect 258224 229316 259276 229344
rect 258224 229304 258230 229316
rect 259270 229304 259276 229316
rect 259328 229304 259334 229356
rect 273226 229276 273254 229452
rect 297082 229440 297088 229452
rect 297140 229440 297146 229492
rect 253906 229248 273254 229276
rect 235074 229168 235080 229220
rect 235132 229208 235138 229220
rect 235902 229208 235908 229220
rect 235132 229180 235908 229208
rect 235132 229168 235138 229180
rect 235902 229168 235908 229180
rect 235960 229168 235966 229220
rect 253934 229168 253940 229220
rect 253992 229208 253998 229220
rect 255130 229208 255136 229220
rect 253992 229180 255136 229208
rect 253992 229168 253998 229180
rect 255130 229168 255136 229180
rect 255188 229168 255194 229220
rect 230842 229100 230848 229152
rect 230900 229140 230906 229152
rect 240042 229140 240048 229152
rect 230900 229112 240048 229140
rect 230900 229100 230906 229112
rect 240042 229100 240048 229112
rect 240100 229100 240106 229152
rect 306098 229100 306104 229152
rect 306156 229140 306162 229152
rect 333974 229140 333980 229152
rect 306156 229112 333980 229140
rect 306156 229100 306162 229112
rect 333974 229100 333980 229112
rect 334032 229100 334038 229152
rect 256878 229032 256884 229084
rect 256936 229072 256942 229084
rect 289354 229072 289360 229084
rect 256936 229044 289360 229072
rect 256936 229032 256942 229044
rect 289354 229032 289360 229044
rect 289412 229032 289418 229084
rect 249242 228964 249248 229016
rect 249300 229004 249306 229016
rect 338574 229004 338580 229016
rect 249300 228976 338580 229004
rect 249300 228964 249306 228976
rect 338574 228964 338580 228976
rect 338632 229004 338638 229016
rect 345014 229004 345020 229016
rect 338632 228976 345020 229004
rect 338632 228964 338638 228976
rect 345014 228964 345020 228976
rect 345072 228964 345078 229016
rect 247678 228896 247684 228948
rect 247736 228936 247742 228948
rect 320542 228936 320548 228948
rect 247736 228908 320548 228936
rect 247736 228896 247742 228908
rect 320542 228896 320548 228908
rect 320600 228896 320606 228948
rect 247034 228828 247040 228880
rect 247092 228868 247098 228880
rect 314930 228868 314936 228880
rect 247092 228840 314936 228868
rect 247092 228828 247098 228840
rect 314930 228828 314936 228840
rect 314988 228828 314994 228880
rect 246850 228760 246856 228812
rect 246908 228800 246914 228812
rect 309410 228800 309416 228812
rect 246908 228772 309416 228800
rect 246908 228760 246914 228772
rect 309410 228760 309416 228772
rect 309468 228760 309474 228812
rect 246022 228692 246028 228744
rect 246080 228732 246086 228744
rect 306466 228732 306472 228744
rect 246080 228704 306472 228732
rect 246080 228692 246086 228704
rect 306466 228692 306472 228704
rect 306524 228692 306530 228744
rect 252830 228624 252836 228676
rect 252888 228664 252894 228676
rect 313090 228664 313096 228676
rect 252888 228636 313096 228664
rect 252888 228624 252894 228636
rect 313090 228624 313096 228636
rect 313148 228624 313154 228676
rect 172514 228556 172520 228608
rect 172572 228596 172578 228608
rect 235074 228596 235080 228608
rect 172572 228568 235080 228596
rect 172572 228556 172578 228568
rect 235074 228556 235080 228568
rect 235132 228556 235138 228608
rect 249150 228556 249156 228608
rect 249208 228596 249214 228608
rect 305638 228596 305644 228608
rect 249208 228568 305644 228596
rect 249208 228556 249214 228568
rect 305638 228556 305644 228568
rect 305696 228556 305702 228608
rect 150434 228488 150440 228540
rect 150492 228528 150498 228540
rect 233878 228528 233884 228540
rect 150492 228500 233884 228528
rect 150492 228488 150498 228500
rect 233878 228488 233884 228500
rect 233936 228488 233942 228540
rect 255958 228488 255964 228540
rect 256016 228528 256022 228540
rect 310514 228528 310520 228540
rect 256016 228500 310520 228528
rect 256016 228488 256022 228500
rect 310514 228488 310520 228500
rect 310572 228488 310578 228540
rect 96614 228420 96620 228472
rect 96672 228460 96678 228472
rect 214650 228460 214656 228472
rect 96672 228432 214656 228460
rect 96672 228420 96678 228432
rect 214650 228420 214656 228432
rect 214708 228420 214714 228472
rect 253290 228420 253296 228472
rect 253348 228460 253354 228472
rect 307938 228460 307944 228472
rect 253348 228432 307944 228460
rect 253348 228420 253354 228432
rect 307938 228420 307944 228432
rect 307996 228420 308002 228472
rect 46934 228352 46940 228404
rect 46992 228392 46998 228404
rect 217870 228392 217876 228404
rect 46992 228364 217876 228392
rect 46992 228352 46998 228364
rect 217870 228352 217876 228364
rect 217928 228352 217934 228404
rect 251910 228352 251916 228404
rect 251968 228392 251974 228404
rect 303614 228392 303620 228404
rect 251968 228364 303620 228392
rect 251968 228352 251974 228364
rect 303614 228352 303620 228364
rect 303672 228352 303678 228404
rect 313090 228352 313096 228404
rect 313148 228392 313154 228404
rect 390646 228392 390652 228404
rect 313148 228364 390652 228392
rect 313148 228352 313154 228364
rect 390646 228352 390652 228364
rect 390704 228352 390710 228404
rect 254670 228284 254676 228336
rect 254728 228324 254734 228336
rect 299566 228324 299572 228336
rect 254728 228296 299572 228324
rect 254728 228284 254734 228296
rect 299566 228284 299572 228296
rect 299624 228284 299630 228336
rect 269850 228256 269856 228268
rect 238726 228228 269856 228256
rect 230750 228080 230756 228132
rect 230808 228120 230814 228132
rect 231302 228120 231308 228132
rect 230808 228092 231308 228120
rect 230808 228080 230814 228092
rect 231302 228080 231308 228092
rect 231360 228120 231366 228132
rect 238726 228120 238754 228228
rect 269850 228216 269856 228228
rect 269908 228216 269914 228268
rect 278774 228216 278780 228268
rect 278832 228256 278838 228268
rect 304074 228256 304080 228268
rect 278832 228228 304080 228256
rect 278832 228216 278838 228228
rect 304074 228216 304080 228228
rect 304132 228216 304138 228268
rect 250070 228148 250076 228200
rect 250128 228188 250134 228200
rect 342254 228188 342260 228200
rect 250128 228160 342260 228188
rect 250128 228148 250134 228160
rect 342254 228148 342260 228160
rect 342312 228148 342318 228200
rect 231360 228092 238754 228120
rect 231360 228080 231366 228092
rect 303614 227944 303620 227996
rect 303672 227984 303678 227996
rect 304258 227984 304264 227996
rect 303672 227956 304264 227984
rect 303672 227944 303678 227956
rect 304258 227944 304264 227956
rect 304316 227944 304322 227996
rect 299566 227740 299572 227792
rect 299624 227780 299630 227792
rect 300210 227780 300216 227792
rect 299624 227752 300216 227780
rect 299624 227740 299630 227752
rect 300210 227740 300216 227752
rect 300268 227740 300274 227792
rect 306466 227740 306472 227792
rect 306524 227780 306530 227792
rect 309134 227780 309140 227792
rect 306524 227752 309140 227780
rect 306524 227740 306530 227752
rect 309134 227740 309140 227752
rect 309192 227740 309198 227792
rect 309410 227740 309416 227792
rect 309468 227780 309474 227792
rect 309870 227780 309876 227792
rect 309468 227752 309876 227780
rect 309468 227740 309474 227752
rect 309870 227740 309876 227752
rect 309928 227740 309934 227792
rect 320542 227740 320548 227792
rect 320600 227780 320606 227792
rect 320818 227780 320824 227792
rect 320600 227752 320824 227780
rect 320600 227740 320606 227752
rect 320818 227740 320824 227752
rect 320876 227740 320882 227792
rect 342254 227740 342260 227792
rect 342312 227780 342318 227792
rect 342898 227780 342904 227792
rect 342312 227752 342904 227780
rect 342312 227740 342318 227752
rect 342898 227740 342904 227752
rect 342956 227740 342962 227792
rect 251726 227672 251732 227724
rect 251784 227712 251790 227724
rect 334158 227712 334164 227724
rect 251784 227684 334164 227712
rect 251784 227672 251790 227684
rect 334158 227672 334164 227684
rect 334216 227712 334222 227724
rect 334526 227712 334532 227724
rect 334216 227684 334532 227712
rect 334216 227672 334222 227684
rect 334526 227672 334532 227684
rect 334584 227672 334590 227724
rect 250438 227604 250444 227656
rect 250496 227644 250502 227656
rect 329926 227644 329932 227656
rect 250496 227616 329932 227644
rect 250496 227604 250502 227616
rect 329926 227604 329932 227616
rect 329984 227604 329990 227656
rect 259178 227536 259184 227588
rect 259236 227576 259242 227588
rect 331306 227576 331312 227588
rect 259236 227548 331312 227576
rect 259236 227536 259242 227548
rect 331306 227536 331312 227548
rect 331364 227536 331370 227588
rect 241330 227468 241336 227520
rect 241388 227508 241394 227520
rect 303982 227508 303988 227520
rect 241388 227480 303988 227508
rect 241388 227468 241394 227480
rect 303982 227468 303988 227480
rect 304040 227468 304046 227520
rect 233050 227400 233056 227452
rect 233108 227440 233114 227452
rect 293126 227440 293132 227452
rect 233108 227412 293132 227440
rect 233108 227400 233114 227412
rect 293126 227400 293132 227412
rect 293184 227400 293190 227452
rect 258534 227332 258540 227384
rect 258592 227372 258598 227384
rect 318518 227372 318524 227384
rect 258592 227344 318524 227372
rect 258592 227332 258598 227344
rect 318518 227332 318524 227344
rect 318576 227332 318582 227384
rect 255314 227264 255320 227316
rect 255372 227304 255378 227316
rect 312722 227304 312728 227316
rect 255372 227276 312728 227304
rect 255372 227264 255378 227276
rect 312722 227264 312728 227276
rect 312780 227264 312786 227316
rect 186314 227196 186320 227248
rect 186372 227236 186378 227248
rect 236638 227236 236644 227248
rect 186372 227208 236644 227236
rect 186372 227196 186378 227208
rect 236638 227196 236644 227208
rect 236696 227196 236702 227248
rect 240318 227196 240324 227248
rect 240376 227236 240382 227248
rect 241330 227236 241336 227248
rect 240376 227208 241336 227236
rect 240376 227196 240382 227208
rect 241330 227196 241336 227208
rect 241388 227196 241394 227248
rect 246758 227196 246764 227248
rect 246816 227236 246822 227248
rect 303246 227236 303252 227248
rect 246816 227208 303252 227236
rect 246816 227196 246822 227208
rect 303246 227196 303252 227208
rect 303304 227196 303310 227248
rect 123478 227128 123484 227180
rect 123536 227168 123542 227180
rect 226518 227168 226524 227180
rect 123536 227140 226524 227168
rect 123536 227128 123542 227140
rect 226518 227128 226524 227140
rect 226576 227128 226582 227180
rect 247310 227128 247316 227180
rect 247368 227168 247374 227180
rect 302050 227168 302056 227180
rect 247368 227140 302056 227168
rect 247368 227128 247374 227140
rect 302050 227128 302056 227140
rect 302108 227128 302114 227180
rect 122098 227060 122104 227112
rect 122156 227100 122162 227112
rect 231026 227100 231032 227112
rect 122156 227072 231032 227100
rect 122156 227060 122162 227072
rect 231026 227060 231032 227072
rect 231084 227060 231090 227112
rect 250806 227060 250812 227112
rect 250864 227100 250870 227112
rect 250990 227100 250996 227112
rect 250864 227072 250996 227100
rect 250864 227060 250870 227072
rect 250990 227060 250996 227072
rect 251048 227060 251054 227112
rect 260650 227060 260656 227112
rect 260708 227100 260714 227112
rect 312906 227100 312912 227112
rect 260708 227072 312912 227100
rect 260708 227060 260714 227072
rect 312906 227060 312912 227072
rect 312964 227060 312970 227112
rect 334158 227060 334164 227112
rect 334216 227100 334222 227112
rect 376018 227100 376024 227112
rect 334216 227072 376024 227100
rect 334216 227060 334222 227072
rect 376018 227060 376024 227072
rect 376076 227060 376082 227112
rect 7650 226992 7656 227044
rect 7708 227032 7714 227044
rect 222930 227032 222936 227044
rect 7708 227004 222936 227032
rect 7708 226992 7714 227004
rect 222930 226992 222936 227004
rect 222988 226992 222994 227044
rect 234154 226992 234160 227044
rect 234212 227032 234218 227044
rect 234212 227004 238754 227032
rect 234212 226992 234218 227004
rect 238726 226964 238754 227004
rect 244550 226992 244556 227044
rect 244608 227032 244614 227044
rect 283006 227032 283012 227044
rect 244608 227004 283012 227032
rect 244608 226992 244614 227004
rect 283006 226992 283012 227004
rect 283064 226992 283070 227044
rect 318518 226992 318524 227044
rect 318576 227032 318582 227044
rect 458174 227032 458180 227044
rect 318576 227004 458180 227032
rect 318576 226992 318582 227004
rect 458174 226992 458180 227004
rect 458232 226992 458238 227044
rect 271322 226964 271328 226976
rect 238726 226936 271328 226964
rect 271322 226924 271328 226936
rect 271380 226924 271386 226976
rect 241054 226856 241060 226908
rect 241112 226896 241118 226908
rect 276750 226896 276756 226908
rect 241112 226868 276756 226896
rect 241112 226856 241118 226868
rect 276750 226856 276756 226868
rect 276808 226856 276814 226908
rect 241698 226788 241704 226840
rect 241756 226828 241762 226840
rect 247034 226828 247040 226840
rect 241756 226800 247040 226828
rect 241756 226788 241762 226800
rect 247034 226788 247040 226800
rect 247092 226828 247098 226840
rect 274082 226828 274088 226840
rect 247092 226800 274088 226828
rect 247092 226788 247098 226800
rect 274082 226788 274088 226800
rect 274140 226788 274146 226840
rect 233694 226652 233700 226704
rect 233752 226692 233758 226704
rect 234154 226692 234160 226704
rect 233752 226664 234160 226692
rect 233752 226652 233758 226664
rect 234154 226652 234160 226664
rect 234212 226652 234218 226704
rect 283006 226380 283012 226432
rect 283064 226420 283070 226432
rect 283742 226420 283748 226432
rect 283064 226392 283748 226420
rect 283064 226380 283070 226392
rect 283742 226380 283748 226392
rect 283800 226380 283806 226432
rect 240134 226312 240140 226364
rect 240192 226352 240198 226364
rect 241054 226352 241060 226364
rect 240192 226324 241060 226352
rect 240192 226312 240198 226324
rect 241054 226312 241060 226324
rect 241112 226312 241118 226364
rect 302050 226312 302056 226364
rect 302108 226352 302114 226364
rect 319438 226352 319444 226364
rect 302108 226324 319444 226352
rect 302108 226312 302114 226324
rect 319438 226312 319444 226324
rect 319496 226312 319502 226364
rect 329926 226312 329932 226364
rect 329984 226352 329990 226364
rect 330570 226352 330576 226364
rect 329984 226324 330576 226352
rect 329984 226312 329990 226324
rect 330570 226312 330576 226324
rect 330628 226312 330634 226364
rect 331306 226312 331312 226364
rect 331364 226352 331370 226364
rect 331950 226352 331956 226364
rect 331364 226324 331956 226352
rect 331364 226312 331370 226324
rect 331950 226312 331956 226324
rect 332008 226312 332014 226364
rect 260190 226244 260196 226296
rect 260248 226284 260254 226296
rect 349246 226284 349252 226296
rect 260248 226256 349252 226284
rect 260248 226244 260254 226256
rect 349246 226244 349252 226256
rect 349304 226244 349310 226296
rect 258442 226176 258448 226228
rect 258500 226216 258506 226228
rect 335538 226216 335544 226228
rect 258500 226188 335544 226216
rect 258500 226176 258506 226188
rect 335538 226176 335544 226188
rect 335596 226216 335602 226228
rect 336090 226216 336096 226228
rect 335596 226188 336096 226216
rect 335596 226176 335602 226188
rect 336090 226176 336096 226188
rect 336148 226176 336154 226228
rect 252738 226108 252744 226160
rect 252796 226148 252802 226160
rect 312814 226148 312820 226160
rect 252796 226120 312820 226148
rect 252796 226108 252802 226120
rect 312814 226108 312820 226120
rect 312872 226108 312878 226160
rect 261202 226040 261208 226092
rect 261260 226080 261266 226092
rect 321186 226080 321192 226092
rect 261260 226052 321192 226080
rect 261260 226040 261266 226052
rect 321186 226040 321192 226052
rect 321244 226040 321250 226092
rect 254210 225972 254216 226024
rect 254268 226012 254274 226024
rect 314010 226012 314016 226024
rect 254268 225984 314016 226012
rect 254268 225972 254274 225984
rect 314010 225972 314016 225984
rect 314068 225972 314074 226024
rect 256970 225904 256976 225956
rect 257028 225944 257034 225956
rect 317138 225944 317144 225956
rect 257028 225916 317144 225944
rect 257028 225904 257034 225916
rect 317138 225904 317144 225916
rect 317196 225944 317202 225956
rect 317322 225944 317328 225956
rect 317196 225916 317328 225944
rect 317196 225904 317202 225916
rect 317322 225904 317328 225916
rect 317380 225904 317386 225956
rect 248598 225836 248604 225888
rect 248656 225876 248662 225888
rect 305270 225876 305276 225888
rect 248656 225848 305276 225876
rect 248656 225836 248662 225848
rect 305270 225836 305276 225848
rect 305328 225836 305334 225888
rect 256142 225768 256148 225820
rect 256200 225808 256206 225820
rect 312538 225808 312544 225820
rect 256200 225780 312544 225808
rect 256200 225768 256206 225780
rect 312538 225768 312544 225780
rect 312596 225768 312602 225820
rect 229370 225700 229376 225752
rect 229428 225740 229434 225752
rect 230014 225740 230020 225752
rect 229428 225712 230020 225740
rect 229428 225700 229434 225712
rect 230014 225700 230020 225712
rect 230072 225700 230078 225752
rect 240042 225700 240048 225752
rect 240100 225740 240106 225752
rect 296162 225740 296168 225752
rect 240100 225712 296168 225740
rect 240100 225700 240106 225712
rect 296162 225700 296168 225712
rect 296220 225700 296226 225752
rect 146294 225632 146300 225684
rect 146352 225672 146358 225684
rect 233970 225672 233976 225684
rect 146352 225644 233976 225672
rect 146352 225632 146358 225644
rect 233970 225632 233976 225644
rect 234028 225632 234034 225684
rect 309778 225632 309784 225684
rect 309836 225672 309842 225684
rect 385678 225672 385684 225684
rect 309836 225644 385684 225672
rect 309836 225632 309842 225644
rect 385678 225632 385684 225644
rect 385736 225632 385742 225684
rect 136634 225564 136640 225616
rect 136692 225604 136698 225616
rect 233050 225604 233056 225616
rect 136692 225576 233056 225604
rect 136692 225564 136698 225576
rect 233050 225564 233056 225576
rect 233108 225564 233114 225616
rect 260374 225564 260380 225616
rect 260432 225604 260438 225616
rect 314838 225604 314844 225616
rect 260432 225576 314844 225604
rect 260432 225564 260438 225576
rect 314838 225564 314844 225576
rect 314896 225564 314902 225616
rect 317322 225564 317328 225616
rect 317380 225604 317386 225616
rect 443638 225604 443644 225616
rect 317380 225576 443644 225604
rect 317380 225564 317386 225576
rect 443638 225564 443644 225576
rect 443696 225564 443702 225616
rect 264330 225496 264336 225548
rect 264388 225536 264394 225548
rect 317966 225536 317972 225548
rect 264388 225508 317972 225536
rect 264388 225496 264394 225508
rect 317966 225496 317972 225508
rect 318024 225536 318030 225548
rect 318702 225536 318708 225548
rect 318024 225508 318708 225536
rect 318024 225496 318030 225508
rect 318702 225496 318708 225508
rect 318760 225496 318766 225548
rect 243538 225428 243544 225480
rect 243596 225468 243602 225480
rect 273254 225468 273260 225480
rect 243596 225440 273260 225468
rect 243596 225428 243602 225440
rect 273254 225428 273260 225440
rect 273312 225428 273318 225480
rect 230014 225360 230020 225412
rect 230072 225400 230078 225412
rect 275830 225400 275836 225412
rect 230072 225372 275836 225400
rect 230072 225360 230078 225372
rect 275830 225360 275836 225372
rect 275888 225360 275894 225412
rect 261662 225292 261668 225344
rect 261720 225332 261726 225344
rect 314286 225332 314292 225344
rect 261720 225304 314292 225332
rect 261720 225292 261726 225304
rect 314286 225292 314292 225304
rect 314344 225292 314350 225344
rect 273254 224952 273260 225004
rect 273312 224992 273318 225004
rect 273990 224992 273996 225004
rect 273312 224964 273996 224992
rect 273312 224952 273318 224964
rect 273990 224952 273996 224964
rect 274048 224952 274054 225004
rect 305270 224952 305276 225004
rect 305328 224992 305334 225004
rect 338114 224992 338120 225004
rect 305328 224964 338120 224992
rect 305328 224952 305334 224964
rect 338114 224952 338120 224964
rect 338172 224952 338178 225004
rect 349246 224952 349252 225004
rect 349304 224992 349310 225004
rect 349798 224992 349804 225004
rect 349304 224964 349804 224992
rect 349304 224952 349310 224964
rect 349798 224952 349804 224964
rect 349856 224952 349862 225004
rect 254762 224884 254768 224936
rect 254820 224924 254826 224936
rect 332778 224924 332784 224936
rect 254820 224896 332784 224924
rect 254820 224884 254826 224896
rect 332778 224884 332784 224896
rect 332836 224924 332842 224936
rect 333054 224924 333060 224936
rect 332836 224896 333060 224924
rect 332836 224884 332842 224896
rect 333054 224884 333060 224896
rect 333112 224884 333118 224936
rect 263686 224816 263692 224868
rect 263744 224856 263750 224868
rect 332870 224856 332876 224868
rect 263744 224828 332876 224856
rect 263744 224816 263750 224828
rect 332870 224816 332876 224828
rect 332928 224816 332934 224868
rect 260926 224748 260932 224800
rect 260984 224788 260990 224800
rect 322474 224788 322480 224800
rect 260984 224760 322480 224788
rect 260984 224748 260990 224760
rect 322474 224748 322480 224760
rect 322532 224748 322538 224800
rect 261018 224680 261024 224732
rect 261076 224720 261082 224732
rect 321002 224720 321008 224732
rect 261076 224692 321008 224720
rect 261076 224680 261082 224692
rect 321002 224680 321008 224692
rect 321060 224680 321066 224732
rect 259914 224612 259920 224664
rect 259972 224652 259978 224664
rect 319530 224652 319536 224664
rect 259972 224624 319536 224652
rect 259972 224612 259978 224624
rect 319530 224612 319536 224624
rect 319588 224612 319594 224664
rect 249978 224544 249984 224596
rect 250036 224584 250042 224596
rect 309318 224584 309324 224596
rect 250036 224556 309324 224584
rect 250036 224544 250042 224556
rect 309318 224544 309324 224556
rect 309376 224584 309382 224596
rect 309376 224556 325694 224584
rect 309376 224544 309382 224556
rect 234890 224476 234896 224528
rect 234948 224516 234954 224528
rect 235626 224516 235632 224528
rect 234948 224488 235632 224516
rect 234948 224476 234954 224488
rect 235626 224476 235632 224488
rect 235684 224516 235690 224528
rect 290550 224516 290556 224528
rect 235684 224488 290556 224516
rect 235684 224476 235690 224488
rect 290550 224476 290556 224488
rect 290608 224476 290614 224528
rect 263134 224408 263140 224460
rect 263192 224448 263198 224460
rect 316770 224448 316776 224460
rect 263192 224420 316776 224448
rect 263192 224408 263198 224420
rect 316770 224408 316776 224420
rect 316828 224408 316834 224460
rect 234798 224340 234804 224392
rect 234856 224380 234862 224392
rect 235534 224380 235540 224392
rect 234856 224352 235540 224380
rect 234856 224340 234862 224352
rect 235534 224340 235540 224352
rect 235592 224380 235598 224392
rect 286594 224380 286600 224392
rect 235592 224352 286600 224380
rect 235592 224340 235598 224352
rect 286594 224340 286600 224352
rect 286652 224340 286658 224392
rect 325666 224380 325694 224556
rect 358814 224380 358820 224392
rect 325666 224352 358820 224380
rect 358814 224340 358820 224352
rect 358872 224340 358878 224392
rect 66898 224272 66904 224324
rect 66956 224312 66962 224324
rect 226334 224312 226340 224324
rect 66956 224284 226340 224312
rect 66956 224272 66962 224284
rect 226334 224272 226340 224284
rect 226392 224272 226398 224324
rect 233510 224272 233516 224324
rect 233568 224312 233574 224324
rect 275462 224312 275468 224324
rect 233568 224284 275468 224312
rect 233568 224272 233574 224284
rect 275462 224272 275468 224284
rect 275520 224272 275526 224324
rect 332778 224272 332784 224324
rect 332836 224312 332842 224324
rect 406378 224312 406384 224324
rect 332836 224284 406384 224312
rect 332836 224272 332842 224284
rect 406378 224272 406384 224284
rect 406436 224272 406442 224324
rect 19978 224204 19984 224256
rect 20036 224244 20042 224256
rect 223574 224244 223580 224256
rect 20036 224216 223580 224244
rect 20036 224204 20042 224216
rect 223574 224204 223580 224216
rect 223632 224204 223638 224256
rect 241514 224204 241520 224256
rect 241572 224244 241578 224256
rect 249518 224244 249524 224256
rect 241572 224216 249524 224244
rect 241572 224204 241578 224216
rect 249518 224204 249524 224216
rect 249576 224244 249582 224256
rect 301406 224244 301412 224256
rect 249576 224216 301412 224244
rect 249576 224204 249582 224216
rect 301406 224204 301412 224216
rect 301464 224204 301470 224256
rect 332870 224204 332876 224256
rect 332928 224244 332934 224256
rect 537478 224244 537484 224256
rect 332928 224216 537484 224244
rect 332928 224204 332934 224216
rect 537478 224204 537484 224216
rect 537536 224204 537542 224256
rect 255498 223524 255504 223576
rect 255556 223564 255562 223576
rect 340966 223564 340972 223576
rect 255556 223536 340972 223564
rect 255556 223524 255562 223536
rect 340966 223524 340972 223536
rect 341024 223564 341030 223576
rect 341518 223564 341524 223576
rect 341024 223536 341524 223564
rect 341024 223524 341030 223536
rect 341518 223524 341524 223536
rect 341576 223524 341582 223576
rect 248506 223456 248512 223508
rect 248564 223496 248570 223508
rect 331214 223496 331220 223508
rect 248564 223468 331220 223496
rect 248564 223456 248570 223468
rect 331214 223456 331220 223468
rect 331272 223496 331278 223508
rect 332042 223496 332048 223508
rect 331272 223468 332048 223496
rect 331272 223456 331278 223468
rect 332042 223456 332048 223468
rect 332100 223456 332106 223508
rect 251266 223388 251272 223440
rect 251324 223428 251330 223440
rect 322934 223428 322940 223440
rect 251324 223400 322940 223428
rect 251324 223388 251330 223400
rect 322934 223388 322940 223400
rect 322992 223388 322998 223440
rect 264606 223320 264612 223372
rect 264664 223360 264670 223372
rect 334250 223360 334256 223372
rect 264664 223332 334256 223360
rect 264664 223320 264670 223332
rect 334250 223320 334256 223332
rect 334308 223360 334314 223372
rect 334802 223360 334808 223372
rect 334308 223332 334808 223360
rect 334308 223320 334314 223332
rect 334802 223320 334808 223332
rect 334860 223320 334866 223372
rect 250990 223252 250996 223304
rect 251048 223292 251054 223304
rect 311342 223292 311348 223304
rect 251048 223264 311348 223292
rect 251048 223252 251054 223264
rect 311342 223252 311348 223264
rect 311400 223252 311406 223304
rect 228358 223184 228364 223236
rect 228416 223224 228422 223236
rect 228818 223224 228824 223236
rect 228416 223196 228824 223224
rect 228416 223184 228422 223196
rect 228818 223184 228824 223196
rect 228876 223224 228882 223236
rect 287606 223224 287612 223236
rect 228876 223196 287612 223224
rect 228876 223184 228882 223196
rect 287606 223184 287612 223196
rect 287664 223184 287670 223236
rect 257798 223116 257804 223168
rect 257856 223156 257862 223168
rect 257856 223128 316034 223156
rect 257856 223116 257862 223128
rect 204254 223048 204260 223100
rect 204312 223088 204318 223100
rect 237650 223088 237656 223100
rect 204312 223060 237656 223088
rect 204312 223048 204318 223060
rect 237650 223048 237656 223060
rect 237708 223048 237714 223100
rect 255130 223048 255136 223100
rect 255188 223088 255194 223100
rect 302878 223088 302884 223100
rect 255188 223060 302884 223088
rect 255188 223048 255194 223060
rect 302878 223048 302884 223060
rect 302936 223048 302942 223100
rect 140774 222980 140780 223032
rect 140832 223020 140838 223032
rect 233418 223020 233424 223032
rect 140832 222992 233424 223020
rect 140832 222980 140838 222992
rect 233418 222980 233424 222992
rect 233476 222980 233482 223032
rect 244090 222980 244096 223032
rect 244148 223020 244154 223032
rect 273162 223020 273168 223032
rect 244148 222992 273168 223020
rect 244148 222980 244154 222992
rect 273162 222980 273168 222992
rect 273220 222980 273226 223032
rect 75914 222912 75920 222964
rect 75972 222952 75978 222964
rect 228358 222952 228364 222964
rect 75972 222924 228364 222952
rect 75972 222912 75978 222924
rect 228358 222912 228364 222924
rect 228416 222912 228422 222964
rect 256878 222912 256884 222964
rect 256936 222952 256942 222964
rect 313274 222952 313280 222964
rect 256936 222924 313280 222952
rect 256936 222912 256942 222924
rect 313274 222912 313280 222924
rect 313332 222912 313338 222964
rect 316006 222952 316034 223128
rect 322934 222980 322940 223032
rect 322992 223020 322998 223032
rect 323578 223020 323584 223032
rect 322992 222992 323584 223020
rect 322992 222980 322998 222992
rect 323578 222980 323584 222992
rect 323636 223020 323642 223032
rect 380894 223020 380900 223032
rect 323636 222992 380900 223020
rect 323636 222980 323642 222992
rect 380894 222980 380900 222992
rect 380952 222980 380958 223032
rect 317046 222952 317052 222964
rect 316006 222924 317052 222952
rect 317046 222912 317052 222924
rect 317104 222952 317110 222964
rect 447778 222952 447784 222964
rect 317104 222924 447784 222952
rect 317104 222912 317110 222924
rect 447778 222912 447784 222924
rect 447836 222912 447842 222964
rect 33134 222844 33140 222896
rect 33192 222884 33198 222896
rect 225046 222884 225052 222896
rect 33192 222856 225052 222884
rect 33192 222844 33198 222856
rect 225046 222844 225052 222856
rect 225104 222844 225110 222896
rect 226610 222844 226616 222896
rect 226668 222884 226674 222896
rect 227070 222884 227076 222896
rect 226668 222856 227076 222884
rect 226668 222844 226674 222856
rect 227070 222844 227076 222856
rect 227128 222884 227134 222896
rect 287422 222884 287428 222896
rect 227128 222856 287428 222884
rect 227128 222844 227134 222856
rect 287422 222844 287428 222856
rect 287480 222844 287486 222896
rect 334802 222844 334808 222896
rect 334860 222884 334866 222896
rect 543734 222884 543740 222896
rect 334860 222856 543740 222884
rect 334860 222844 334866 222856
rect 543734 222844 543740 222856
rect 543792 222844 543798 222896
rect 254394 222776 254400 222828
rect 254452 222816 254458 222828
rect 255130 222816 255136 222828
rect 254452 222788 255136 222816
rect 254452 222776 254458 222788
rect 255130 222776 255136 222788
rect 255188 222816 255194 222828
rect 256878 222816 256884 222828
rect 255188 222788 256884 222816
rect 255188 222776 255194 222788
rect 256878 222776 256884 222788
rect 256936 222776 256942 222828
rect 229278 222096 229284 222148
rect 229336 222136 229342 222148
rect 230106 222136 230112 222148
rect 229336 222108 230112 222136
rect 229336 222096 229342 222108
rect 230106 222096 230112 222108
rect 230164 222096 230170 222148
rect 241146 222096 241152 222148
rect 241204 222136 241210 222148
rect 241514 222136 241520 222148
rect 241204 222108 241520 222136
rect 241204 222096 241210 222108
rect 241514 222096 241520 222108
rect 241572 222096 241578 222148
rect 249886 222096 249892 222148
rect 249944 222136 249950 222148
rect 338482 222136 338488 222148
rect 249944 222108 338488 222136
rect 249944 222096 249950 222108
rect 338482 222096 338488 222108
rect 338540 222136 338546 222148
rect 339402 222136 339408 222148
rect 338540 222108 339408 222136
rect 338540 222096 338546 222108
rect 339402 222096 339408 222108
rect 339460 222096 339466 222148
rect 259638 222028 259644 222080
rect 259696 222068 259702 222080
rect 329834 222068 329840 222080
rect 259696 222040 329840 222068
rect 259696 222028 259702 222040
rect 329834 222028 329840 222040
rect 329892 222068 329898 222080
rect 330294 222068 330300 222080
rect 329892 222040 330300 222068
rect 329892 222028 329898 222040
rect 330294 222028 330300 222040
rect 330352 222028 330358 222080
rect 236086 221960 236092 222012
rect 236144 222000 236150 222012
rect 295702 222000 295708 222012
rect 236144 221972 295708 222000
rect 236144 221960 236150 221972
rect 295702 221960 295708 221972
rect 295760 221960 295766 222012
rect 254118 221892 254124 221944
rect 254176 221932 254182 221944
rect 313274 221932 313280 221944
rect 254176 221904 313280 221932
rect 254176 221892 254182 221904
rect 313274 221892 313280 221904
rect 313332 221892 313338 221944
rect 237558 221824 237564 221876
rect 237616 221864 237622 221876
rect 296070 221864 296076 221876
rect 237616 221836 296076 221864
rect 237616 221824 237622 221836
rect 296070 221824 296076 221836
rect 296128 221824 296134 221876
rect 223850 221756 223856 221808
rect 223908 221796 223914 221808
rect 224126 221796 224132 221808
rect 223908 221768 224132 221796
rect 223908 221756 223914 221768
rect 224126 221756 224132 221768
rect 224184 221796 224190 221808
rect 282362 221796 282368 221808
rect 224184 221768 282368 221796
rect 224184 221756 224190 221768
rect 282362 221756 282368 221768
rect 282420 221756 282426 221808
rect 237190 221688 237196 221740
rect 237248 221728 237254 221740
rect 287882 221728 287888 221740
rect 237248 221700 287888 221728
rect 237248 221688 237254 221700
rect 287882 221688 287888 221700
rect 287940 221688 287946 221740
rect 230106 221620 230112 221672
rect 230164 221660 230170 221672
rect 278222 221660 278228 221672
rect 230164 221632 278228 221660
rect 230164 221620 230170 221632
rect 278222 221620 278228 221632
rect 278280 221620 278286 221672
rect 273162 221552 273168 221604
rect 273220 221592 273226 221604
rect 305178 221592 305184 221604
rect 273220 221564 305184 221592
rect 273220 221552 273226 221564
rect 305178 221552 305184 221564
rect 305236 221552 305242 221604
rect 339402 221552 339408 221604
rect 339460 221592 339466 221604
rect 362954 221592 362960 221604
rect 339460 221564 362960 221592
rect 339460 221552 339466 221564
rect 362954 221552 362960 221564
rect 363012 221552 363018 221604
rect 107654 221484 107660 221536
rect 107712 221524 107718 221536
rect 230474 221524 230480 221536
rect 107712 221496 230480 221524
rect 107712 221484 107718 221496
rect 230474 221484 230480 221496
rect 230532 221484 230538 221536
rect 241514 221484 241520 221536
rect 241572 221524 241578 221536
rect 297358 221524 297364 221536
rect 241572 221496 297364 221524
rect 241572 221484 241578 221496
rect 297358 221484 297364 221496
rect 297416 221484 297422 221536
rect 313274 221484 313280 221536
rect 313332 221524 313338 221536
rect 314470 221524 314476 221536
rect 313332 221496 314476 221524
rect 313332 221484 313338 221496
rect 314470 221484 314476 221496
rect 314528 221524 314534 221536
rect 411898 221524 411904 221536
rect 314528 221496 411904 221524
rect 314528 221484 314534 221496
rect 411898 221484 411904 221496
rect 411956 221484 411962 221536
rect 17954 221416 17960 221468
rect 18012 221456 18018 221468
rect 224126 221456 224132 221468
rect 18012 221428 224132 221456
rect 18012 221416 18018 221428
rect 224126 221416 224132 221428
rect 224184 221416 224190 221468
rect 264606 221416 264612 221468
rect 264664 221456 264670 221468
rect 323762 221456 323768 221468
rect 264664 221428 323768 221456
rect 264664 221416 264670 221428
rect 323762 221416 323768 221428
rect 323820 221416 323826 221468
rect 330294 221416 330300 221468
rect 330352 221456 330358 221468
rect 478138 221456 478144 221468
rect 330352 221428 478144 221456
rect 330352 221416 330358 221428
rect 478138 221416 478144 221428
rect 478196 221416 478202 221468
rect 222378 220736 222384 220788
rect 222436 220776 222442 220788
rect 222930 220776 222936 220788
rect 222436 220748 222936 220776
rect 222436 220736 222442 220748
rect 222930 220736 222936 220748
rect 222988 220736 222994 220788
rect 226978 220736 226984 220788
rect 227036 220776 227042 220788
rect 227254 220776 227260 220788
rect 227036 220748 227260 220776
rect 227036 220736 227042 220748
rect 227254 220736 227260 220748
rect 227312 220736 227318 220788
rect 228082 220736 228088 220788
rect 228140 220776 228146 220788
rect 228542 220776 228548 220788
rect 228140 220748 228548 220776
rect 228140 220736 228146 220748
rect 228542 220736 228548 220748
rect 228600 220736 228606 220788
rect 249794 220736 249800 220788
rect 249852 220776 249858 220788
rect 336826 220776 336832 220788
rect 249852 220748 336832 220776
rect 249852 220736 249858 220748
rect 336826 220736 336832 220748
rect 336884 220776 336890 220788
rect 338022 220776 338028 220788
rect 336884 220748 338028 220776
rect 336884 220736 336890 220748
rect 338022 220736 338028 220748
rect 338080 220736 338086 220788
rect 255406 220668 255412 220720
rect 255464 220708 255470 220720
rect 340874 220708 340880 220720
rect 255464 220680 340880 220708
rect 255464 220668 255470 220680
rect 340874 220668 340880 220680
rect 340932 220668 340938 220720
rect 266538 220600 266544 220652
rect 266596 220640 266602 220652
rect 338666 220640 338672 220652
rect 266596 220612 338672 220640
rect 266596 220600 266602 220612
rect 338666 220600 338672 220612
rect 338724 220640 338730 220652
rect 339402 220640 339408 220652
rect 338724 220612 339408 220640
rect 338724 220600 338730 220612
rect 339402 220600 339408 220612
rect 339460 220600 339466 220652
rect 228174 220532 228180 220584
rect 228232 220572 228238 220584
rect 290274 220572 290280 220584
rect 228232 220544 290280 220572
rect 228232 220532 228238 220544
rect 290274 220532 290280 220544
rect 290332 220532 290338 220584
rect 180794 220464 180800 220516
rect 180852 220504 180858 220516
rect 236086 220504 236092 220516
rect 180852 220476 236092 220504
rect 180852 220464 180858 220476
rect 236086 220464 236092 220476
rect 236144 220464 236150 220516
rect 256418 220464 256424 220516
rect 256476 220504 256482 220516
rect 315850 220504 315856 220516
rect 256476 220476 315856 220504
rect 256476 220464 256482 220476
rect 315850 220464 315856 220476
rect 315908 220464 315914 220516
rect 340874 220464 340880 220516
rect 340932 220504 340938 220516
rect 341610 220504 341616 220516
rect 340932 220476 341616 220504
rect 340932 220464 340938 220476
rect 341610 220464 341616 220476
rect 341668 220464 341674 220516
rect 226334 220396 226340 220448
rect 226392 220436 226398 220448
rect 227162 220436 227168 220448
rect 226392 220408 227168 220436
rect 226392 220396 226398 220408
rect 227162 220396 227168 220408
rect 227220 220436 227226 220448
rect 286318 220436 286324 220448
rect 227220 220408 286324 220436
rect 227220 220396 227226 220408
rect 286318 220396 286324 220408
rect 286376 220396 286382 220448
rect 226978 220328 226984 220380
rect 227036 220368 227042 220380
rect 284938 220368 284944 220380
rect 227036 220340 284944 220368
rect 227036 220328 227042 220340
rect 284938 220328 284944 220340
rect 284996 220328 285002 220380
rect 228542 220260 228548 220312
rect 228600 220300 228606 220312
rect 286410 220300 286416 220312
rect 228600 220272 286416 220300
rect 228600 220260 228606 220272
rect 286410 220260 286416 220272
rect 286468 220260 286474 220312
rect 222930 220192 222936 220244
rect 222988 220232 222994 220244
rect 282914 220232 282920 220244
rect 222988 220204 282920 220232
rect 222988 220192 222994 220204
rect 282914 220192 282920 220204
rect 282972 220192 282978 220244
rect 338022 220192 338028 220244
rect 338080 220232 338086 220244
rect 353938 220232 353944 220244
rect 338080 220204 353944 220232
rect 338080 220192 338086 220204
rect 353938 220192 353944 220204
rect 353996 220192 354002 220244
rect 129734 220124 129740 220176
rect 129792 220164 129798 220176
rect 232958 220164 232964 220176
rect 129792 220136 232964 220164
rect 129792 220124 129798 220136
rect 232958 220124 232964 220136
rect 233016 220124 233022 220176
rect 244550 220124 244556 220176
rect 244608 220164 244614 220176
rect 285582 220164 285588 220176
rect 244608 220136 285588 220164
rect 244608 220124 244614 220136
rect 285582 220124 285588 220136
rect 285640 220124 285646 220176
rect 318702 220124 318708 220176
rect 318760 220164 318766 220176
rect 426434 220164 426440 220176
rect 318760 220136 426440 220164
rect 318760 220124 318766 220136
rect 426434 220124 426440 220136
rect 426492 220124 426498 220176
rect 64874 220056 64880 220108
rect 64932 220096 64938 220108
rect 226334 220096 226340 220108
rect 64932 220068 226340 220096
rect 64932 220056 64938 220068
rect 226334 220056 226340 220068
rect 226392 220056 226398 220108
rect 339402 220056 339408 220108
rect 339460 220096 339466 220108
rect 568574 220096 568580 220108
rect 339460 220068 568580 220096
rect 339460 220056 339466 220068
rect 568574 220056 568580 220068
rect 568632 220056 568638 220108
rect 260834 219376 260840 219428
rect 260892 219416 260898 219428
rect 332686 219416 332692 219428
rect 260892 219388 332692 219416
rect 260892 219376 260898 219388
rect 332686 219376 332692 219388
rect 332744 219376 332750 219428
rect 258350 219308 258356 219360
rect 258408 219348 258414 219360
rect 323394 219348 323400 219360
rect 258408 219320 323400 219348
rect 258408 219308 258414 219320
rect 323394 219308 323400 219320
rect 323452 219308 323458 219360
rect 224310 219240 224316 219292
rect 224368 219280 224374 219292
rect 283558 219280 283564 219292
rect 224368 219252 283564 219280
rect 224368 219240 224374 219252
rect 283558 219240 283564 219252
rect 283616 219240 283622 219292
rect 230290 219172 230296 219224
rect 230348 219212 230354 219224
rect 287698 219212 287704 219224
rect 230348 219184 287704 219212
rect 230348 219172 230354 219184
rect 287698 219172 287704 219184
rect 287756 219172 287762 219224
rect 260742 219104 260748 219156
rect 260800 219144 260806 219156
rect 319990 219144 319996 219156
rect 260800 219116 319996 219144
rect 260800 219104 260806 219116
rect 319990 219104 319996 219116
rect 320048 219104 320054 219156
rect 231578 219036 231584 219088
rect 231636 219076 231642 219088
rect 283650 219076 283656 219088
rect 231636 219048 283656 219076
rect 231636 219036 231642 219048
rect 283650 219036 283656 219048
rect 283708 219036 283714 219088
rect 230198 218968 230204 219020
rect 230256 219008 230262 219020
rect 280890 219008 280896 219020
rect 230256 218980 280896 219008
rect 230256 218968 230262 218980
rect 280890 218968 280896 218980
rect 280948 218968 280954 219020
rect 253474 218900 253480 218952
rect 253532 218940 253538 218952
rect 303430 218940 303436 218952
rect 253532 218912 303436 218940
rect 253532 218900 253538 218912
rect 303430 218900 303436 218912
rect 303488 218900 303494 218952
rect 147674 218832 147680 218884
rect 147732 218872 147738 218884
rect 233326 218872 233332 218884
rect 147732 218844 233332 218872
rect 147732 218832 147738 218844
rect 233326 218832 233332 218844
rect 233384 218832 233390 218884
rect 244458 218832 244464 218884
rect 244516 218872 244522 218884
rect 288342 218872 288348 218884
rect 244516 218844 288348 218872
rect 244516 218832 244522 218844
rect 288342 218832 288348 218844
rect 288400 218832 288406 218884
rect 100754 218764 100760 218816
rect 100812 218804 100818 218816
rect 230290 218804 230296 218816
rect 100812 218776 230296 218804
rect 100812 218764 100818 218776
rect 230290 218764 230296 218776
rect 230348 218764 230354 218816
rect 323394 218764 323400 218816
rect 323452 218804 323458 218816
rect 462314 218804 462320 218816
rect 323452 218776 462320 218804
rect 323452 218764 323458 218776
rect 462314 218764 462320 218776
rect 462372 218764 462378 218816
rect 35894 218696 35900 218748
rect 35952 218736 35958 218748
rect 225414 218736 225420 218748
rect 35952 218708 225420 218736
rect 35952 218696 35958 218708
rect 225414 218696 225420 218708
rect 225472 218696 225478 218748
rect 332686 218696 332692 218748
rect 332744 218736 332750 218748
rect 500954 218736 500960 218748
rect 332744 218708 500960 218736
rect 332744 218696 332750 218708
rect 500954 218696 500960 218708
rect 501012 218696 501018 218748
rect 288342 218016 288348 218068
rect 288400 218056 288406 218068
rect 289078 218056 289084 218068
rect 288400 218028 289084 218056
rect 288400 218016 288406 218028
rect 289078 218016 289084 218028
rect 289136 218016 289142 218068
rect 303430 218016 303436 218068
rect 303488 218056 303494 218068
rect 394694 218056 394700 218068
rect 303488 218028 394700 218056
rect 303488 218016 303494 218028
rect 394694 218016 394700 218028
rect 394752 218016 394758 218068
rect 254026 217948 254032 218000
rect 254084 217988 254090 218000
rect 338298 217988 338304 218000
rect 254084 217960 338304 217988
rect 254084 217948 254090 217960
rect 338298 217948 338304 217960
rect 338356 217948 338362 218000
rect 266814 217880 266820 217932
rect 266872 217920 266878 217932
rect 338390 217920 338396 217932
rect 266872 217892 338396 217920
rect 266872 217880 266878 217892
rect 338390 217880 338396 217892
rect 338448 217880 338454 217932
rect 245838 217812 245844 217864
rect 245896 217852 245902 217864
rect 300118 217852 300124 217864
rect 245896 217824 300124 217852
rect 245896 217812 245902 217824
rect 300118 217812 300124 217824
rect 300176 217812 300182 217864
rect 187694 217472 187700 217524
rect 187752 217512 187758 217524
rect 237190 217512 237196 217524
rect 187752 217484 237196 217512
rect 187752 217472 187758 217484
rect 237190 217472 237196 217484
rect 237248 217472 237254 217524
rect 151814 217404 151820 217456
rect 151872 217444 151878 217456
rect 233970 217444 233976 217456
rect 151872 217416 233976 217444
rect 151872 217404 151878 217416
rect 233970 217404 233976 217416
rect 234028 217404 234034 217456
rect 78674 217336 78680 217388
rect 78732 217376 78738 217388
rect 227990 217376 227996 217388
rect 78732 217348 227996 217376
rect 78732 217336 78738 217348
rect 227990 217336 227996 217348
rect 228048 217336 228054 217388
rect 338298 217336 338304 217388
rect 338356 217376 338362 217388
rect 415394 217376 415400 217388
rect 338356 217348 415400 217376
rect 338356 217336 338362 217348
rect 415394 217336 415400 217348
rect 415452 217336 415458 217388
rect 26234 217268 26240 217320
rect 26292 217308 26298 217320
rect 224310 217308 224316 217320
rect 26292 217280 224316 217308
rect 26292 217268 26298 217280
rect 224310 217268 224316 217280
rect 224368 217268 224374 217320
rect 248230 217268 248236 217320
rect 248288 217308 248294 217320
rect 322934 217308 322940 217320
rect 248288 217280 322940 217308
rect 248288 217268 248294 217280
rect 322934 217268 322940 217280
rect 322992 217268 322998 217320
rect 338390 217268 338396 217320
rect 338448 217308 338454 217320
rect 565078 217308 565084 217320
rect 338448 217280 565084 217308
rect 338448 217268 338454 217280
rect 565078 217268 565084 217280
rect 565136 217268 565142 217320
rect 249334 216588 249340 216640
rect 249392 216628 249398 216640
rect 338206 216628 338212 216640
rect 249392 216600 338212 216628
rect 249392 216588 249398 216600
rect 338206 216588 338212 216600
rect 338264 216628 338270 216640
rect 339402 216628 339408 216640
rect 338264 216600 339408 216628
rect 338264 216588 338270 216600
rect 339402 216588 339408 216600
rect 339460 216588 339466 216640
rect 266446 216520 266452 216572
rect 266504 216560 266510 216572
rect 327166 216560 327172 216572
rect 266504 216532 327172 216560
rect 266504 216520 266510 216532
rect 327166 216520 327172 216532
rect 327224 216560 327230 216572
rect 328362 216560 328368 216572
rect 327224 216532 328368 216560
rect 327224 216520 327230 216532
rect 328362 216520 328368 216532
rect 328420 216520 328426 216572
rect 224862 216452 224868 216504
rect 224920 216492 224926 216504
rect 282178 216492 282184 216504
rect 224920 216464 282184 216492
rect 224920 216452 224926 216464
rect 282178 216452 282184 216464
rect 282236 216452 282242 216504
rect 225046 216112 225052 216164
rect 225104 216152 225110 216164
rect 239582 216152 239588 216164
rect 225104 216124 239588 216152
rect 225104 216112 225110 216124
rect 239582 216112 239588 216124
rect 239640 216112 239646 216164
rect 118694 216044 118700 216096
rect 118752 216084 118758 216096
rect 231578 216084 231584 216096
rect 118752 216056 231584 216084
rect 118752 216044 118758 216056
rect 231578 216044 231584 216056
rect 231636 216044 231642 216096
rect 339402 216044 339408 216096
rect 339460 216084 339466 216096
rect 349246 216084 349252 216096
rect 339460 216056 349252 216084
rect 339460 216044 339466 216056
rect 349246 216044 349252 216056
rect 349304 216044 349310 216096
rect 46198 215976 46204 216028
rect 46256 216016 46262 216028
rect 224954 216016 224960 216028
rect 46256 215988 224960 216016
rect 46256 215976 46262 215988
rect 224954 215976 224960 215988
rect 225012 215976 225018 216028
rect 315850 215976 315856 216028
rect 315908 216016 315914 216028
rect 430574 216016 430580 216028
rect 315908 215988 430580 216016
rect 315908 215976 315914 215988
rect 430574 215976 430580 215988
rect 430632 215976 430638 216028
rect 11054 215908 11060 215960
rect 11112 215948 11118 215960
rect 222194 215948 222200 215960
rect 11112 215920 222200 215948
rect 11112 215908 11118 215920
rect 222194 215908 222200 215920
rect 222252 215908 222258 215960
rect 244182 215908 244188 215960
rect 244240 215948 244246 215960
rect 266354 215948 266360 215960
rect 244240 215920 266360 215948
rect 244240 215908 244246 215920
rect 266354 215908 266360 215920
rect 266412 215908 266418 215960
rect 328362 215908 328368 215960
rect 328420 215948 328426 215960
rect 575474 215948 575480 215960
rect 328420 215920 575480 215948
rect 328420 215908 328426 215920
rect 575474 215908 575480 215920
rect 575532 215908 575538 215960
rect 224310 215296 224316 215348
rect 224368 215336 224374 215348
rect 224862 215336 224868 215348
rect 224368 215308 224868 215336
rect 224368 215296 224374 215308
rect 224862 215296 224868 215308
rect 224920 215296 224926 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 91738 215268 91744 215280
rect 3384 215240 91744 215268
rect 3384 215228 3390 215240
rect 91738 215228 91744 215240
rect 91796 215228 91802 215280
rect 256786 215228 256792 215280
rect 256844 215268 256850 215280
rect 334066 215268 334072 215280
rect 256844 215240 334072 215268
rect 256844 215228 256850 215240
rect 334066 215228 334072 215240
rect 334124 215228 334130 215280
rect 252186 215160 252192 215212
rect 252244 215200 252250 215212
rect 328086 215200 328092 215212
rect 252244 215172 328092 215200
rect 252244 215160 252250 215172
rect 328086 215160 328092 215172
rect 328144 215200 328150 215212
rect 328362 215200 328368 215212
rect 328144 215172 328368 215200
rect 328144 215160 328150 215172
rect 328362 215160 328368 215172
rect 328420 215160 328426 215212
rect 264974 215092 264980 215144
rect 265032 215132 265038 215144
rect 324314 215132 324320 215144
rect 265032 215104 324320 215132
rect 265032 215092 265038 215104
rect 324314 215092 324320 215104
rect 324372 215092 324378 215144
rect 168374 214684 168380 214736
rect 168432 214724 168438 214736
rect 235442 214724 235448 214736
rect 168432 214696 235448 214724
rect 168432 214684 168438 214696
rect 235442 214684 235448 214696
rect 235500 214684 235506 214736
rect 328362 214684 328368 214736
rect 328420 214724 328426 214736
rect 378778 214724 378784 214736
rect 328420 214696 378784 214724
rect 328420 214684 328426 214696
rect 378778 214684 378784 214696
rect 378836 214684 378842 214736
rect 91094 214616 91100 214668
rect 91152 214656 91158 214668
rect 230198 214656 230204 214668
rect 91152 214628 230204 214656
rect 91152 214616 91158 214628
rect 230198 214616 230204 214628
rect 230256 214616 230262 214668
rect 334066 214616 334072 214668
rect 334124 214656 334130 214668
rect 451274 214656 451280 214668
rect 334124 214628 451280 214656
rect 334124 214616 334130 214628
rect 451274 214616 451280 214628
rect 451332 214616 451338 214668
rect 50338 214548 50344 214600
rect 50396 214588 50402 214600
rect 225230 214588 225236 214600
rect 50396 214560 225236 214588
rect 50396 214548 50402 214560
rect 225230 214548 225236 214560
rect 225288 214548 225294 214600
rect 242710 214548 242716 214600
rect 242768 214588 242774 214600
rect 253198 214588 253204 214600
rect 242768 214560 253204 214588
rect 242768 214548 242774 214560
rect 253198 214548 253204 214560
rect 253256 214548 253262 214600
rect 324314 214548 324320 214600
rect 324372 214588 324378 214600
rect 547138 214588 547144 214600
rect 324372 214560 547144 214588
rect 324372 214548 324378 214560
rect 547138 214548 547144 214560
rect 547196 214548 547202 214600
rect 253566 213868 253572 213920
rect 253624 213908 253630 213920
rect 320726 213908 320732 213920
rect 253624 213880 320732 213908
rect 253624 213868 253630 213880
rect 320726 213868 320732 213880
rect 320784 213868 320790 213920
rect 256694 213800 256700 213852
rect 256752 213840 256758 213852
rect 307662 213840 307668 213852
rect 256752 213812 307668 213840
rect 256752 213800 256758 213812
rect 307662 213800 307668 213812
rect 307720 213800 307726 213852
rect 205634 213256 205640 213308
rect 205692 213296 205698 213308
rect 237558 213296 237564 213308
rect 205692 213268 237564 213296
rect 205692 213256 205698 213268
rect 237558 213256 237564 213268
rect 237616 213256 237622 213308
rect 320726 213256 320732 213308
rect 320784 213296 320790 213308
rect 398926 213296 398932 213308
rect 320784 213268 398932 213296
rect 320784 213256 320790 213268
rect 398926 213256 398932 213268
rect 398984 213256 398990 213308
rect 28994 213188 29000 213240
rect 29052 213228 29058 213240
rect 224034 213228 224040 213240
rect 29052 213200 224040 213228
rect 29052 213188 29058 213200
rect 224034 213188 224040 213200
rect 224092 213188 224098 213240
rect 307662 213188 307668 213240
rect 307720 213228 307726 213240
rect 454678 213228 454684 213240
rect 307720 213200 454684 213228
rect 307720 213188 307726 213200
rect 454678 213188 454684 213200
rect 454736 213188 454742 213240
rect 262214 212440 262220 212492
rect 262272 212480 262278 212492
rect 328546 212480 328552 212492
rect 262272 212452 328552 212480
rect 262272 212440 262278 212452
rect 328546 212440 328552 212452
rect 328604 212480 328610 212492
rect 329742 212480 329748 212492
rect 328604 212452 329748 212480
rect 328604 212440 328610 212452
rect 329742 212440 329748 212452
rect 329800 212440 329806 212492
rect 258074 212372 258080 212424
rect 258132 212412 258138 212424
rect 318426 212412 318432 212424
rect 258132 212384 318432 212412
rect 258132 212372 258138 212384
rect 318426 212372 318432 212384
rect 318484 212412 318490 212424
rect 318702 212412 318708 212424
rect 318484 212384 318708 212412
rect 318484 212372 318490 212384
rect 318702 212372 318708 212384
rect 318760 212372 318766 212424
rect 162854 211896 162860 211948
rect 162912 211936 162918 211948
rect 235626 211936 235632 211948
rect 162912 211908 235632 211936
rect 162912 211896 162918 211908
rect 235626 211896 235632 211908
rect 235684 211896 235690 211948
rect 55858 211828 55864 211880
rect 55916 211868 55922 211880
rect 226978 211868 226984 211880
rect 55916 211840 226984 211868
rect 55916 211828 55922 211840
rect 226978 211828 226984 211840
rect 227036 211828 227042 211880
rect 318702 211828 318708 211880
rect 318760 211868 318766 211880
rect 465074 211868 465080 211880
rect 318760 211840 465080 211868
rect 318760 211828 318766 211840
rect 465074 211828 465080 211840
rect 465132 211828 465138 211880
rect 40034 211760 40040 211812
rect 40092 211800 40098 211812
rect 225506 211800 225512 211812
rect 40092 211772 225512 211800
rect 40092 211760 40098 211772
rect 225506 211760 225512 211772
rect 225564 211760 225570 211812
rect 329742 211760 329748 211812
rect 329800 211800 329806 211812
rect 518894 211800 518900 211812
rect 329800 211772 518900 211800
rect 329800 211760 329806 211772
rect 518894 211760 518900 211772
rect 518952 211760 518958 211812
rect 253934 211080 253940 211132
rect 253992 211120 253998 211132
rect 336734 211120 336740 211132
rect 253992 211092 336740 211120
rect 253992 211080 253998 211092
rect 336734 211080 336740 211092
rect 336792 211120 336798 211132
rect 338022 211120 338028 211132
rect 336792 211092 338028 211120
rect 336792 211080 336798 211092
rect 338022 211080 338028 211092
rect 338080 211080 338086 211132
rect 248138 211012 248144 211064
rect 248196 211052 248202 211064
rect 307202 211052 307208 211064
rect 248196 211024 307208 211052
rect 248196 211012 248202 211024
rect 307202 211012 307208 211024
rect 307260 211052 307266 211064
rect 307662 211052 307668 211064
rect 307260 211024 307668 211052
rect 307260 211012 307266 211024
rect 307662 211012 307668 211024
rect 307720 211012 307726 211064
rect 259546 210944 259552 210996
rect 259604 210984 259610 210996
rect 318794 210984 318800 210996
rect 259604 210956 318800 210984
rect 259604 210944 259610 210956
rect 318794 210944 318800 210956
rect 318852 210984 318858 210996
rect 320082 210984 320088 210996
rect 318852 210956 320088 210984
rect 318852 210944 318858 210956
rect 320082 210944 320088 210956
rect 320140 210944 320146 210996
rect 166994 210536 167000 210588
rect 167052 210576 167058 210588
rect 235534 210576 235540 210588
rect 167052 210548 235540 210576
rect 167052 210536 167058 210548
rect 235534 210536 235540 210548
rect 235592 210536 235598 210588
rect 86954 210468 86960 210520
rect 87012 210508 87018 210520
rect 230106 210508 230112 210520
rect 87012 210480 230112 210508
rect 87012 210468 87018 210480
rect 230106 210468 230112 210480
rect 230164 210468 230170 210520
rect 338022 210468 338028 210520
rect 338080 210508 338086 210520
rect 417418 210508 417424 210520
rect 338080 210480 417424 210508
rect 338080 210468 338086 210480
rect 417418 210468 417424 210480
rect 417476 210468 417482 210520
rect 2774 210400 2780 210452
rect 2832 210440 2838 210452
rect 223022 210440 223028 210452
rect 2832 210412 223028 210440
rect 2832 210400 2838 210412
rect 223022 210400 223028 210412
rect 223080 210400 223086 210452
rect 307662 210400 307668 210452
rect 307720 210440 307726 210452
rect 318058 210440 318064 210452
rect 307720 210412 318064 210440
rect 307720 210400 307726 210412
rect 318058 210400 318064 210412
rect 318116 210400 318122 210452
rect 320082 210400 320088 210452
rect 320140 210440 320146 210452
rect 476114 210440 476120 210452
rect 320140 210412 476120 210440
rect 320140 210400 320146 210412
rect 476114 210400 476120 210412
rect 476172 210400 476178 210452
rect 138658 209108 138664 209160
rect 138716 209148 138722 209160
rect 232866 209148 232872 209160
rect 138716 209120 232872 209148
rect 138716 209108 138722 209120
rect 232866 209108 232872 209120
rect 232924 209108 232930 209160
rect 244366 209108 244372 209160
rect 244424 209148 244430 209160
rect 292574 209148 292580 209160
rect 244424 209120 292580 209148
rect 244424 209108 244430 209120
rect 292574 209108 292580 209120
rect 292632 209108 292638 209160
rect 341610 209108 341616 209160
rect 341668 209148 341674 209160
rect 425698 209148 425704 209160
rect 341668 209120 425704 209148
rect 341668 209108 341674 209120
rect 425698 209108 425704 209120
rect 425756 209108 425762 209160
rect 22094 209040 22100 209092
rect 22152 209080 22158 209092
rect 224494 209080 224500 209092
rect 22152 209052 224500 209080
rect 22152 209040 22158 209052
rect 224494 209040 224500 209052
rect 224552 209040 224558 209092
rect 264514 209040 264520 209092
rect 264572 209080 264578 209092
rect 530578 209080 530584 209092
rect 264572 209052 530584 209080
rect 264572 209040 264578 209052
rect 530578 209040 530584 209052
rect 530636 209040 530642 209092
rect 245746 208292 245752 208344
rect 245804 208332 245810 208344
rect 305086 208332 305092 208344
rect 245804 208304 305092 208332
rect 245804 208292 245810 208304
rect 305086 208292 305092 208304
rect 305144 208292 305150 208344
rect 305086 207884 305092 207936
rect 305144 207924 305150 207936
rect 306282 207924 306288 207936
rect 305144 207896 306288 207924
rect 305144 207884 305150 207896
rect 306282 207884 306288 207896
rect 306340 207924 306346 207936
rect 307018 207924 307024 207936
rect 306340 207896 307024 207924
rect 306340 207884 306346 207896
rect 307018 207884 307024 207896
rect 307076 207884 307082 207936
rect 190454 207680 190460 207732
rect 190512 207720 190518 207732
rect 236730 207720 236736 207732
rect 190512 207692 236736 207720
rect 190512 207680 190518 207692
rect 236730 207680 236736 207692
rect 236788 207680 236794 207732
rect 67634 207612 67640 207664
rect 67692 207652 67698 207664
rect 221642 207652 221648 207664
rect 67692 207624 221648 207652
rect 67692 207612 67698 207624
rect 221642 207612 221648 207624
rect 221700 207612 221706 207664
rect 341518 207612 341524 207664
rect 341576 207652 341582 207664
rect 436738 207652 436744 207664
rect 341576 207624 436744 207652
rect 341576 207612 341582 207624
rect 436738 207612 436744 207624
rect 436796 207612 436802 207664
rect 233970 207544 233976 207596
rect 234028 207584 234034 207596
rect 239490 207584 239496 207596
rect 234028 207556 239496 207584
rect 234028 207544 234034 207556
rect 239490 207544 239496 207556
rect 239548 207544 239554 207596
rect 269942 206932 269948 206984
rect 270000 206972 270006 206984
rect 580166 206972 580172 206984
rect 270000 206944 580172 206972
rect 270000 206932 270006 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 201586 206388 201592 206440
rect 201644 206428 201650 206440
rect 237466 206428 237472 206440
rect 201644 206400 237472 206428
rect 201644 206388 201650 206400
rect 237466 206388 237472 206400
rect 237524 206388 237530 206440
rect 155954 206320 155960 206372
rect 156012 206360 156018 206372
rect 234154 206360 234160 206372
rect 156012 206332 234160 206360
rect 156012 206320 156018 206332
rect 234154 206320 234160 206332
rect 234212 206320 234218 206372
rect 55214 206252 55220 206304
rect 55272 206292 55278 206304
rect 226886 206292 226892 206304
rect 55272 206264 226892 206292
rect 55272 206252 55278 206264
rect 226886 206252 226892 206264
rect 226944 206252 226950 206304
rect 258258 205572 258264 205624
rect 258316 205612 258322 205624
rect 328454 205612 328460 205624
rect 258316 205584 328460 205612
rect 258316 205572 258322 205584
rect 328454 205572 328460 205584
rect 328512 205612 328518 205624
rect 329742 205612 329748 205624
rect 328512 205584 329748 205612
rect 328512 205572 328518 205584
rect 329742 205572 329748 205584
rect 329800 205572 329806 205624
rect 265986 205504 265992 205556
rect 266044 205544 266050 205556
rect 324866 205544 324872 205556
rect 266044 205516 324872 205544
rect 266044 205504 266050 205516
rect 324866 205504 324872 205516
rect 324924 205544 324930 205556
rect 325326 205544 325332 205556
rect 324924 205516 325332 205544
rect 324924 205504 324930 205516
rect 325326 205504 325332 205516
rect 325384 205504 325390 205556
rect 121454 204960 121460 205012
rect 121512 205000 121518 205012
rect 231946 205000 231952 205012
rect 121512 204972 231952 205000
rect 121512 204960 121518 204972
rect 231946 204960 231952 204972
rect 232004 204960 232010 205012
rect 329742 204960 329748 205012
rect 329800 205000 329806 205012
rect 461578 205000 461584 205012
rect 329800 204972 461584 205000
rect 329800 204960 329806 204972
rect 461578 204960 461584 204972
rect 461636 204960 461642 205012
rect 80054 204892 80060 204944
rect 80112 204932 80118 204944
rect 228726 204932 228732 204944
rect 80112 204904 228732 204932
rect 80112 204892 80118 204904
rect 228726 204892 228732 204904
rect 228784 204892 228790 204944
rect 324866 204892 324872 204944
rect 324924 204932 324930 204944
rect 553394 204932 553400 204944
rect 324924 204904 553400 204932
rect 324924 204892 324930 204904
rect 553394 204892 553400 204904
rect 553452 204892 553458 204944
rect 258166 204212 258172 204264
rect 258224 204252 258230 204264
rect 335354 204252 335360 204264
rect 258224 204224 335360 204252
rect 258224 204212 258230 204224
rect 335354 204212 335360 204224
rect 335412 204252 335418 204264
rect 336642 204252 336648 204264
rect 335412 204224 336648 204252
rect 335412 204212 335418 204224
rect 336642 204212 336648 204224
rect 336700 204212 336706 204264
rect 8294 203532 8300 203584
rect 8352 203572 8358 203584
rect 222930 203572 222936 203584
rect 8352 203544 222936 203572
rect 8352 203532 8358 203544
rect 222930 203532 222936 203544
rect 222988 203532 222994 203584
rect 336642 203532 336648 203584
rect 336700 203572 336706 203584
rect 472618 203572 472624 203584
rect 336700 203544 472624 203572
rect 336700 203532 336706 203544
rect 472618 203532 472624 203544
rect 472676 203532 472682 203584
rect 21358 202104 21364 202156
rect 21416 202144 21422 202156
rect 222746 202144 222752 202156
rect 21416 202116 222752 202144
rect 21416 202104 21422 202116
rect 222746 202104 222752 202116
rect 222804 202104 222810 202156
rect 126238 200744 126244 200796
rect 126296 200784 126302 200796
rect 232774 200784 232780 200796
rect 126296 200756 232780 200784
rect 126296 200744 126302 200756
rect 232774 200744 232780 200756
rect 232832 200744 232838 200796
rect 31018 199384 31024 199436
rect 31076 199424 31082 199436
rect 223942 199424 223948 199436
rect 31076 199396 223948 199424
rect 31076 199384 31082 199396
rect 223942 199384 223948 199396
rect 224000 199384 224006 199436
rect 165614 198024 165620 198076
rect 165672 198064 165678 198076
rect 235350 198064 235356 198076
rect 165672 198036 235356 198064
rect 165672 198024 165678 198036
rect 235350 198024 235356 198036
rect 235408 198024 235414 198076
rect 65518 197956 65524 198008
rect 65576 197996 65582 198008
rect 227070 197996 227076 198008
rect 65576 197968 227076 197996
rect 65576 197956 65582 197968
rect 227070 197956 227076 197968
rect 227128 197956 227134 198008
rect 176746 196596 176752 196648
rect 176804 196636 176810 196648
rect 236638 196636 236644 196648
rect 176804 196608 236644 196636
rect 176804 196596 176810 196608
rect 236638 196596 236644 196608
rect 236696 196596 236702 196648
rect 249426 196596 249432 196648
rect 249484 196636 249490 196648
rect 340966 196636 340972 196648
rect 249484 196608 340972 196636
rect 249484 196596 249490 196608
rect 340966 196596 340972 196608
rect 341024 196596 341030 196648
rect 75178 195236 75184 195288
rect 75236 195276 75242 195288
rect 228542 195276 228548 195288
rect 75236 195248 228548 195276
rect 75236 195236 75242 195248
rect 228542 195236 228548 195248
rect 228600 195236 228606 195288
rect 250806 195236 250812 195288
rect 250864 195276 250870 195288
rect 357526 195276 357532 195288
rect 250864 195248 357532 195276
rect 250864 195236 250870 195248
rect 357526 195236 357532 195248
rect 357584 195236 357590 195288
rect 39298 193808 39304 193860
rect 39356 193848 39362 193860
rect 225138 193848 225144 193860
rect 39356 193820 225144 193848
rect 39356 193808 39362 193820
rect 225138 193808 225144 193820
rect 225196 193808 225202 193860
rect 577590 193128 577596 193180
rect 577648 193168 577654 193180
rect 579614 193168 579620 193180
rect 577648 193140 579620 193168
rect 577648 193128 577654 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 133874 192516 133880 192568
rect 133932 192556 133938 192568
rect 232682 192556 232688 192568
rect 133932 192528 232688 192556
rect 133932 192516 133938 192528
rect 232682 192516 232688 192528
rect 232740 192516 232746 192568
rect 46290 192448 46296 192500
rect 46348 192488 46354 192500
rect 225782 192488 225788 192500
rect 46348 192460 225788 192488
rect 46348 192448 46354 192460
rect 225782 192448 225788 192460
rect 225840 192448 225846 192500
rect 93946 191088 93952 191140
rect 94004 191128 94010 191140
rect 230014 191128 230020 191140
rect 94004 191100 230020 191128
rect 94004 191088 94010 191100
rect 230014 191088 230020 191100
rect 230072 191088 230078 191140
rect 14458 189728 14464 189780
rect 14516 189768 14522 189780
rect 222654 189768 222660 189780
rect 14516 189740 222660 189768
rect 14516 189728 14522 189740
rect 222654 189728 222660 189740
rect 222712 189728 222718 189780
rect 255038 189728 255044 189780
rect 255096 189768 255102 189780
rect 415486 189768 415492 189780
rect 255096 189740 415492 189768
rect 255096 189728 255102 189740
rect 415486 189728 415492 189740
rect 415544 189728 415550 189780
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 213454 189020 213460 189032
rect 3568 188992 213460 189020
rect 3568 188980 3574 188992
rect 213454 188980 213460 188992
rect 213512 188980 213518 189032
rect 112438 186940 112444 186992
rect 112496 186980 112502 186992
rect 231302 186980 231308 186992
rect 112496 186952 231308 186980
rect 112496 186940 112502 186952
rect 231302 186940 231308 186952
rect 231360 186940 231366 186992
rect 263318 186940 263324 186992
rect 263376 186980 263382 186992
rect 521654 186980 521660 186992
rect 263376 186952 521660 186980
rect 263376 186940 263382 186952
rect 521654 186940 521660 186952
rect 521712 186940 521718 186992
rect 115934 185580 115940 185632
rect 115992 185620 115998 185632
rect 231486 185620 231492 185632
rect 115992 185592 231492 185620
rect 115992 185580 115998 185592
rect 231486 185580 231492 185592
rect 231544 185580 231550 185632
rect 264606 185580 264612 185632
rect 264664 185620 264670 185632
rect 535454 185620 535460 185632
rect 264664 185592 535460 185620
rect 264664 185580 264670 185592
rect 535454 185580 535460 185592
rect 535512 185580 535518 185632
rect 32398 184152 32404 184204
rect 32456 184192 32462 184204
rect 223666 184192 223672 184204
rect 32456 184164 223672 184192
rect 32456 184152 32462 184164
rect 223666 184152 223672 184164
rect 223724 184152 223730 184204
rect 264698 184152 264704 184204
rect 264756 184192 264762 184204
rect 539686 184192 539692 184204
rect 264756 184164 539692 184192
rect 264756 184152 264762 184164
rect 539686 184152 539692 184164
rect 539744 184152 539750 184204
rect 222194 181500 222200 181552
rect 222252 181540 222258 181552
rect 239398 181540 239404 181552
rect 222252 181512 239404 181540
rect 222252 181500 222258 181512
rect 239398 181500 239404 181512
rect 239456 181500 239462 181552
rect 9674 181432 9680 181484
rect 9732 181472 9738 181484
rect 222562 181472 222568 181484
rect 9732 181444 222568 181472
rect 9732 181432 9738 181444
rect 222562 181432 222568 181444
rect 222620 181432 222626 181484
rect 264790 181432 264796 181484
rect 264848 181472 264854 181484
rect 542354 181472 542360 181484
rect 264848 181444 542360 181472
rect 264848 181432 264854 181444
rect 542354 181432 542360 181444
rect 542412 181432 542418 181484
rect 49694 180072 49700 180124
rect 49752 180112 49758 180124
rect 225322 180112 225328 180124
rect 49752 180084 225328 180112
rect 49752 180072 49758 180084
rect 225322 180072 225328 180084
rect 225380 180072 225386 180124
rect 265710 180072 265716 180124
rect 265768 180112 265774 180124
rect 559558 180112 559564 180124
rect 265768 180084 559564 180112
rect 265768 180072 265774 180084
rect 559558 180072 559564 180084
rect 559616 180072 559622 180124
rect 577498 179324 577504 179376
rect 577556 179364 577562 179376
rect 579706 179364 579712 179376
rect 577556 179336 579712 179364
rect 577556 179324 577562 179336
rect 579706 179324 579712 179336
rect 579764 179324 579770 179376
rect 70394 178644 70400 178696
rect 70452 178684 70458 178696
rect 228450 178684 228456 178696
rect 70452 178656 228456 178684
rect 70452 178644 70458 178656
rect 228450 178644 228456 178656
rect 228508 178644 228514 178696
rect 54478 177284 54484 177336
rect 54536 177324 54542 177336
rect 226794 177324 226800 177336
rect 54536 177296 226800 177324
rect 54536 177284 54542 177296
rect 226794 177284 226800 177296
rect 226852 177284 226858 177336
rect 266170 177284 266176 177336
rect 266228 177324 266234 177336
rect 564526 177324 564532 177336
rect 266228 177296 564532 177324
rect 266228 177284 266234 177296
rect 564526 177284 564532 177296
rect 564584 177284 564590 177336
rect 81434 175924 81440 175976
rect 81492 175964 81498 175976
rect 220262 175964 220268 175976
rect 81492 175936 220268 175964
rect 81492 175924 81498 175936
rect 220262 175924 220268 175936
rect 220320 175924 220326 175976
rect 267366 175924 267372 175976
rect 267424 175964 267430 175976
rect 563698 175964 563704 175976
rect 267424 175936 563704 175964
rect 267424 175924 267430 175936
rect 563698 175924 563704 175936
rect 563756 175924 563762 175976
rect 15838 174496 15844 174548
rect 15896 174536 15902 174548
rect 222470 174536 222476 174548
rect 15896 174508 222476 174536
rect 15896 174496 15902 174508
rect 222470 174496 222476 174508
rect 222528 174496 222534 174548
rect 267550 174496 267556 174548
rect 267608 174536 267614 174548
rect 571334 174536 571340 174548
rect 267608 174508 571340 174536
rect 267608 174496 267614 174508
rect 571334 174496 571340 174508
rect 571392 174496 571398 174548
rect 90358 173136 90364 173188
rect 90416 173176 90422 173188
rect 229922 173176 229928 173188
rect 90416 173148 229928 173176
rect 90416 173136 90422 173148
rect 229922 173136 229928 173148
rect 229980 173136 229986 173188
rect 267274 173136 267280 173188
rect 267332 173176 267338 173188
rect 578234 173176 578240 173188
rect 267332 173148 578240 173176
rect 267332 173136 267338 173148
rect 578234 173136 578240 173148
rect 578292 173136 578298 173188
rect 85666 171776 85672 171828
rect 85724 171816 85730 171828
rect 220170 171816 220176 171828
rect 85724 171788 220176 171816
rect 85724 171776 85730 171788
rect 220170 171776 220176 171788
rect 220228 171776 220234 171828
rect 255130 171776 255136 171828
rect 255188 171816 255194 171828
rect 411254 171816 411260 171828
rect 255188 171788 411260 171816
rect 255188 171776 255194 171788
rect 411254 171776 411260 171788
rect 411312 171776 411318 171828
rect 97258 170348 97264 170400
rect 97316 170388 97322 170400
rect 229830 170388 229836 170400
rect 97316 170360 229836 170388
rect 97316 170348 97322 170360
rect 229830 170348 229836 170360
rect 229888 170348 229894 170400
rect 267642 170348 267648 170400
rect 267700 170388 267706 170400
rect 574094 170388 574100 170400
rect 267700 170360 574100 170388
rect 267700 170348 267706 170360
rect 574094 170348 574100 170360
rect 574152 170348 574158 170400
rect 19334 168988 19340 169040
rect 19392 169028 19398 169040
rect 218974 169028 218980 169040
rect 19392 169000 218980 169028
rect 19392 168988 19398 169000
rect 218974 168988 218980 169000
rect 219032 168988 219038 169040
rect 31754 167628 31760 167680
rect 31812 167668 31818 167680
rect 224402 167668 224408 167680
rect 31812 167640 224408 167668
rect 31812 167628 31818 167640
rect 224402 167628 224408 167640
rect 224460 167628 224466 167680
rect 137278 166268 137284 166320
rect 137336 166308 137342 166320
rect 232590 166308 232596 166320
rect 137336 166280 232596 166308
rect 137336 166268 137342 166280
rect 232590 166268 232596 166280
rect 232648 166268 232654 166320
rect 35986 164840 35992 164892
rect 36044 164880 36050 164892
rect 215294 164880 215300 164892
rect 36044 164852 215300 164880
rect 36044 164840 36050 164852
rect 215294 164840 215300 164852
rect 215352 164840 215358 164892
rect 250898 164840 250904 164892
rect 250956 164880 250962 164892
rect 361574 164880 361580 164892
rect 250956 164852 361580 164880
rect 250956 164840 250962 164852
rect 361574 164840 361580 164852
rect 361632 164840 361638 164892
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 199378 164200 199384 164212
rect 3292 164172 199384 164200
rect 3292 164160 3298 164172
rect 199378 164160 199384 164172
rect 199436 164160 199442 164212
rect 155310 162120 155316 162172
rect 155368 162160 155374 162172
rect 234062 162160 234068 162172
rect 155368 162132 234068 162160
rect 155368 162120 155374 162132
rect 234062 162120 234068 162132
rect 234120 162120 234126 162172
rect 241606 162120 241612 162172
rect 241664 162160 241670 162172
rect 251266 162160 251272 162172
rect 241664 162132 251272 162160
rect 241664 162120 241670 162132
rect 251266 162120 251272 162132
rect 251324 162120 251330 162172
rect 42794 160692 42800 160744
rect 42852 160732 42858 160744
rect 206370 160732 206376 160744
rect 42852 160704 206376 160732
rect 42852 160692 42858 160704
rect 206370 160692 206376 160704
rect 206428 160692 206434 160744
rect 79318 159332 79324 159384
rect 79376 159372 79382 159384
rect 228358 159372 228364 159384
rect 79376 159344 228364 159372
rect 79376 159332 79382 159344
rect 228358 159332 228364 159344
rect 228416 159332 228422 159384
rect 127066 157972 127072 158024
rect 127124 158012 127130 158024
rect 232498 158012 232504 158024
rect 127124 157984 232504 158012
rect 127124 157972 127130 157984
rect 232498 157972 232504 157984
rect 232556 157972 232562 158024
rect 53834 155184 53840 155236
rect 53892 155224 53898 155236
rect 227346 155224 227352 155236
rect 53892 155196 227352 155224
rect 53892 155184 53898 155196
rect 227346 155184 227352 155196
rect 227404 155184 227410 155236
rect 334618 153144 334624 153196
rect 334676 153184 334682 153196
rect 580166 153184 580172 153196
rect 334676 153156 580172 153184
rect 334676 153144 334682 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 257982 149676 257988 149728
rect 258040 149716 258046 149728
rect 454034 149716 454040 149728
rect 258040 149688 454040 149716
rect 258040 149676 258046 149688
rect 454034 149676 454040 149688
rect 454092 149676 454098 149728
rect 260742 145528 260748 145580
rect 260800 145568 260806 145580
rect 478874 145568 478880 145580
rect 260800 145540 478880 145568
rect 260800 145528 260806 145540
rect 478874 145528 478880 145540
rect 478932 145528 478938 145580
rect 263410 144168 263416 144220
rect 263468 144208 263474 144220
rect 511994 144208 512000 144220
rect 263468 144180 512000 144208
rect 263468 144168 263474 144180
rect 511994 144168 512000 144180
rect 512052 144168 512058 144220
rect 263502 141380 263508 141432
rect 263560 141420 263566 141432
rect 519538 141420 519544 141432
rect 263560 141392 519544 141420
rect 263560 141380 263566 141392
rect 519538 141380 519544 141392
rect 519596 141380 519602 141432
rect 2866 137912 2872 137964
rect 2924 137952 2930 137964
rect 203518 137952 203524 137964
rect 2924 137924 203524 137952
rect 2924 137912 2930 137924
rect 203518 137912 203524 137924
rect 203576 137912 203582 137964
rect 266262 137232 266268 137284
rect 266320 137272 266326 137284
rect 555510 137272 555516 137284
rect 266320 137244 555516 137272
rect 266320 137232 266326 137244
rect 555510 137232 555516 137244
rect 555568 137232 555574 137284
rect 222010 126216 222016 126268
rect 222068 126256 222074 126268
rect 580350 126256 580356 126268
rect 222068 126228 580356 126256
rect 222068 126216 222074 126228
rect 580350 126216 580356 126228
rect 580408 126216 580414 126268
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 211798 111772 211804 111784
rect 3476 111744 211804 111772
rect 3476 111732 3482 111744
rect 211798 111732 211804 111744
rect 211856 111732 211862 111784
rect 280062 100648 280068 100700
rect 280120 100688 280126 100700
rect 579614 100688 579620 100700
rect 280120 100660 579620 100688
rect 280120 100648 280126 100660
rect 579614 100648 579620 100660
rect 579672 100648 579678 100700
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 197998 97968 198004 97980
rect 3476 97940 198004 97968
rect 3476 97928 3482 97940
rect 197998 97928 198004 97940
rect 198056 97928 198062 97980
rect 11146 90312 11152 90364
rect 11204 90352 11210 90364
rect 209038 90352 209044 90364
rect 11204 90324 209044 90352
rect 11204 90312 11210 90324
rect 209038 90312 209044 90324
rect 209096 90312 209102 90364
rect 222102 87592 222108 87644
rect 222160 87632 222166 87644
rect 580258 87632 580264 87644
rect 222160 87604 580264 87632
rect 222160 87592 222166 87604
rect 580258 87592 580264 87604
rect 580316 87592 580322 87644
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 192478 85524 192484 85536
rect 3200 85496 192484 85524
rect 3200 85484 3206 85496
rect 192478 85484 192484 85496
rect 192536 85484 192542 85536
rect 331858 73108 331864 73160
rect 331916 73148 331922 73160
rect 580166 73148 580172 73160
rect 331916 73120 580172 73148
rect 331916 73108 331922 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 186958 71720 186964 71732
rect 3476 71692 186964 71720
rect 3476 71680 3482 71692
rect 186958 71680 186964 71692
rect 187016 71680 187022 71732
rect 280798 60664 280804 60716
rect 280856 60704 280862 60716
rect 580166 60704 580172 60716
rect 280856 60676 580172 60704
rect 280856 60664 280862 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 195238 59344 195244 59356
rect 3108 59316 195244 59344
rect 3108 59304 3114 59316
rect 195238 59304 195244 59316
rect 195296 59304 195302 59356
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 206278 45540 206284 45552
rect 3476 45512 206284 45540
rect 3476 45500 3482 45512
rect 206278 45500 206284 45512
rect 206336 45500 206342 45552
rect 242802 33736 242808 33788
rect 242860 33776 242866 33788
rect 255314 33776 255320 33788
rect 242860 33748 255320 33776
rect 242860 33736 242866 33748
rect 255314 33736 255320 33748
rect 255372 33736 255378 33788
rect 3418 32988 3424 33040
rect 3476 33028 3482 33040
rect 7558 33028 7564 33040
rect 3476 33000 7564 33028
rect 3476 32988 3482 33000
rect 7558 32988 7564 33000
rect 7616 32988 7622 33040
rect 264882 29588 264888 29640
rect 264940 29628 264946 29640
rect 527818 29628 527824 29640
rect 264940 29600 527824 29628
rect 264940 29588 264946 29600
rect 527818 29588 527824 29600
rect 527876 29588 527882 29640
rect 19426 24080 19432 24132
rect 19484 24120 19490 24132
rect 188338 24120 188344 24132
rect 19484 24092 188344 24120
rect 19484 24080 19490 24092
rect 188338 24080 188344 24092
rect 188396 24080 188402 24132
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 222838 22760 222844 22772
rect 15252 22732 222844 22760
rect 15252 22720 15258 22732
rect 222838 22720 222844 22732
rect 222896 22720 222902 22772
rect 27614 21360 27620 21412
rect 27672 21400 27678 21412
rect 213362 21400 213368 21412
rect 27672 21372 213368 21400
rect 27672 21360 27678 21372
rect 213362 21360 213368 21372
rect 213420 21360 213426 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 43438 20652 43444 20664
rect 3476 20624 43444 20652
rect 3476 20612 3482 20624
rect 43438 20612 43444 20624
rect 43496 20612 43502 20664
rect 418798 20612 418804 20664
rect 418856 20652 418862 20664
rect 580166 20652 580172 20664
rect 418856 20624 580172 20652
rect 418856 20612 418862 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 214558 18612 214564 18624
rect 23532 18584 214564 18612
rect 23532 18572 23538 18584
rect 214558 18572 214564 18584
rect 214616 18572 214622 18624
rect 99374 17212 99380 17264
rect 99432 17252 99438 17264
rect 217410 17252 217416 17264
rect 99432 17224 217416 17252
rect 99432 17212 99438 17224
rect 217410 17212 217416 17224
rect 217468 17212 217474 17264
rect 149514 14424 149520 14476
rect 149572 14464 149578 14476
rect 233878 14464 233884 14476
rect 149572 14436 233884 14464
rect 149572 14424 149578 14436
rect 233878 14424 233884 14436
rect 233936 14424 233942 14476
rect 255222 14424 255228 14476
rect 255280 14464 255286 14476
rect 422570 14464 422576 14476
rect 255280 14436 422576 14464
rect 255280 14424 255286 14436
rect 422570 14424 422576 14436
rect 422628 14424 422634 14476
rect 25314 13064 25320 13116
rect 25372 13104 25378 13116
rect 224126 13104 224132 13116
rect 25372 13076 224132 13104
rect 25372 13064 25378 13076
rect 224126 13064 224132 13076
rect 224184 13064 224190 13116
rect 126974 11772 126980 11824
rect 127032 11812 127038 11824
rect 128170 11812 128176 11824
rect 127032 11784 128176 11812
rect 127032 11772 127038 11784
rect 128170 11772 128176 11784
rect 128228 11772 128234 11824
rect 176654 11772 176660 11824
rect 176712 11812 176718 11824
rect 177850 11812 177856 11824
rect 176712 11784 177856 11812
rect 176712 11772 176718 11784
rect 177850 11772 177856 11784
rect 177908 11772 177914 11824
rect 201494 11772 201500 11824
rect 201552 11812 201558 11824
rect 202690 11812 202696 11824
rect 201552 11784 202696 11812
rect 201552 11772 201558 11784
rect 202690 11772 202696 11784
rect 202748 11772 202754 11824
rect 39114 11704 39120 11756
rect 39172 11744 39178 11756
rect 224310 11744 224316 11756
rect 39172 11716 224316 11744
rect 39172 11704 39178 11716
rect 224310 11704 224316 11716
rect 224368 11704 224374 11756
rect 110506 10276 110512 10328
rect 110564 10316 110570 10328
rect 230934 10316 230940 10328
rect 110564 10288 230940 10316
rect 110564 10276 110570 10288
rect 230934 10276 230940 10288
rect 230992 10276 230998 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 84470 8916 84476 8968
rect 84528 8956 84534 8968
rect 227806 8956 227812 8968
rect 84528 8928 227812 8956
rect 84528 8916 84534 8928
rect 227806 8916 227812 8928
rect 227864 8916 227870 8968
rect 250990 8916 250996 8968
rect 251048 8956 251054 8968
rect 369394 8956 369400 8968
rect 251048 8928 369400 8956
rect 251048 8916 251054 8928
rect 369394 8916 369400 8928
rect 369452 8916 369458 8968
rect 103330 7556 103336 7608
rect 103388 7596 103394 7608
rect 229738 7596 229744 7608
rect 103388 7568 229744 7596
rect 103388 7556 103394 7568
rect 229738 7556 229744 7568
rect 229796 7556 229802 7608
rect 249610 7556 249616 7608
rect 249668 7596 249674 7608
rect 344554 7596 344560 7608
rect 249668 7568 344560 7596
rect 249668 7556 249674 7568
rect 344554 7556 344560 7568
rect 344612 7556 344618 7608
rect 355318 7556 355324 7608
rect 355376 7596 355382 7608
rect 474550 7596 474556 7608
rect 355376 7568 474556 7596
rect 355376 7556 355382 7568
rect 474550 7556 474556 7568
rect 474608 7556 474614 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 116578 6848 116584 6860
rect 3476 6820 116584 6848
rect 3476 6808 3482 6820
rect 116578 6808 116584 6820
rect 116636 6808 116642 6860
rect 336090 6468 336096 6520
rect 336148 6508 336154 6520
rect 460382 6508 460388 6520
rect 336148 6480 460388 6508
rect 336148 6468 336154 6480
rect 460382 6468 460388 6480
rect 460440 6468 460446 6520
rect 252646 6400 252652 6452
rect 252704 6440 252710 6452
rect 394234 6440 394240 6452
rect 252704 6412 394240 6440
rect 252704 6400 252710 6412
rect 394234 6400 394240 6412
rect 394292 6400 394298 6452
rect 253842 6332 253848 6384
rect 253900 6372 253906 6384
rect 397730 6372 397736 6384
rect 253900 6344 397736 6372
rect 253900 6332 253906 6344
rect 397730 6332 397736 6344
rect 397788 6332 397794 6384
rect 256510 6264 256516 6316
rect 256568 6304 256574 6316
rect 429654 6304 429660 6316
rect 256568 6276 429660 6304
rect 256568 6264 256574 6276
rect 429654 6264 429660 6276
rect 429712 6264 429718 6316
rect 256602 6196 256608 6248
rect 256660 6236 256666 6248
rect 433242 6236 433248 6248
rect 256660 6208 433248 6236
rect 256660 6196 256666 6208
rect 433242 6196 433248 6208
rect 433300 6196 433306 6248
rect 117590 6128 117596 6180
rect 117648 6168 117654 6180
rect 231118 6168 231124 6180
rect 117648 6140 231124 6168
rect 117648 6128 117654 6140
rect 231118 6128 231124 6140
rect 231176 6128 231182 6180
rect 259362 6128 259368 6180
rect 259420 6168 259426 6180
rect 461578 6168 461584 6180
rect 259420 6140 461584 6168
rect 259420 6128 259426 6140
rect 461578 6128 461584 6140
rect 461636 6128 461642 6180
rect 475378 5516 475384 5568
rect 475436 5556 475442 5568
rect 478046 5556 478052 5568
rect 475436 5528 478052 5556
rect 475436 5516 475442 5528
rect 478046 5516 478052 5528
rect 478104 5516 478110 5568
rect 78582 4768 78588 4820
rect 78640 4808 78646 4820
rect 227898 4808 227904 4820
rect 78640 4780 227904 4808
rect 78640 4768 78646 4780
rect 227898 4768 227904 4780
rect 227956 4768 227962 4820
rect 349798 4768 349804 4820
rect 349856 4808 349862 4820
rect 449802 4808 449808 4820
rect 349856 4780 449808 4808
rect 349856 4768 349862 4780
rect 449802 4768 449808 4780
rect 449860 4768 449866 4820
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 46198 4128 46204 4140
rect 45520 4100 46204 4128
rect 45520 4088 45526 4100
rect 46198 4088 46204 4100
rect 46256 4088 46262 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 199102 4088 199108 4140
rect 199160 4128 199166 4140
rect 216122 4128 216128 4140
rect 199160 4100 216128 4128
rect 199160 4088 199166 4100
rect 216122 4088 216128 4100
rect 216180 4088 216186 4140
rect 248322 4088 248328 4140
rect 248380 4128 248386 4140
rect 249978 4128 249984 4140
rect 248380 4100 249984 4128
rect 248380 4088 248386 4100
rect 249978 4088 249984 4100
rect 250036 4088 250042 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 318518 4128 318524 4140
rect 315356 4100 318524 4128
rect 315356 4088 315362 4100
rect 318518 4088 318524 4100
rect 318576 4088 318582 4140
rect 330570 4088 330576 4140
rect 330628 4128 330634 4140
rect 336274 4128 336280 4140
rect 330628 4100 336280 4128
rect 330628 4088 330634 4100
rect 336274 4088 336280 4100
rect 336332 4088 336338 4140
rect 353938 4088 353944 4140
rect 353996 4128 354002 4140
rect 353996 4100 354674 4128
rect 353996 4088 354002 4100
rect 193306 4020 193312 4072
rect 193364 4060 193370 4072
rect 213270 4060 213276 4072
rect 193364 4032 213276 4060
rect 193364 4020 193370 4032
rect 213270 4020 213276 4032
rect 213328 4020 213334 4072
rect 251082 4020 251088 4072
rect 251140 4060 251146 4072
rect 260650 4060 260656 4072
rect 251140 4032 260656 4060
rect 251140 4020 251146 4032
rect 260650 4020 260656 4032
rect 260708 4020 260714 4072
rect 275922 4020 275928 4072
rect 275980 4060 275986 4072
rect 278314 4060 278320 4072
rect 275980 4032 278320 4060
rect 275980 4020 275986 4032
rect 278314 4020 278320 4032
rect 278372 4020 278378 4072
rect 329190 4020 329196 4072
rect 329248 4060 329254 4072
rect 329248 4032 331720 4060
rect 329248 4020 329254 4032
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 7650 3992 7656 4004
rect 2924 3964 7656 3992
rect 2924 3952 2930 3964
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 92750 3952 92756 4004
rect 92808 3992 92814 4004
rect 95878 3992 95884 4004
rect 92808 3964 95884 3992
rect 92808 3952 92814 3964
rect 95878 3952 95884 3964
rect 95936 3952 95942 4004
rect 171962 3952 171968 4004
rect 172020 3992 172026 4004
rect 215938 3992 215944 4004
rect 172020 3964 215944 3992
rect 172020 3952 172026 3964
rect 215938 3952 215944 3964
rect 215996 3952 216002 4004
rect 244918 3952 244924 4004
rect 244976 3992 244982 4004
rect 257062 3992 257068 4004
rect 244976 3964 257068 3992
rect 244976 3952 244982 3964
rect 257062 3952 257068 3964
rect 257120 3952 257126 4004
rect 279418 3952 279424 4004
rect 279476 3992 279482 4004
rect 288986 3992 288992 4004
rect 279476 3964 288992 3992
rect 279476 3952 279482 3964
rect 288986 3952 288992 3964
rect 289044 3952 289050 4004
rect 319438 3952 319444 4004
rect 319496 3992 319502 4004
rect 331582 3992 331588 4004
rect 319496 3964 331588 3992
rect 319496 3952 319502 3964
rect 331582 3952 331588 3964
rect 331640 3952 331646 4004
rect 331692 3992 331720 4032
rect 331950 4020 331956 4072
rect 332008 4060 332014 4072
rect 335906 4060 335912 4072
rect 332008 4032 335912 4060
rect 332008 4020 332014 4032
rect 335906 4020 335912 4032
rect 335964 4020 335970 4072
rect 335998 4020 336004 4072
rect 336056 4060 336062 4072
rect 336056 4032 340092 4060
rect 336056 4020 336062 4032
rect 339862 3992 339868 4004
rect 331692 3964 339868 3992
rect 339862 3952 339868 3964
rect 339920 3952 339926 4004
rect 340064 3992 340092 4032
rect 342898 4020 342904 4072
rect 342956 4060 342962 4072
rect 354030 4060 354036 4072
rect 342956 4032 354036 4060
rect 342956 4020 342962 4032
rect 354030 4020 354036 4032
rect 354088 4020 354094 4072
rect 354646 4060 354674 4100
rect 378778 4088 378784 4140
rect 378836 4128 378842 4140
rect 384758 4128 384764 4140
rect 378836 4100 384764 4128
rect 378836 4088 378842 4100
rect 384758 4088 384764 4100
rect 384816 4088 384822 4140
rect 411990 4088 411996 4140
rect 412048 4128 412054 4140
rect 413094 4128 413100 4140
rect 412048 4100 413100 4128
rect 412048 4088 412054 4100
rect 413094 4088 413100 4100
rect 413152 4088 413158 4140
rect 425698 4088 425704 4140
rect 425756 4128 425762 4140
rect 434438 4128 434444 4140
rect 425756 4100 434444 4128
rect 425756 4088 425762 4100
rect 434438 4088 434444 4100
rect 434496 4088 434502 4140
rect 478138 4088 478144 4140
rect 478196 4128 478202 4140
rect 480530 4128 480536 4140
rect 478196 4100 480536 4128
rect 478196 4088 478202 4100
rect 480530 4088 480536 4100
rect 480588 4088 480594 4140
rect 508498 4088 508504 4140
rect 508556 4128 508562 4140
rect 510062 4128 510068 4140
rect 508556 4100 510068 4128
rect 508556 4088 508562 4100
rect 510062 4088 510068 4100
rect 510120 4088 510126 4140
rect 527818 4088 527824 4140
rect 527876 4128 527882 4140
rect 530118 4128 530124 4140
rect 527876 4100 530124 4128
rect 527876 4088 527882 4100
rect 530118 4088 530124 4100
rect 530176 4088 530182 4140
rect 367002 4060 367008 4072
rect 354646 4032 367008 4060
rect 367002 4020 367008 4032
rect 367060 4020 367066 4072
rect 357434 3992 357440 4004
rect 340064 3964 357440 3992
rect 357434 3952 357440 3964
rect 357492 3952 357498 4004
rect 547138 3952 547144 4004
rect 547196 3992 547202 4004
rect 550266 3992 550272 4004
rect 547196 3964 550272 3992
rect 547196 3952 547202 3964
rect 550266 3952 550272 3964
rect 550324 3952 550330 4004
rect 563698 3952 563704 4004
rect 563756 3992 563762 4004
rect 568022 3992 568028 4004
rect 563756 3964 568028 3992
rect 563756 3952 563762 3964
rect 568022 3952 568028 3964
rect 568080 3952 568086 4004
rect 168466 3884 168472 3936
rect 168524 3924 168530 3936
rect 215570 3924 215576 3936
rect 168524 3896 215576 3924
rect 168524 3884 168530 3896
rect 215570 3884 215576 3896
rect 215628 3884 215634 3936
rect 252278 3884 252284 3936
rect 252336 3924 252342 3936
rect 372890 3924 372896 3936
rect 252336 3896 372896 3924
rect 252336 3884 252342 3896
rect 372890 3884 372896 3896
rect 372948 3884 372954 3936
rect 402514 3924 402520 3936
rect 383626 3896 402520 3924
rect 52546 3816 52552 3868
rect 52604 3856 52610 3868
rect 55858 3856 55864 3868
rect 52604 3828 55864 3856
rect 52604 3816 52610 3828
rect 55858 3816 55864 3828
rect 55916 3816 55922 3868
rect 62022 3816 62028 3868
rect 62080 3856 62086 3868
rect 66898 3856 66904 3868
rect 62080 3828 66904 3856
rect 62080 3816 62086 3828
rect 66898 3816 66904 3828
rect 66956 3816 66962 3868
rect 164878 3816 164884 3868
rect 164936 3856 164942 3868
rect 220354 3856 220360 3868
rect 164936 3828 220360 3856
rect 164936 3816 164942 3828
rect 220354 3816 220360 3828
rect 220412 3816 220418 3868
rect 252462 3816 252468 3868
rect 252520 3856 252526 3868
rect 376478 3856 376484 3868
rect 252520 3828 376484 3856
rect 252520 3816 252526 3828
rect 376478 3816 376484 3828
rect 376536 3816 376542 3868
rect 161290 3748 161296 3800
rect 161348 3788 161354 3800
rect 218698 3788 218704 3800
rect 161348 3760 218704 3788
rect 161348 3748 161354 3760
rect 218698 3748 218704 3760
rect 218756 3748 218762 3800
rect 249702 3748 249708 3800
rect 249760 3788 249766 3800
rect 259362 3788 259368 3800
rect 249760 3760 259368 3788
rect 249760 3748 249766 3760
rect 259362 3748 259368 3760
rect 259420 3748 259426 3800
rect 265342 3788 265348 3800
rect 259932 3760 265348 3788
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 46290 3720 46296 3732
rect 41932 3692 46296 3720
rect 41932 3680 41938 3692
rect 46290 3680 46296 3692
rect 46348 3680 46354 3732
rect 135254 3680 135260 3732
rect 135312 3720 135318 3732
rect 138658 3720 138664 3732
rect 135312 3692 138664 3720
rect 135312 3680 135318 3692
rect 138658 3680 138664 3692
rect 138716 3680 138722 3732
rect 155402 3680 155408 3732
rect 155460 3720 155466 3732
rect 218790 3720 218796 3732
rect 155460 3692 218796 3720
rect 155460 3680 155466 3692
rect 218790 3680 218796 3692
rect 218848 3680 218854 3732
rect 252370 3680 252376 3732
rect 252428 3720 252434 3732
rect 253474 3720 253480 3732
rect 252428 3692 253480 3720
rect 252428 3680 252434 3692
rect 253474 3680 253480 3692
rect 253532 3680 253538 3732
rect 253658 3680 253664 3732
rect 253716 3720 253722 3732
rect 259822 3720 259828 3732
rect 253716 3692 259828 3720
rect 253716 3680 253722 3692
rect 259822 3680 259828 3692
rect 259880 3680 259886 3732
rect 57238 3612 57244 3664
rect 57296 3652 57302 3664
rect 57296 3624 64874 3652
rect 57296 3612 57302 3624
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 10318 3584 10324 3596
rect 1728 3556 10324 3584
rect 1728 3544 1734 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 10428 3556 14596 3584
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 10428 3516 10456 3556
rect 7708 3488 10456 3516
rect 7708 3476 7714 3488
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14568 3516 14596 3556
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15838 3584 15844 3596
rect 14792 3556 15844 3584
rect 14792 3544 14798 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 46658 3544 46664 3596
rect 46716 3584 46722 3596
rect 46716 3556 50568 3584
rect 46716 3544 46722 3556
rect 21358 3516 21364 3528
rect 14568 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21818 3476 21824 3528
rect 21876 3516 21882 3528
rect 25498 3516 25504 3528
rect 21876 3488 25504 3516
rect 21876 3476 21882 3488
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 31294 3476 31300 3528
rect 31352 3516 31358 3528
rect 32398 3516 32404 3528
rect 31352 3488 32404 3516
rect 31352 3476 31358 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 39298 3516 39304 3528
rect 38436 3488 39304 3516
rect 38436 3476 38442 3488
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 50338 3516 50344 3528
rect 49016 3488 50344 3516
rect 49016 3476 49022 3488
rect 50338 3476 50344 3488
rect 50396 3476 50402 3528
rect 50540 3516 50568 3556
rect 53742 3544 53748 3596
rect 53800 3584 53806 3596
rect 54478 3584 54484 3596
rect 53800 3556 54484 3584
rect 53800 3544 53806 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 62758 3584 62764 3596
rect 59688 3556 62764 3584
rect 59688 3544 59694 3556
rect 62758 3544 62764 3556
rect 62816 3544 62822 3596
rect 64846 3584 64874 3624
rect 69106 3612 69112 3664
rect 69164 3652 69170 3664
rect 71038 3652 71044 3664
rect 69164 3624 71044 3652
rect 69164 3612 69170 3624
rect 71038 3612 71044 3624
rect 71096 3612 71102 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 97258 3652 97264 3664
rect 96304 3624 97264 3652
rect 96304 3612 96310 3624
rect 97258 3612 97264 3624
rect 97316 3612 97322 3664
rect 109310 3612 109316 3664
rect 109368 3652 109374 3664
rect 112438 3652 112444 3664
rect 109368 3624 112444 3652
rect 109368 3612 109374 3624
rect 112438 3612 112444 3624
rect 112496 3612 112502 3664
rect 121086 3612 121092 3664
rect 121144 3652 121150 3664
rect 122098 3652 122104 3664
rect 121144 3624 122104 3652
rect 121144 3612 121150 3624
rect 122098 3612 122104 3624
rect 122156 3612 122162 3664
rect 123478 3612 123484 3664
rect 123536 3652 123542 3664
rect 152458 3652 152464 3664
rect 123536 3624 152464 3652
rect 123536 3612 123542 3624
rect 152458 3612 152464 3624
rect 152516 3612 152522 3664
rect 160094 3612 160100 3664
rect 160152 3652 160158 3664
rect 235258 3652 235264 3664
rect 160152 3624 235264 3652
rect 160152 3612 160158 3624
rect 235258 3612 235264 3624
rect 235316 3612 235322 3664
rect 246850 3612 246856 3664
rect 246908 3652 246914 3664
rect 259932 3652 259960 3760
rect 265342 3748 265348 3760
rect 265400 3748 265406 3800
rect 278130 3748 278136 3800
rect 278188 3788 278194 3800
rect 383626 3788 383654 3896
rect 402514 3884 402520 3896
rect 402572 3884 402578 3936
rect 537478 3884 537484 3936
rect 537536 3924 537542 3936
rect 540790 3924 540796 3936
rect 537536 3896 540796 3924
rect 537536 3884 537542 3896
rect 540790 3884 540796 3896
rect 540848 3884 540854 3936
rect 390554 3856 390560 3868
rect 278188 3760 383654 3788
rect 385512 3828 390560 3856
rect 278188 3748 278194 3760
rect 260006 3680 260012 3732
rect 260064 3720 260070 3732
rect 385512 3720 385540 3828
rect 390554 3816 390560 3828
rect 390612 3816 390618 3868
rect 574738 3816 574744 3868
rect 574796 3856 574802 3868
rect 577406 3856 577412 3868
rect 574796 3828 577412 3856
rect 574796 3816 574802 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 260064 3692 385540 3720
rect 260064 3680 260070 3692
rect 385678 3680 385684 3732
rect 385736 3720 385742 3732
rect 388254 3720 388260 3732
rect 385736 3692 388260 3720
rect 385736 3680 385742 3692
rect 388254 3680 388260 3692
rect 388312 3680 388318 3732
rect 400858 3680 400864 3732
rect 400916 3720 400922 3732
rect 531314 3720 531320 3732
rect 400916 3692 531320 3720
rect 400916 3680 400922 3692
rect 531314 3680 531320 3692
rect 531372 3680 531378 3732
rect 246908 3624 259960 3652
rect 246908 3612 246914 3624
rect 260098 3612 260104 3664
rect 260156 3652 260162 3664
rect 261754 3652 261760 3664
rect 260156 3624 261760 3652
rect 260156 3612 260162 3624
rect 261754 3612 261760 3624
rect 261812 3612 261818 3664
rect 269758 3612 269764 3664
rect 269816 3652 269822 3664
rect 274818 3652 274824 3664
rect 269816 3624 274824 3652
rect 269816 3612 269822 3624
rect 274818 3612 274824 3624
rect 274876 3612 274882 3664
rect 285398 3652 285404 3664
rect 274928 3624 285404 3652
rect 123386 3584 123392 3596
rect 64846 3556 123392 3584
rect 123386 3544 123392 3556
rect 123444 3544 123450 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 210418 3584 210424 3596
rect 129424 3556 210424 3584
rect 129424 3544 129430 3556
rect 210418 3544 210424 3556
rect 210476 3544 210482 3596
rect 213178 3544 213184 3596
rect 213236 3544 213242 3596
rect 226426 3544 226432 3596
rect 226484 3584 226490 3596
rect 233970 3584 233976 3596
rect 226484 3556 233976 3584
rect 226484 3544 226490 3556
rect 233970 3544 233976 3556
rect 234028 3544 234034 3596
rect 242986 3544 242992 3596
rect 243044 3584 243050 3596
rect 243044 3556 244228 3584
rect 243044 3544 243050 3556
rect 175918 3516 175924 3528
rect 50540 3488 175924 3516
rect 175918 3476 175924 3488
rect 175976 3476 175982 3528
rect 186130 3476 186136 3528
rect 186188 3516 186194 3528
rect 213196 3516 213224 3544
rect 186188 3488 213224 3516
rect 186188 3476 186194 3488
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 238018 3516 238024 3528
rect 215720 3488 238024 3516
rect 215720 3476 215726 3488
rect 238018 3476 238024 3488
rect 238076 3476 238082 3528
rect 241330 3476 241336 3528
rect 241388 3516 241394 3528
rect 244090 3516 244096 3528
rect 241388 3488 244096 3516
rect 241388 3476 241394 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 244200 3516 244228 3556
rect 246942 3544 246948 3596
rect 247000 3584 247006 3596
rect 270862 3584 270868 3596
rect 247000 3556 270868 3584
rect 247000 3544 247006 3556
rect 270862 3544 270868 3556
rect 270920 3544 270926 3596
rect 271138 3544 271144 3596
rect 271196 3584 271202 3596
rect 274928 3584 274956 3624
rect 285398 3612 285404 3624
rect 285456 3612 285462 3664
rect 291838 3612 291844 3664
rect 291896 3652 291902 3664
rect 306742 3652 306748 3664
rect 291896 3624 306748 3652
rect 291896 3612 291902 3624
rect 306742 3612 306748 3624
rect 306800 3612 306806 3664
rect 313918 3612 313924 3664
rect 313976 3652 313982 3664
rect 317322 3652 317328 3664
rect 313976 3624 317328 3652
rect 313976 3612 313982 3624
rect 317322 3612 317328 3624
rect 317380 3612 317386 3664
rect 330478 3612 330484 3664
rect 330536 3652 330542 3664
rect 485222 3652 485228 3664
rect 330536 3624 485228 3652
rect 330536 3612 330542 3624
rect 485222 3612 485228 3624
rect 485280 3612 485286 3664
rect 493318 3612 493324 3664
rect 493376 3652 493382 3664
rect 552658 3652 552664 3664
rect 493376 3624 552664 3652
rect 493376 3612 493382 3624
rect 552658 3612 552664 3624
rect 552716 3612 552722 3664
rect 271196 3556 274956 3584
rect 271196 3544 271202 3556
rect 275278 3544 275284 3596
rect 275336 3584 275342 3596
rect 275336 3556 277394 3584
rect 275336 3544 275342 3556
rect 267734 3516 267740 3528
rect 244200 3488 267740 3516
rect 267734 3476 267740 3488
rect 267792 3476 267798 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 272426 3516 272432 3528
rect 271288 3488 272432 3516
rect 271288 3476 271294 3488
rect 272426 3476 272432 3488
rect 272484 3476 272490 3528
rect 273898 3476 273904 3528
rect 273956 3516 273962 3528
rect 276014 3516 276020 3528
rect 273956 3488 276020 3516
rect 273956 3476 273962 3488
rect 276014 3476 276020 3488
rect 276072 3476 276078 3528
rect 277366 3516 277394 3556
rect 278038 3544 278044 3596
rect 278096 3584 278102 3596
rect 296070 3584 296076 3596
rect 278096 3556 296076 3584
rect 278096 3544 278102 3556
rect 296070 3544 296076 3556
rect 296128 3544 296134 3596
rect 298738 3544 298744 3596
rect 298796 3584 298802 3596
rect 298796 3556 311112 3584
rect 298796 3544 298802 3556
rect 277366 3488 289032 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 217318 3448 217324 3460
rect 6512 3420 217324 3448
rect 6512 3408 6518 3420
rect 217318 3408 217324 3420
rect 217376 3408 217382 3460
rect 226334 3408 226340 3460
rect 226392 3448 226398 3460
rect 227530 3448 227536 3460
rect 226392 3420 227536 3448
rect 226392 3408 226398 3420
rect 227530 3408 227536 3420
rect 227588 3408 227594 3460
rect 229830 3408 229836 3460
rect 229888 3448 229894 3460
rect 240778 3448 240784 3460
rect 229888 3420 240784 3448
rect 229888 3408 229894 3420
rect 240778 3408 240784 3420
rect 240836 3408 240842 3460
rect 241422 3408 241428 3460
rect 241480 3448 241486 3460
rect 242894 3448 242900 3460
rect 241480 3420 242900 3448
rect 241480 3408 241486 3420
rect 242894 3408 242900 3420
rect 242952 3408 242958 3460
rect 245562 3408 245568 3460
rect 245620 3448 245626 3460
rect 287790 3448 287796 3460
rect 245620 3420 287796 3448
rect 245620 3408 245626 3420
rect 287790 3408 287796 3420
rect 287848 3408 287854 3460
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 90358 3380 90364 3392
rect 89220 3352 90364 3380
rect 89220 3340 89226 3352
rect 90358 3340 90364 3352
rect 90416 3340 90422 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 114002 3340 114008 3392
rect 114060 3380 114066 3392
rect 115198 3380 115204 3392
rect 114060 3352 115204 3380
rect 114060 3340 114066 3352
rect 115198 3340 115204 3352
rect 115256 3340 115262 3392
rect 136450 3340 136456 3392
rect 136508 3380 136514 3392
rect 137278 3380 137284 3392
rect 136508 3352 137284 3380
rect 136508 3340 136514 3352
rect 137278 3340 137284 3352
rect 137336 3340 137342 3392
rect 153010 3340 153016 3392
rect 153068 3380 153074 3392
rect 155218 3380 155224 3392
rect 153068 3352 155224 3380
rect 153068 3340 153074 3352
rect 155218 3340 155224 3352
rect 155276 3340 155282 3392
rect 168374 3340 168380 3392
rect 168432 3380 168438 3392
rect 169570 3380 169576 3392
rect 168432 3352 169576 3380
rect 168432 3340 168438 3352
rect 169570 3340 169576 3352
rect 169628 3340 169634 3392
rect 193214 3340 193220 3392
rect 193272 3380 193278 3392
rect 194410 3380 194416 3392
rect 193272 3352 194416 3380
rect 193272 3340 193278 3352
rect 194410 3340 194416 3352
rect 194468 3340 194474 3392
rect 249518 3340 249524 3392
rect 249576 3380 249582 3392
rect 251174 3380 251180 3392
rect 249576 3352 251180 3380
rect 249576 3340 249582 3352
rect 251174 3340 251180 3352
rect 251232 3340 251238 3392
rect 253198 3340 253204 3392
rect 253256 3380 253262 3392
rect 254670 3380 254676 3392
rect 253256 3352 254676 3380
rect 253256 3340 253262 3352
rect 254670 3340 254676 3352
rect 254728 3340 254734 3392
rect 259362 3340 259368 3392
rect 259420 3380 259426 3392
rect 264146 3380 264152 3392
rect 259420 3352 264152 3380
rect 259420 3340 259426 3352
rect 264146 3340 264152 3352
rect 264204 3340 264210 3392
rect 289004 3380 289032 3488
rect 289078 3476 289084 3528
rect 289136 3516 289142 3528
rect 290182 3516 290188 3528
rect 289136 3488 290188 3516
rect 289136 3476 289142 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 300118 3476 300124 3528
rect 300176 3516 300182 3528
rect 301958 3516 301964 3528
rect 300176 3488 301964 3516
rect 300176 3476 300182 3488
rect 301958 3476 301964 3488
rect 302016 3476 302022 3528
rect 307018 3476 307024 3528
rect 307076 3516 307082 3528
rect 309042 3516 309048 3528
rect 307076 3488 309048 3516
rect 307076 3476 307082 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 311084 3516 311112 3556
rect 311158 3544 311164 3596
rect 311216 3584 311222 3596
rect 312630 3584 312636 3596
rect 311216 3556 312636 3584
rect 311216 3544 311222 3556
rect 312630 3544 312636 3556
rect 312688 3544 312694 3596
rect 327718 3544 327724 3596
rect 327776 3544 327782 3596
rect 329098 3544 329104 3596
rect 329156 3584 329162 3596
rect 495894 3584 495900 3596
rect 329156 3556 495900 3584
rect 329156 3544 329162 3556
rect 495894 3544 495900 3556
rect 495952 3544 495958 3596
rect 498194 3544 498200 3596
rect 498252 3584 498258 3596
rect 499022 3584 499028 3596
rect 498252 3556 499028 3584
rect 498252 3544 498258 3556
rect 499022 3544 499028 3556
rect 499080 3544 499086 3596
rect 500218 3544 500224 3596
rect 500276 3584 500282 3596
rect 502886 3584 502892 3596
rect 500276 3556 502892 3584
rect 500276 3544 500282 3556
rect 502886 3544 502892 3556
rect 502944 3544 502950 3596
rect 502978 3544 502984 3596
rect 503036 3584 503042 3596
rect 505370 3584 505376 3596
rect 503036 3556 505376 3584
rect 503036 3544 503042 3556
rect 505370 3544 505376 3556
rect 505428 3544 505434 3596
rect 554038 3544 554044 3596
rect 554096 3584 554102 3596
rect 556154 3584 556160 3596
rect 554096 3556 556160 3584
rect 554096 3544 554102 3556
rect 556154 3544 556160 3556
rect 556212 3544 556218 3596
rect 313826 3516 313832 3528
rect 311084 3488 313832 3516
rect 313826 3476 313832 3488
rect 313884 3476 313890 3528
rect 318058 3476 318064 3528
rect 318116 3516 318122 3528
rect 319714 3516 319720 3528
rect 318116 3488 319720 3516
rect 318116 3476 318122 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 320818 3476 320824 3528
rect 320876 3516 320882 3528
rect 325602 3516 325608 3528
rect 320876 3488 325608 3516
rect 320876 3476 320882 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 327736 3516 327764 3544
rect 517146 3516 517152 3528
rect 327736 3488 517152 3516
rect 517146 3476 517152 3488
rect 517204 3476 517210 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 526438 3476 526444 3528
rect 526496 3516 526502 3528
rect 527818 3516 527824 3528
rect 526496 3488 527824 3516
rect 526496 3476 526502 3488
rect 527818 3476 527824 3488
rect 527876 3476 527882 3528
rect 536190 3476 536196 3528
rect 536248 3516 536254 3528
rect 537202 3516 537208 3528
rect 536248 3488 537208 3516
rect 536248 3476 536254 3488
rect 537202 3476 537208 3488
rect 537260 3476 537266 3528
rect 540238 3476 540244 3528
rect 540296 3516 540302 3528
rect 547874 3516 547880 3528
rect 540296 3488 547880 3516
rect 540296 3476 540302 3488
rect 547874 3476 547880 3488
rect 547932 3476 547938 3528
rect 555510 3476 555516 3528
rect 555568 3516 555574 3528
rect 557350 3516 557356 3528
rect 555568 3488 557356 3516
rect 555568 3476 555574 3488
rect 557350 3476 557356 3488
rect 557408 3476 557414 3528
rect 559558 3476 559564 3528
rect 559616 3516 559622 3528
rect 560846 3516 560852 3528
rect 559616 3488 560852 3516
rect 559616 3476 559622 3488
rect 560846 3476 560852 3488
rect 560904 3476 560910 3528
rect 289170 3408 289176 3460
rect 289228 3448 289234 3460
rect 291378 3448 291384 3460
rect 289228 3420 291384 3448
rect 289228 3408 289234 3420
rect 291378 3408 291384 3420
rect 291436 3408 291442 3460
rect 295978 3408 295984 3460
rect 296036 3448 296042 3460
rect 296036 3420 296714 3448
rect 296036 3408 296042 3420
rect 292574 3380 292580 3392
rect 289004 3352 292580 3380
rect 292574 3340 292580 3352
rect 292632 3340 292638 3392
rect 296686 3380 296714 3420
rect 299566 3408 299572 3460
rect 299624 3448 299630 3460
rect 300762 3448 300768 3460
rect 299624 3420 300768 3448
rect 299624 3408 299630 3420
rect 300762 3408 300768 3420
rect 300820 3408 300826 3460
rect 305638 3408 305644 3460
rect 305696 3448 305702 3460
rect 329190 3448 329196 3460
rect 305696 3420 329196 3448
rect 305696 3408 305702 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 329282 3408 329288 3460
rect 329340 3448 329346 3460
rect 520734 3448 520740 3460
rect 329340 3420 520740 3448
rect 329340 3408 329346 3420
rect 520734 3408 520740 3420
rect 520792 3408 520798 3460
rect 529198 3408 529204 3460
rect 529256 3448 529262 3460
rect 554958 3448 554964 3460
rect 529256 3420 554964 3448
rect 529256 3408 529262 3420
rect 554958 3408 554964 3420
rect 555016 3408 555022 3460
rect 555418 3408 555424 3460
rect 555476 3448 555482 3460
rect 562042 3448 562048 3460
rect 555476 3420 562048 3448
rect 555476 3408 555482 3420
rect 562042 3408 562048 3420
rect 562100 3408 562106 3460
rect 565078 3408 565084 3460
rect 565136 3448 565142 3460
rect 572714 3448 572720 3460
rect 565136 3420 572720 3448
rect 565136 3408 565142 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 299658 3380 299664 3392
rect 296686 3352 299664 3380
rect 299658 3340 299664 3352
rect 299716 3340 299722 3392
rect 324958 3340 324964 3392
rect 325016 3380 325022 3392
rect 326798 3380 326804 3392
rect 325016 3352 326804 3380
rect 325016 3340 325022 3352
rect 326798 3340 326804 3352
rect 326856 3340 326862 3392
rect 332042 3340 332048 3392
rect 332100 3380 332106 3392
rect 342162 3380 342168 3392
rect 332100 3352 342168 3380
rect 332100 3340 332106 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357526 3340 357532 3392
rect 357584 3380 357590 3392
rect 358722 3380 358728 3392
rect 357584 3352 358728 3380
rect 357584 3340 357590 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 376018 3340 376024 3392
rect 376076 3380 376082 3392
rect 377674 3380 377680 3392
rect 376076 3352 377680 3380
rect 376076 3340 376082 3352
rect 377674 3340 377680 3352
rect 377732 3340 377738 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 422938 3340 422944 3392
rect 422996 3380 423002 3392
rect 424962 3380 424968 3392
rect 422996 3352 424968 3380
rect 422996 3340 423002 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 436738 3340 436744 3392
rect 436796 3380 436802 3392
rect 437934 3380 437940 3392
rect 436796 3352 437940 3380
rect 436796 3340 436802 3352
rect 437934 3340 437940 3352
rect 437992 3340 437998 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 443638 3340 443644 3392
rect 443696 3380 443702 3392
rect 445018 3380 445024 3392
rect 443696 3352 445024 3380
rect 443696 3340 443702 3352
rect 445018 3340 445024 3352
rect 445076 3340 445082 3392
rect 456886 3340 456892 3392
rect 456944 3380 456950 3392
rect 458082 3380 458088 3392
rect 456944 3352 458088 3380
rect 456944 3340 456950 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 461670 3340 461676 3392
rect 461728 3380 461734 3392
rect 469858 3380 469864 3392
rect 461728 3352 469864 3380
rect 461728 3340 461734 3352
rect 469858 3340 469864 3352
rect 469916 3340 469922 3392
rect 77386 3272 77392 3324
rect 77444 3312 77450 3324
rect 79318 3312 79324 3324
rect 77444 3284 79324 3312
rect 77444 3272 77450 3284
rect 79318 3272 79324 3284
rect 79376 3272 79382 3324
rect 335906 3272 335912 3324
rect 335964 3312 335970 3324
rect 343358 3312 343364 3324
rect 335964 3284 343364 3312
rect 335964 3272 335970 3284
rect 343358 3272 343364 3284
rect 343416 3272 343422 3324
rect 417510 3272 417516 3324
rect 417568 3312 417574 3324
rect 420178 3312 420184 3324
rect 417568 3284 420184 3312
rect 417568 3272 417574 3284
rect 420178 3272 420184 3284
rect 420236 3272 420242 3324
rect 421558 3272 421564 3324
rect 421616 3312 421622 3324
rect 423766 3312 423772 3324
rect 421616 3284 423772 3312
rect 421616 3272 421622 3284
rect 423766 3272 423772 3284
rect 423824 3272 423830 3324
rect 454678 3272 454684 3324
rect 454736 3312 454742 3324
rect 455690 3312 455696 3324
rect 454736 3284 455696 3312
rect 454736 3272 454742 3284
rect 455690 3272 455696 3284
rect 455748 3272 455754 3324
rect 562318 3272 562324 3324
rect 562376 3312 562382 3324
rect 565630 3312 565636 3324
rect 562376 3284 565636 3312
rect 562376 3272 562382 3284
rect 565630 3272 565636 3284
rect 565688 3272 565694 3324
rect 27706 3204 27712 3256
rect 27764 3244 27770 3256
rect 31018 3244 31024 3256
rect 27764 3216 31024 3244
rect 27764 3204 27770 3216
rect 31018 3204 31024 3216
rect 31076 3204 31082 3256
rect 243630 3204 243636 3256
rect 243688 3244 243694 3256
rect 248782 3244 248788 3256
rect 243688 3216 248788 3244
rect 243688 3204 243694 3216
rect 248782 3204 248788 3216
rect 248840 3204 248846 3256
rect 519630 3204 519636 3256
rect 519688 3244 519694 3256
rect 525426 3244 525432 3256
rect 519688 3216 525432 3244
rect 519688 3204 519694 3216
rect 525426 3204 525432 3216
rect 525484 3204 525490 3256
rect 64322 3136 64328 3188
rect 64380 3176 64386 3188
rect 65518 3176 65524 3188
rect 64380 3148 65524 3176
rect 64380 3136 64386 3148
rect 65518 3136 65524 3148
rect 65576 3136 65582 3188
rect 124674 3136 124680 3188
rect 124732 3176 124738 3188
rect 126238 3176 126244 3188
rect 124732 3148 126244 3176
rect 124732 3136 124738 3148
rect 126238 3136 126244 3148
rect 126296 3136 126302 3188
rect 309870 3136 309876 3188
rect 309928 3176 309934 3188
rect 315022 3176 315028 3188
rect 309928 3148 315028 3176
rect 309928 3136 309934 3148
rect 315022 3136 315028 3148
rect 315080 3136 315086 3188
rect 512638 3136 512644 3188
rect 512696 3176 512702 3188
rect 515950 3176 515956 3188
rect 512696 3148 515956 3176
rect 512696 3136 512702 3148
rect 515950 3136 515956 3148
rect 516008 3136 516014 3188
rect 223942 3068 223948 3120
rect 224000 3108 224006 3120
rect 226978 3108 226984 3120
rect 224000 3080 226984 3108
rect 224000 3068 224006 3080
rect 226978 3068 226984 3080
rect 227036 3068 227042 3120
rect 273162 3068 273168 3120
rect 273220 3108 273226 3120
rect 277118 3108 277124 3120
rect 273220 3080 277124 3108
rect 273220 3068 273226 3080
rect 277118 3068 277124 3080
rect 277176 3068 277182 3120
rect 406378 3068 406384 3120
rect 406436 3108 406442 3120
rect 409598 3108 409604 3120
rect 406436 3080 409604 3108
rect 406436 3068 406442 3080
rect 409598 3068 409604 3080
rect 409656 3068 409662 3120
rect 542998 3068 543004 3120
rect 543056 3108 543062 3120
rect 545482 3108 545488 3120
rect 543056 3080 545488 3108
rect 543056 3068 543062 3080
rect 545482 3068 545488 3080
rect 545540 3068 545546 3120
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 19978 3040 19984 3052
rect 17092 3012 19984 3040
rect 17092 3000 17098 3012
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 154206 3000 154212 3052
rect 154264 3040 154270 3052
rect 155310 3040 155316 3052
rect 154264 3012 155316 3040
rect 154264 3000 154270 3012
rect 155310 3000 155316 3012
rect 155368 3000 155374 3052
rect 351270 3000 351276 3052
rect 351328 3040 351334 3052
rect 352834 3040 352840 3052
rect 351328 3012 352840 3040
rect 351328 3000 351334 3012
rect 352834 3000 352840 3012
rect 352892 3000 352898 3052
rect 447778 3000 447784 3052
rect 447836 3040 447842 3052
rect 448606 3040 448612 3052
rect 447836 3012 448612 3040
rect 447836 3000 447842 3012
rect 448606 3000 448612 3012
rect 448664 3000 448670 3052
rect 472618 3000 472624 3052
rect 472676 3040 472682 3052
rect 473446 3040 473452 3052
rect 472676 3012 473452 3040
rect 472676 3000 472682 3012
rect 473446 3000 473452 3012
rect 473504 3000 473510 3052
rect 530578 3000 530584 3052
rect 530636 3040 530642 3052
rect 532510 3040 532516 3052
rect 530636 3012 532516 3040
rect 530636 3000 530642 3012
rect 532510 3000 532516 3012
rect 532568 3000 532574 3052
rect 189718 2932 189724 2984
rect 189776 2972 189782 2984
rect 191098 2972 191104 2984
rect 189776 2944 191104 2972
rect 189776 2932 189782 2944
rect 191098 2932 191104 2944
rect 191156 2932 191162 2984
rect 358078 2864 358084 2916
rect 358136 2904 358142 2916
rect 361114 2904 361120 2916
rect 358136 2876 361120 2904
rect 358136 2864 358142 2876
rect 361114 2864 361120 2876
rect 361172 2864 361178 2916
rect 511350 2864 511356 2916
rect 511408 2904 511414 2916
rect 513558 2904 513564 2916
rect 511408 2876 513564 2904
rect 511408 2864 511414 2876
rect 513558 2864 513564 2876
rect 513616 2864 513622 2916
rect 398834 2592 398840 2644
rect 398892 2632 398898 2644
rect 400122 2632 400128 2644
rect 398892 2604 400128 2632
rect 398892 2592 398898 2604
rect 400122 2592 400128 2604
rect 400180 2592 400186 2644
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 283840 700272 283892 700324
rect 305000 700272 305052 700324
rect 340144 700272 340196 700324
rect 348792 700272 348844 700324
rect 403624 700272 403676 700324
rect 413652 700272 413704 700324
rect 414664 700272 414716 700324
rect 478512 700272 478564 700324
rect 154120 700068 154172 700120
rect 155224 700068 155276 700120
rect 8116 699660 8168 699712
rect 10324 699660 10376 699712
rect 24308 699660 24360 699712
rect 26884 699660 26936 699712
rect 89168 699660 89220 699712
rect 90364 699660 90416 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 526444 699660 526496 699712
rect 527180 699660 527232 699712
rect 218980 698912 219032 698964
rect 306380 698912 306432 698964
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 299664 696940 299716 696992
rect 580172 696940 580224 696992
rect 300124 683204 300176 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 310520 683136 310572 683188
rect 3516 670692 3568 670744
rect 310612 670692 310664 670744
rect 330484 670692 330536 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 310704 656888 310756 656940
rect 323584 643084 323636 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 289084 632068 289136 632120
rect 298744 630640 298796 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 302884 618264 302936 618316
rect 363604 616836 363656 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 291844 605820 291896 605872
rect 324964 590656 325016 590708
rect 579804 590656 579856 590708
rect 334624 576852 334676 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 313280 565836 313332 565888
rect 319444 563048 319496 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 46204 553392 46256 553444
rect 320824 536800 320876 536852
rect 580172 536800 580224 536852
rect 2780 527144 2832 527196
rect 4804 527144 4856 527196
rect 329104 524424 329156 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 250444 514768 250496 514820
rect 318064 510620 318116 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 14464 500964 14516 501016
rect 322204 484372 322256 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 7564 474716 7616 474768
rect 399484 470568 399536 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 314752 462340 314804 462392
rect 3148 448536 3200 448588
rect 15844 448536 15896 448588
rect 295984 447788 296036 447840
rect 399484 447788 399536 447840
rect 294604 430584 294656 430636
rect 579896 430584 579948 430636
rect 3516 422288 3568 422340
rect 151084 422288 151136 422340
rect 294696 418140 294748 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 309600 409844 309652 409896
rect 26884 407736 26936 407788
rect 309140 407736 309192 407788
rect 250444 406376 250496 406428
rect 314844 406376 314896 406428
rect 294788 404336 294840 404388
rect 580172 404336 580224 404388
rect 309600 403588 309652 403640
rect 316040 403588 316092 403640
rect 304264 402228 304316 402280
rect 340144 402228 340196 402280
rect 302976 400868 303028 400920
rect 414664 400868 414716 400920
rect 298836 399440 298888 399492
rect 334624 399440 334676 399492
rect 304356 398080 304408 398132
rect 403624 398080 403676 398132
rect 3516 397468 3568 397520
rect 305644 397468 305696 397520
rect 297364 396720 297416 396772
rect 329104 396720 329156 396772
rect 302884 395360 302936 395412
rect 311900 395360 311952 395412
rect 14464 395292 14516 395344
rect 313372 395292 313424 395344
rect 201500 394000 201552 394052
rect 306472 394000 306524 394052
rect 301504 393932 301556 393984
rect 542360 393932 542412 393984
rect 304448 392640 304500 392692
rect 331220 392640 331272 392692
rect 155224 392572 155276 392624
rect 307760 392572 307812 392624
rect 15844 391212 15896 391264
rect 255320 391212 255372 391264
rect 302884 391212 302936 391264
rect 396724 391212 396776 391264
rect 255320 390532 255372 390584
rect 314936 390532 314988 390584
rect 303252 389784 303304 389836
rect 462320 389784 462372 389836
rect 298928 388492 298980 388544
rect 323584 388492 323636 388544
rect 10324 388424 10376 388476
rect 309232 388424 309284 388476
rect 296076 387132 296128 387184
rect 322204 387132 322256 387184
rect 136640 387064 136692 387116
rect 307852 387064 307904 387116
rect 296720 385636 296772 385688
rect 324964 385636 325016 385688
rect 151084 384344 151136 384396
rect 316132 384344 316184 384396
rect 301044 384276 301096 384328
rect 526444 384276 526496 384328
rect 245660 382984 245712 383036
rect 266360 382984 266412 383036
rect 305552 383052 305604 383104
rect 303344 382984 303396 383036
rect 429200 382984 429252 383036
rect 71780 382916 71832 382968
rect 307944 382916 307996 382968
rect 301780 381488 301832 381540
rect 494060 381488 494112 381540
rect 291844 380196 291896 380248
rect 312084 380196 312136 380248
rect 299756 380128 299808 380180
rect 330484 380128 330536 380180
rect 292580 378156 292632 378208
rect 580172 378156 580224 378208
rect 297088 377476 297140 377528
rect 320824 377476 320876 377528
rect 298928 377408 298980 377460
rect 363604 377408 363656 377460
rect 262128 376728 262180 376780
rect 322388 376728 322440 376780
rect 296628 376116 296680 376168
rect 318064 376116 318116 376168
rect 303160 376048 303212 376100
rect 558920 376048 558972 376100
rect 3424 375980 3476 376032
rect 312820 375980 312872 376032
rect 275100 375844 275152 375896
rect 306380 375844 306432 375896
rect 236644 375776 236696 375828
rect 294696 375776 294748 375828
rect 294880 375776 294932 375828
rect 249800 375708 249852 375760
rect 309140 375708 309192 375760
rect 239404 375640 239456 375692
rect 298836 375640 298888 375692
rect 244280 375572 244332 375624
rect 304264 375572 304316 375624
rect 304724 375572 304776 375624
rect 238760 375504 238812 375556
rect 298744 375504 298796 375556
rect 240140 375436 240192 375488
rect 300308 375436 300360 375488
rect 236000 375368 236052 375420
rect 297364 375368 297416 375420
rect 298744 375368 298796 375420
rect 299388 375368 299440 375420
rect 306380 375368 306432 375420
rect 306932 375368 306984 375420
rect 309140 375368 309192 375420
rect 310244 375368 310296 375420
rect 262496 374892 262548 374944
rect 323124 374892 323176 374944
rect 278596 374824 278648 374876
rect 296076 374824 296128 374876
rect 297824 374824 297876 374876
rect 319444 374824 319496 374876
rect 277952 374756 278004 374808
rect 304540 374756 304592 374808
rect 275744 374688 275796 374740
rect 304356 374688 304408 374740
rect 278504 374620 278556 374672
rect 295892 374620 295944 374672
rect 253204 374552 253256 374604
rect 294788 374552 294840 374604
rect 295524 374552 295576 374604
rect 580264 374620 580316 374672
rect 275192 374484 275244 374536
rect 319076 374484 319128 374536
rect 255964 374416 256016 374468
rect 299756 374416 299808 374468
rect 257344 374348 257396 374400
rect 300768 374348 300820 374400
rect 303160 374348 303212 374400
rect 313280 374348 313332 374400
rect 313464 374348 313516 374400
rect 259644 374280 259696 374332
rect 319812 374280 319864 374332
rect 264888 374212 264940 374264
rect 325332 374212 325384 374264
rect 234712 374144 234764 374196
rect 294604 374144 294656 374196
rect 260104 374076 260156 374128
rect 320180 374076 320232 374128
rect 281080 374008 281132 374060
rect 297824 374008 297876 374060
rect 295800 373600 295852 373652
rect 296076 373600 296128 373652
rect 294328 373532 294380 373584
rect 294788 373532 294840 373584
rect 230480 373328 230532 373380
rect 291568 373328 291620 373380
rect 304448 373328 304500 373380
rect 364340 373328 364392 373380
rect 234620 373260 234672 373312
rect 248420 373260 248472 373312
rect 262404 373192 262456 373244
rect 313740 373192 313792 373244
rect 258816 373124 258868 373176
rect 317328 373124 317380 373176
rect 257436 373056 257488 373108
rect 317236 373056 317288 373108
rect 229100 372988 229152 373040
rect 288992 372988 289044 373040
rect 577596 372988 577648 373040
rect 258724 372920 258776 372972
rect 318800 372920 318852 372972
rect 262312 372852 262364 372904
rect 322940 372852 322992 372904
rect 259552 372784 259604 372836
rect 320548 372784 320600 372836
rect 261024 372716 261076 372768
rect 321652 372716 321704 372768
rect 275928 372648 275980 372700
rect 323492 372648 323544 372700
rect 3424 372580 3476 372632
rect 256700 372580 256752 372632
rect 257436 372580 257488 372632
rect 281172 372580 281224 372632
rect 295524 372580 295576 372632
rect 307760 372512 307812 372564
rect 308036 372512 308088 372564
rect 245752 372172 245804 372224
rect 305000 372172 305052 372224
rect 305828 372172 305880 372224
rect 245016 372104 245068 372156
rect 292212 372104 292264 372156
rect 363604 372104 363656 372156
rect 243544 372036 243596 372088
rect 288256 372036 288308 372088
rect 289268 372036 289320 372088
rect 577504 372036 577556 372088
rect 279516 371968 279568 372020
rect 290556 371968 290608 372020
rect 313740 371968 313792 372020
rect 322020 371968 322072 372020
rect 280804 371900 280856 371952
rect 314752 371900 314804 371952
rect 315764 371900 315816 371952
rect 280896 371832 280948 371884
rect 316040 371832 316092 371884
rect 316868 371832 316920 371884
rect 280436 371764 280488 371816
rect 317972 371764 318024 371816
rect 279424 371696 279476 371748
rect 321284 371696 321336 371748
rect 280988 371628 281040 371680
rect 313464 371628 313516 371680
rect 280252 371560 280304 371612
rect 324596 371560 324648 371612
rect 247684 371492 247736 371544
rect 293684 371492 293736 371544
rect 293960 371492 294012 371544
rect 336004 371492 336056 371544
rect 250444 371424 250496 371476
rect 308036 371424 308088 371476
rect 308864 371424 308916 371476
rect 316132 371424 316184 371476
rect 317328 371424 317380 371476
rect 318340 371424 318392 371476
rect 290556 371356 290608 371408
rect 299480 371356 299532 371408
rect 282000 371288 282052 371340
rect 291844 371288 291896 371340
rect 299296 371288 299348 371340
rect 314844 371356 314896 371408
rect 242164 371220 242216 371272
rect 289268 371220 289320 371272
rect 314568 371220 314620 371272
rect 319444 371220 319496 371272
rect 319536 371220 319588 371272
rect 323860 371220 323912 371272
rect 241520 370744 241572 370796
rect 302240 370744 302292 370796
rect 303252 370744 303304 370796
rect 260196 370676 260248 370728
rect 314568 370676 314620 370728
rect 229192 370608 229244 370660
rect 290004 370608 290056 370660
rect 293684 370608 293736 370660
rect 236092 370540 236144 370592
rect 297088 370540 297140 370592
rect 231952 370472 232004 370524
rect 292948 370472 293000 370524
rect 293776 370472 293828 370524
rect 302332 370608 302384 370660
rect 580356 370608 580408 370660
rect 299480 370540 299532 370592
rect 580540 370540 580592 370592
rect 580172 370472 580224 370524
rect 244924 370404 244976 370456
rect 296628 370404 296680 370456
rect 231860 370336 231912 370388
rect 292672 370336 292724 370388
rect 329104 370336 329156 370388
rect 242900 370268 242952 370320
rect 302884 370268 302936 370320
rect 245844 370200 245896 370252
rect 306564 370200 306616 370252
rect 247040 370132 247092 370184
rect 307668 370132 307720 370184
rect 277860 370064 277912 370116
rect 293178 370064 293230 370116
rect 329196 370064 329248 370116
rect 282276 369996 282328 370048
rect 317604 369996 317656 370048
rect 281356 369928 281408 369980
rect 281448 369860 281500 369912
rect 288532 369860 288584 369912
rect 291568 369928 291620 369980
rect 330484 369928 330536 369980
rect 290740 369860 290792 369912
rect 290464 369656 290516 369708
rect 345664 369860 345716 369912
rect 291936 369588 291988 369640
rect 292212 369588 292264 369640
rect 282368 369384 282420 369436
rect 284116 369384 284168 369436
rect 282184 369316 282236 369368
rect 290004 369384 290056 369436
rect 308864 369452 308916 369504
rect 255412 369248 255464 369300
rect 245936 369180 245988 369232
rect 248420 369180 248472 369232
rect 282460 369180 282512 369232
rect 229284 369112 229336 369164
rect 282184 369112 282236 369164
rect 292304 369384 292356 369436
rect 293316 369384 293368 369436
rect 306288 369384 306340 369436
rect 326252 369384 326304 369436
rect 329012 369384 329064 369436
rect 233240 368500 233292 368552
rect 282460 368772 282512 368824
rect 264244 366324 264296 366376
rect 280252 366324 280304 366376
rect 258356 364352 258408 364404
rect 280436 364352 280488 364404
rect 223764 360204 223816 360256
rect 280712 360204 280764 360256
rect 226340 358776 226392 358828
rect 280068 358776 280120 358828
rect 280712 358776 280764 358828
rect 3424 358028 3476 358080
rect 258356 358028 258408 358080
rect 252560 356668 252612 356720
rect 280988 356668 281040 356720
rect 329196 353200 329248 353252
rect 579620 353200 579672 353252
rect 3332 345040 3384 345092
rect 256792 345040 256844 345092
rect 230572 327700 230624 327752
rect 279516 327700 279568 327752
rect 261484 326340 261536 326392
rect 279424 326340 279476 326392
rect 329104 325592 329156 325644
rect 580172 325592 580224 325644
rect 256884 324912 256936 324964
rect 280896 324912 280948 324964
rect 255504 323552 255556 323604
rect 280804 323552 280856 323604
rect 225052 322192 225104 322244
rect 279976 322192 280028 322244
rect 280804 322192 280856 322244
rect 281908 320968 281960 321020
rect 282276 320696 282328 320748
rect 283702 320696 283754 320748
rect 282184 320628 282236 320680
rect 211068 320560 211120 320612
rect 285818 320560 285870 320612
rect 272616 320492 272668 320544
rect 281908 320492 281960 320544
rect 302930 320628 302982 320680
rect 248512 320424 248564 320476
rect 249984 320356 250036 320408
rect 282184 320356 282236 320408
rect 219164 320288 219216 320340
rect 292442 320288 292494 320340
rect 275652 320220 275704 320272
rect 219348 320152 219400 320204
rect 280712 320084 280764 320136
rect 224868 319676 224920 319728
rect 284622 320016 284674 320068
rect 287014 320016 287066 320068
rect 282000 319880 282052 319932
rect 283334 319880 283386 319932
rect 283518 319880 283570 319932
rect 283748 319880 283800 319932
rect 283978 319880 284030 319932
rect 284346 319880 284398 319932
rect 284806 319880 284858 319932
rect 284898 319880 284950 319932
rect 281724 319812 281776 319864
rect 282690 319812 282742 319864
rect 283196 319676 283248 319728
rect 284760 319744 284812 319796
rect 284484 319676 284536 319728
rect 286370 319812 286422 319864
rect 286508 319744 286560 319796
rect 285036 319676 285088 319728
rect 285956 319676 286008 319728
rect 287474 319880 287526 319932
rect 289498 319880 289550 319932
rect 290050 319880 290102 319932
rect 291614 319880 291666 319932
rect 292718 319880 292770 319932
rect 287520 319744 287572 319796
rect 289452 319744 289504 319796
rect 290004 319744 290056 319796
rect 291568 319676 291620 319728
rect 269764 319608 269816 319660
rect 293822 319880 293874 319932
rect 294558 319880 294610 319932
rect 295202 319880 295254 319932
rect 295294 319880 295346 319932
rect 293914 319812 293966 319864
rect 294328 319812 294380 319864
rect 293776 319744 293828 319796
rect 295156 319676 295208 319728
rect 293868 319608 293920 319660
rect 293960 319608 294012 319660
rect 295754 319880 295806 319932
rect 295524 319676 295576 319728
rect 296306 319880 296358 319932
rect 296582 319880 296634 319932
rect 264336 319540 264388 319592
rect 296536 319540 296588 319592
rect 252744 319472 252796 319524
rect 298330 319880 298382 319932
rect 298698 319880 298750 319932
rect 298790 319880 298842 319932
rect 299250 319880 299302 319932
rect 298284 319676 298336 319728
rect 299158 319812 299210 319864
rect 298744 319608 298796 319660
rect 298560 319540 298612 319592
rect 237472 319404 237524 319456
rect 295340 319404 295392 319456
rect 295708 319404 295760 319456
rect 296076 319404 296128 319456
rect 300078 319812 300130 319864
rect 299388 319540 299440 319592
rect 301274 319880 301326 319932
rect 301366 319880 301418 319932
rect 301734 319880 301786 319932
rect 301918 319880 301970 319932
rect 303298 319880 303350 319932
rect 303482 319880 303534 319932
rect 301458 319812 301510 319864
rect 301320 319744 301372 319796
rect 301412 319676 301464 319728
rect 300216 319540 300268 319592
rect 300768 319540 300820 319592
rect 301596 319540 301648 319592
rect 301872 319676 301924 319728
rect 302700 319676 302752 319728
rect 303758 319880 303810 319932
rect 304034 319880 304086 319932
rect 303804 319744 303856 319796
rect 303436 319676 303488 319728
rect 302424 319608 302476 319660
rect 302608 319608 302660 319660
rect 301964 319540 302016 319592
rect 302148 319540 302200 319592
rect 304264 319540 304316 319592
rect 304862 319880 304914 319932
rect 305230 319880 305282 319932
rect 305322 319880 305374 319932
rect 305506 319880 305558 319932
rect 304770 319812 304822 319864
rect 305414 319812 305466 319864
rect 305184 319744 305236 319796
rect 305276 319744 305328 319796
rect 305368 319676 305420 319728
rect 304724 319540 304776 319592
rect 299296 319404 299348 319456
rect 300860 319404 300912 319456
rect 301044 319404 301096 319456
rect 301320 319404 301372 319456
rect 301596 319404 301648 319456
rect 305368 319404 305420 319456
rect 305966 319880 306018 319932
rect 306518 319880 306570 319932
rect 306702 319880 306754 319932
rect 305920 319608 305972 319660
rect 306472 319608 306524 319660
rect 308496 319880 308548 319932
rect 309094 319880 309146 319932
rect 308312 319812 308364 319864
rect 308956 319608 309008 319660
rect 327632 320764 327684 320816
rect 328184 320628 328236 320680
rect 338580 320560 338632 320612
rect 327724 320424 327776 320476
rect 336740 320424 336792 320476
rect 338304 320356 338356 320408
rect 309278 319880 309330 319932
rect 309370 319880 309422 319932
rect 309554 319880 309606 319932
rect 309830 319880 309882 319932
rect 310290 319880 310342 319932
rect 310934 319880 310986 319932
rect 311118 319880 311170 319932
rect 311486 319880 311538 319932
rect 309324 319744 309376 319796
rect 309784 319744 309836 319796
rect 309692 319676 309744 319728
rect 310244 319676 310296 319728
rect 311256 319676 311308 319728
rect 309232 319608 309284 319660
rect 309876 319608 309928 319660
rect 306932 319540 306984 319592
rect 307484 319540 307536 319592
rect 310888 319472 310940 319524
rect 311854 319812 311906 319864
rect 312314 319880 312366 319932
rect 313050 319880 313102 319932
rect 313418 319880 313470 319932
rect 313786 319880 313838 319932
rect 312590 319812 312642 319864
rect 312682 319812 312734 319864
rect 312774 319812 312826 319864
rect 312866 319812 312918 319864
rect 312268 319744 312320 319796
rect 312544 319676 312596 319728
rect 312360 319608 312412 319660
rect 312728 319608 312780 319660
rect 313096 319608 313148 319660
rect 311900 319540 311952 319592
rect 312820 319540 312872 319592
rect 309968 319404 310020 319456
rect 310152 319404 310204 319456
rect 310796 319404 310848 319456
rect 251456 319336 251508 319388
rect 311348 319336 311400 319388
rect 311624 319404 311676 319456
rect 312268 319404 312320 319456
rect 312636 319404 312688 319456
rect 312912 319404 312964 319456
rect 313280 319404 313332 319456
rect 313464 319404 313516 319456
rect 313878 319812 313930 319864
rect 314062 319812 314114 319864
rect 336832 320288 336884 320340
rect 327632 320220 327684 320272
rect 335820 320220 335872 320272
rect 327540 320152 327592 320204
rect 335912 320152 335964 320204
rect 321698 320084 321750 320136
rect 331404 320084 331456 320136
rect 320870 320016 320922 320068
rect 332968 320016 333020 320068
rect 314798 319880 314850 319932
rect 315442 319880 315494 319932
rect 315626 319880 315678 319932
rect 316914 319880 316966 319932
rect 317006 319880 317058 319932
rect 319582 319880 319634 319932
rect 314200 319540 314252 319592
rect 313924 319472 313976 319524
rect 315304 319608 315356 319660
rect 316408 319812 316460 319864
rect 316638 319812 316690 319864
rect 316224 319676 316276 319728
rect 317144 319744 317196 319796
rect 315672 319608 315724 319660
rect 316040 319608 316092 319660
rect 318202 319812 318254 319864
rect 318892 319812 318944 319864
rect 319260 319812 319312 319864
rect 320318 319812 320370 319864
rect 320686 319880 320738 319932
rect 320594 319812 320646 319864
rect 333060 319948 333112 320000
rect 323538 319880 323590 319932
rect 323216 319744 323268 319796
rect 320272 319676 320324 319728
rect 320364 319676 320416 319728
rect 338212 319744 338264 319796
rect 320640 319608 320692 319660
rect 328460 319608 328512 319660
rect 314660 319336 314712 319388
rect 243084 319268 243136 319320
rect 302516 319268 302568 319320
rect 309784 319268 309836 319320
rect 316040 319268 316092 319320
rect 248696 319200 248748 319252
rect 309324 319200 309376 319252
rect 311716 319200 311768 319252
rect 311900 319200 311952 319252
rect 248604 319132 248656 319184
rect 309232 319132 309284 319184
rect 322112 319472 322164 319524
rect 323032 319472 323084 319524
rect 323492 319472 323544 319524
rect 340880 319676 340932 319728
rect 316500 319404 316552 319456
rect 325884 319404 325936 319456
rect 326068 319404 326120 319456
rect 322388 319336 322440 319388
rect 336004 319404 336056 319456
rect 580448 319404 580500 319456
rect 337016 319336 337068 319388
rect 283472 319064 283524 319116
rect 292120 319064 292172 319116
rect 275284 318996 275336 319048
rect 294604 318996 294656 319048
rect 295708 318996 295760 319048
rect 296444 318996 296496 319048
rect 296536 318996 296588 319048
rect 310704 319064 310756 319116
rect 338488 319268 338540 319320
rect 321284 319200 321336 319252
rect 331588 319200 331640 319252
rect 314292 318996 314344 319048
rect 332876 319132 332928 319184
rect 272984 318928 273036 318980
rect 297364 318928 297416 318980
rect 309048 318928 309100 318980
rect 331220 319064 331272 319116
rect 325332 318996 325384 319048
rect 325516 318996 325568 319048
rect 326068 318996 326120 319048
rect 326620 318996 326672 319048
rect 322572 318928 322624 318980
rect 331956 318928 332008 318980
rect 279884 318860 279936 318912
rect 295524 318860 295576 318912
rect 318248 318860 318300 318912
rect 318432 318860 318484 318912
rect 320272 318860 320324 318912
rect 330392 318860 330444 318912
rect 3424 318792 3476 318844
rect 278044 318792 278096 318844
rect 284208 318792 284260 318844
rect 286692 318792 286744 318844
rect 286876 318792 286928 318844
rect 288716 318792 288768 318844
rect 289728 318792 289780 318844
rect 290924 318792 290976 318844
rect 291108 318792 291160 318844
rect 292120 318792 292172 318844
rect 258172 318724 258224 318776
rect 258816 318724 258868 318776
rect 285036 318724 285088 318776
rect 285220 318724 285272 318776
rect 286324 318724 286376 318776
rect 287520 318724 287572 318776
rect 289452 318724 289504 318776
rect 289636 318724 289688 318776
rect 292948 318792 293000 318844
rect 293868 318792 293920 318844
rect 298100 318792 298152 318844
rect 298284 318792 298336 318844
rect 302976 318792 303028 318844
rect 303252 318792 303304 318844
rect 322204 318792 322256 318844
rect 330024 318792 330076 318844
rect 293040 318724 293092 318776
rect 293316 318724 293368 318776
rect 293684 318724 293736 318776
rect 279608 318656 279660 318708
rect 301044 318724 301096 318776
rect 318432 318724 318484 318776
rect 318800 318724 318852 318776
rect 319904 318724 319956 318776
rect 329840 318724 329892 318776
rect 294052 318656 294104 318708
rect 294788 318656 294840 318708
rect 295892 318656 295944 318708
rect 300768 318656 300820 318708
rect 319996 318656 320048 318708
rect 330116 318656 330168 318708
rect 277584 318588 277636 318640
rect 278412 318588 278464 318640
rect 282184 318588 282236 318640
rect 285404 318588 285456 318640
rect 287796 318588 287848 318640
rect 294972 318588 295024 318640
rect 298284 318588 298336 318640
rect 299388 318588 299440 318640
rect 301044 318588 301096 318640
rect 303804 318588 303856 318640
rect 312084 318588 312136 318640
rect 323492 318588 323544 318640
rect 324964 318588 325016 318640
rect 325608 318588 325660 318640
rect 326344 318588 326396 318640
rect 334532 318588 334584 318640
rect 272892 318520 272944 318572
rect 294052 318520 294104 318572
rect 295156 318520 295208 318572
rect 295616 318520 295668 318572
rect 300860 318520 300912 318572
rect 317328 318520 317380 318572
rect 329104 318520 329156 318572
rect 247224 318452 247276 318504
rect 282828 318452 282880 318504
rect 238852 318384 238904 318436
rect 282276 318384 282328 318436
rect 282644 318384 282696 318436
rect 296628 318452 296680 318504
rect 302056 318452 302108 318504
rect 317972 318452 318024 318504
rect 325608 318452 325660 318504
rect 325792 318452 325844 318504
rect 335728 318452 335780 318504
rect 289452 318384 289504 318436
rect 209688 318316 209740 318368
rect 283748 318316 283800 318368
rect 284852 318316 284904 318368
rect 285128 318316 285180 318368
rect 291936 318316 291988 318368
rect 294420 318316 294472 318368
rect 295156 318384 295208 318436
rect 303436 318384 303488 318436
rect 317420 318384 317472 318436
rect 326528 318384 326580 318436
rect 297088 318316 297140 318368
rect 300860 318316 300912 318368
rect 302240 318316 302292 318368
rect 318892 318316 318944 318368
rect 335544 318316 335596 318368
rect 212264 318248 212316 318300
rect 286232 318248 286284 318300
rect 292120 318248 292172 318300
rect 299940 318248 299992 318300
rect 300216 318248 300268 318300
rect 300768 318248 300820 318300
rect 311808 318248 311860 318300
rect 326344 318248 326396 318300
rect 218980 318112 219032 318164
rect 287244 318180 287296 318232
rect 288808 318180 288860 318232
rect 289268 318180 289320 318232
rect 290740 318180 290792 318232
rect 298100 318180 298152 318232
rect 299296 318180 299348 318232
rect 306656 318180 306708 318232
rect 319352 318180 319404 318232
rect 286232 318112 286284 318164
rect 286784 318112 286836 318164
rect 219072 318044 219124 318096
rect 287796 318044 287848 318096
rect 287244 317976 287296 318028
rect 295984 318112 296036 318164
rect 300216 318112 300268 318164
rect 302792 318112 302844 318164
rect 316592 318112 316644 318164
rect 294052 318044 294104 318096
rect 301780 318044 301832 318096
rect 288808 317976 288860 318028
rect 289084 317976 289136 318028
rect 295340 317976 295392 318028
rect 301504 317976 301556 318028
rect 309784 317976 309836 318028
rect 312544 317976 312596 318028
rect 313372 317976 313424 318028
rect 278136 317908 278188 317960
rect 295432 317908 295484 317960
rect 303436 317908 303488 317960
rect 304356 317908 304408 317960
rect 311808 317908 311860 317960
rect 314016 317908 314068 317960
rect 322388 317908 322440 317960
rect 326436 318180 326488 318232
rect 340972 318180 341024 318232
rect 326528 318112 326580 318164
rect 349252 318112 349304 318164
rect 354680 318044 354732 318096
rect 325608 317976 325660 318028
rect 330576 317976 330628 318028
rect 326436 317908 326488 317960
rect 286784 317840 286836 317892
rect 293408 317840 293460 317892
rect 293868 317840 293920 317892
rect 298468 317840 298520 317892
rect 312268 317840 312320 317892
rect 326528 317840 326580 317892
rect 283748 317772 283800 317824
rect 292304 317772 292356 317824
rect 294788 317772 294840 317824
rect 298744 317772 298796 317824
rect 300032 317772 300084 317824
rect 300308 317772 300360 317824
rect 301412 317772 301464 317824
rect 302884 317772 302936 317824
rect 221740 317704 221792 317756
rect 296628 317704 296680 317756
rect 297364 317704 297416 317756
rect 301136 317704 301188 317756
rect 301228 317704 301280 317756
rect 303804 317772 303856 317824
rect 276940 317636 276992 317688
rect 295340 317636 295392 317688
rect 296260 317636 296312 317688
rect 299572 317636 299624 317688
rect 301964 317636 302016 317688
rect 307116 317704 307168 317756
rect 303988 317636 304040 317688
rect 305276 317636 305328 317688
rect 305828 317636 305880 317688
rect 320732 317636 320784 317688
rect 321376 317636 321428 317688
rect 280620 317568 280672 317620
rect 283748 317568 283800 317620
rect 283932 317568 283984 317620
rect 290648 317568 290700 317620
rect 293408 317568 293460 317620
rect 295064 317568 295116 317620
rect 296076 317568 296128 317620
rect 298376 317568 298428 317620
rect 300308 317568 300360 317620
rect 306104 317568 306156 317620
rect 306288 317568 306340 317620
rect 308496 317568 308548 317620
rect 308956 317568 309008 317620
rect 323400 317568 323452 317620
rect 327816 317568 327868 317620
rect 283656 317500 283708 317552
rect 289544 317500 289596 317552
rect 272800 317432 272852 317484
rect 295892 317500 295944 317552
rect 298192 317500 298244 317552
rect 300124 317500 300176 317552
rect 303068 317500 303120 317552
rect 305460 317500 305512 317552
rect 305828 317500 305880 317552
rect 308036 317500 308088 317552
rect 313280 317500 313332 317552
rect 320732 317500 320784 317552
rect 324412 317500 324464 317552
rect 327632 317500 327684 317552
rect 295340 317432 295392 317484
rect 297272 317432 297324 317484
rect 298836 317432 298888 317484
rect 300492 317432 300544 317484
rect 303804 317432 303856 317484
rect 303988 317432 304040 317484
rect 307576 317432 307628 317484
rect 308220 317432 308272 317484
rect 308956 317432 309008 317484
rect 309600 317432 309652 317484
rect 314568 317432 314620 317484
rect 315120 317432 315172 317484
rect 315672 317432 315724 317484
rect 317972 317432 318024 317484
rect 326160 317432 326212 317484
rect 327540 317432 327592 317484
rect 279792 317364 279844 317416
rect 302148 317364 302200 317416
rect 318708 317364 318760 317416
rect 323400 317364 323452 317416
rect 274180 317296 274232 317348
rect 296352 317296 296404 317348
rect 322940 317296 322992 317348
rect 328736 317296 328788 317348
rect 274272 317228 274324 317280
rect 296812 317228 296864 317280
rect 271420 317092 271472 317144
rect 295800 317092 295852 317144
rect 295984 317092 296036 317144
rect 305644 317092 305696 317144
rect 273996 317024 274048 317076
rect 303620 317024 303672 317076
rect 317696 317024 317748 317076
rect 334072 317024 334124 317076
rect 273168 316956 273220 317008
rect 303712 316956 303764 317008
rect 308864 316956 308916 317008
rect 328828 316956 328880 317008
rect 271512 316888 271564 316940
rect 302608 316888 302660 316940
rect 308312 316888 308364 316940
rect 329932 316888 329984 316940
rect 277308 316820 277360 316872
rect 313740 316820 313792 316872
rect 316684 316820 316736 316872
rect 336924 316820 336976 316872
rect 218796 316752 218848 316804
rect 294604 316752 294656 316804
rect 295248 316752 295300 316804
rect 305000 316752 305052 316804
rect 213368 316684 213420 316736
rect 293868 316684 293920 316736
rect 296628 316684 296680 316736
rect 282828 316616 282880 316668
rect 303436 316616 303488 316668
rect 308312 316684 308364 316736
rect 310796 316684 310848 316736
rect 364340 316752 364392 316804
rect 323584 316684 323636 316736
rect 400864 316684 400916 316736
rect 320456 316616 320508 316668
rect 276848 316548 276900 316600
rect 293960 316548 294012 316600
rect 280988 316480 281040 316532
rect 292396 316480 292448 316532
rect 271328 316412 271380 316464
rect 294328 316412 294380 316464
rect 325240 316412 325292 316464
rect 324964 316276 325016 316328
rect 327908 316276 327960 316328
rect 284300 316208 284352 316260
rect 284852 316208 284904 316260
rect 309600 316208 309652 316260
rect 310244 316208 310296 316260
rect 322204 316208 322256 316260
rect 323584 316208 323636 316260
rect 324044 316208 324096 316260
rect 284760 316140 284812 316192
rect 285496 316140 285548 316192
rect 306840 316140 306892 316192
rect 307024 316140 307076 316192
rect 323860 316140 323912 316192
rect 324136 316140 324188 316192
rect 325056 316140 325108 316192
rect 325240 316140 325292 316192
rect 493324 316208 493376 316260
rect 534080 316140 534132 316192
rect 283104 316072 283156 316124
rect 284116 316072 284168 316124
rect 284668 316072 284720 316124
rect 285588 316072 285640 316124
rect 287336 316072 287388 316124
rect 287888 316072 287940 316124
rect 288532 316072 288584 316124
rect 289360 316072 289412 316124
rect 290188 316072 290240 316124
rect 290464 316072 290516 316124
rect 283012 316004 283064 316056
rect 283840 316004 283892 316056
rect 284852 316004 284904 316056
rect 285312 316004 285364 316056
rect 285680 316004 285732 316056
rect 286876 316004 286928 316056
rect 287244 316004 287296 316056
rect 288164 316004 288216 316056
rect 288624 316004 288676 316056
rect 289176 316004 289228 316056
rect 289912 316004 289964 316056
rect 290740 316004 290792 316056
rect 291476 316004 291528 316056
rect 292028 316004 292080 316056
rect 275560 315936 275612 315988
rect 290648 315936 290700 315988
rect 276756 315868 276808 315920
rect 295616 316072 295668 316124
rect 309416 316072 309468 316124
rect 310244 316072 310296 316124
rect 311532 316072 311584 316124
rect 311716 316072 311768 316124
rect 315488 316072 315540 316124
rect 315764 316072 315816 316124
rect 323584 316072 323636 316124
rect 324044 316072 324096 316124
rect 325148 316072 325200 316124
rect 547972 316072 548024 316124
rect 294236 316004 294288 316056
rect 294512 316004 294564 316056
rect 294604 316004 294656 316056
rect 301044 316004 301096 316056
rect 303896 316004 303948 316056
rect 304816 316004 304868 316056
rect 306564 316004 306616 316056
rect 306840 316004 306892 316056
rect 307668 316004 307720 316056
rect 310796 316004 310848 316056
rect 311164 316004 311216 316056
rect 318800 316004 318852 316056
rect 319444 316004 319496 316056
rect 320180 316004 320232 316056
rect 320640 316004 320692 316056
rect 321652 316004 321704 316056
rect 322480 316004 322532 316056
rect 322848 316004 322900 316056
rect 327448 316004 327500 316056
rect 327908 316004 327960 316056
rect 554044 316004 554096 316056
rect 292856 315936 292908 315988
rect 293776 315936 293828 315988
rect 299756 315936 299808 315988
rect 300492 315936 300544 315988
rect 302516 315936 302568 315988
rect 303160 315936 303212 315988
rect 303804 315936 303856 315988
rect 304632 315936 304684 315988
rect 306380 315936 306432 315988
rect 306656 315936 306708 315988
rect 307392 315936 307444 315988
rect 308404 315936 308456 315988
rect 308864 315936 308916 315988
rect 310520 315936 310572 315988
rect 311532 315936 311584 315988
rect 312084 315936 312136 315988
rect 312452 315936 312504 315988
rect 312728 315936 312780 315988
rect 313004 315936 313056 315988
rect 313648 315936 313700 315988
rect 314292 315936 314344 315988
rect 315396 315936 315448 315988
rect 315764 315936 315816 315988
rect 319168 315936 319220 315988
rect 319720 315936 319772 315988
rect 320456 315936 320508 315988
rect 321008 315936 321060 315988
rect 321560 315936 321612 315988
rect 322756 315936 322808 315988
rect 324688 315936 324740 315988
rect 324872 315936 324924 315988
rect 325792 315936 325844 315988
rect 326252 315936 326304 315988
rect 327080 315936 327132 315988
rect 327264 315936 327316 315988
rect 306564 315868 306616 315920
rect 307300 315868 307352 315920
rect 308128 315868 308180 315920
rect 308772 315868 308824 315920
rect 309324 315868 309376 315920
rect 310336 315868 310388 315920
rect 321744 315868 321796 315920
rect 321928 315868 321980 315920
rect 323308 315868 323360 315920
rect 323952 315868 324004 315920
rect 274364 315800 274416 315852
rect 272708 315732 272760 315784
rect 292580 315732 292632 315784
rect 292764 315800 292816 315852
rect 293224 315800 293276 315852
rect 294420 315800 294472 315852
rect 294880 315800 294932 315852
rect 306196 315800 306248 315852
rect 307944 315800 307996 315852
rect 312452 315800 312504 315852
rect 312728 315800 312780 315852
rect 313464 315800 313516 315852
rect 314108 315800 314160 315852
rect 315212 315800 315264 315852
rect 315580 315800 315632 315852
rect 320548 315800 320600 315852
rect 321192 315800 321244 315852
rect 294052 315732 294104 315784
rect 294328 315732 294380 315784
rect 294696 315732 294748 315784
rect 307024 315732 307076 315784
rect 309416 315732 309468 315784
rect 312360 315732 312412 315784
rect 313188 315732 313240 315784
rect 274088 315664 274140 315716
rect 292396 315664 292448 315716
rect 293040 315664 293092 315716
rect 301688 315664 301740 315716
rect 306380 315664 306432 315716
rect 310888 315664 310940 315716
rect 271236 315596 271288 315648
rect 292304 315596 292356 315648
rect 294696 315596 294748 315648
rect 303528 315596 303580 315648
rect 307668 315596 307720 315648
rect 317788 315664 317840 315716
rect 311992 315596 312044 315648
rect 313188 315596 313240 315648
rect 268384 315528 268436 315580
rect 293960 315528 294012 315580
rect 294052 315528 294104 315580
rect 299940 315528 299992 315580
rect 302884 315528 302936 315580
rect 314844 315528 314896 315580
rect 272524 315460 272576 315512
rect 233056 315392 233108 315444
rect 282920 315392 282972 315444
rect 283564 315392 283616 315444
rect 284392 315392 284444 315444
rect 287612 315392 287664 315444
rect 288256 315392 288308 315444
rect 290004 315392 290056 315444
rect 290372 315392 290424 315444
rect 316776 315460 316828 315512
rect 293960 315392 294012 315444
rect 302056 315392 302108 315444
rect 308496 315392 308548 315444
rect 331312 315392 331364 315444
rect 217692 315324 217744 315376
rect 280160 315324 280212 315376
rect 287704 315324 287756 315376
rect 287980 315324 288032 315376
rect 288348 315324 288400 315376
rect 290280 315324 290332 315376
rect 292304 315324 292356 315376
rect 294696 315324 294748 315376
rect 309968 315324 310020 315376
rect 336004 315324 336056 315376
rect 215024 315256 215076 315308
rect 284300 315256 284352 315308
rect 284392 315256 284444 315308
rect 285036 315256 285088 315308
rect 287152 315256 287204 315308
rect 288256 315256 288308 315308
rect 288440 315256 288492 315308
rect 289544 315256 289596 315308
rect 291844 315256 291896 315308
rect 306104 315256 306156 315308
rect 279700 315188 279752 315240
rect 300676 315188 300728 315240
rect 303160 315188 303212 315240
rect 311072 315188 311124 315240
rect 367100 315256 367152 315308
rect 278688 315120 278740 315172
rect 295156 315120 295208 315172
rect 282920 315052 282972 315104
rect 288900 315052 288952 315104
rect 292580 315052 292632 315104
rect 299388 315052 299440 315104
rect 286416 314984 286468 315036
rect 287888 314984 287940 315036
rect 312636 314712 312688 314764
rect 396080 314712 396132 314764
rect 313924 314644 313976 314696
rect 407120 314644 407172 314696
rect 276664 314576 276716 314628
rect 290556 314576 290608 314628
rect 269856 314508 269908 314560
rect 290464 314508 290516 314560
rect 299112 314508 299164 314560
rect 299296 314508 299348 314560
rect 274548 314440 274600 314492
rect 295248 314440 295300 314492
rect 279424 314372 279476 314424
rect 304264 314372 304316 314424
rect 320916 314372 320968 314424
rect 328920 314372 328972 314424
rect 280896 314304 280948 314356
rect 315948 314304 316000 314356
rect 270040 314236 270092 314288
rect 319260 314236 319312 314288
rect 286876 314168 286928 314220
rect 298744 314168 298796 314220
rect 220544 314100 220596 314152
rect 292212 314100 292264 314152
rect 218888 314032 218940 314084
rect 291936 314032 291988 314084
rect 216312 313964 216364 314016
rect 297824 313964 297876 314016
rect 319628 314032 319680 314084
rect 330300 314032 330352 314084
rect 431960 313964 432012 314016
rect 216404 313896 216456 313948
rect 221832 313828 221884 313880
rect 286692 313828 286744 313880
rect 291660 313896 291712 313948
rect 292488 313896 292540 313948
rect 316960 313896 317012 313948
rect 441620 313896 441672 313948
rect 297732 313760 297784 313812
rect 315488 313760 315540 313812
rect 316960 313760 317012 313812
rect 290648 313624 290700 313676
rect 291200 313624 291252 313676
rect 300124 313352 300176 313404
rect 306012 313352 306064 313404
rect 315304 313352 315356 313404
rect 422944 313352 422996 313404
rect 268568 313284 268620 313336
rect 314108 313284 314160 313336
rect 315396 313284 315448 313336
rect 427820 313284 427872 313336
rect 293224 313216 293276 313268
rect 296536 313216 296588 313268
rect 313280 313216 313332 313268
rect 313832 313216 313884 313268
rect 296168 313148 296220 313200
rect 300032 313148 300084 313200
rect 271696 313080 271748 313132
rect 304540 313080 304592 313132
rect 278412 313012 278464 313064
rect 312820 313012 312872 313064
rect 275376 312944 275428 312996
rect 318064 312944 318116 312996
rect 252468 312876 252520 312928
rect 311348 312876 311400 312928
rect 235632 312808 235684 312860
rect 296444 312808 296496 312860
rect 297456 312808 297508 312860
rect 321100 312808 321152 312860
rect 235908 312740 235960 312792
rect 295892 312740 295944 312792
rect 309692 312740 309744 312792
rect 342260 312740 342312 312792
rect 216036 312672 216088 312724
rect 282552 312672 282604 312724
rect 216128 312604 216180 312656
rect 284024 312604 284076 312656
rect 215944 312536 215996 312588
rect 282552 312536 282604 312588
rect 315028 312672 315080 312724
rect 321100 312672 321152 312724
rect 500224 312672 500276 312724
rect 322296 312604 322348 312656
rect 511264 312604 511316 312656
rect 320916 312536 320968 312588
rect 323032 312536 323084 312588
rect 526444 312536 526496 312588
rect 286508 312468 286560 312520
rect 302976 312060 303028 312112
rect 303160 312060 303212 312112
rect 213828 311924 213880 311976
rect 288440 311992 288492 312044
rect 217508 311856 217560 311908
rect 292580 311924 292632 311976
rect 320824 311924 320876 311976
rect 322296 311924 322348 311976
rect 291936 311856 291988 311908
rect 293592 311856 293644 311908
rect 313280 311856 313332 311908
rect 409880 311856 409932 311908
rect 279516 311584 279568 311636
rect 288256 311584 288308 311636
rect 277216 311516 277268 311568
rect 303068 311516 303120 311568
rect 224592 311448 224644 311500
rect 283012 311448 283064 311500
rect 300124 311448 300176 311500
rect 300308 311448 300360 311500
rect 251088 311380 251140 311432
rect 309508 311380 309560 311432
rect 249616 311312 249668 311364
rect 309232 311312 309284 311364
rect 250996 311244 251048 311296
rect 310612 311244 310664 311296
rect 250720 311176 250772 311228
rect 311532 311176 311584 311228
rect 221648 311108 221700 311160
rect 280988 311108 281040 311160
rect 281264 311108 281316 311160
rect 282644 311108 282696 311160
rect 289452 311108 289504 311160
rect 294604 311108 294656 311160
rect 294788 311108 294840 311160
rect 298744 311108 298796 311160
rect 299112 311108 299164 311160
rect 300952 311108 301004 311160
rect 301964 311108 302016 311160
rect 314108 311108 314160 311160
rect 414020 311108 414072 311160
rect 284668 311040 284720 311092
rect 312360 310564 312412 310616
rect 312636 310564 312688 310616
rect 391940 310564 391992 310616
rect 324412 310496 324464 310548
rect 324780 310496 324832 310548
rect 543004 310496 543056 310548
rect 289176 310428 289228 310480
rect 293316 310428 293368 310480
rect 289268 310360 289320 310412
rect 295340 310360 295392 310412
rect 276020 310292 276072 310344
rect 285680 310292 285732 310344
rect 278228 310224 278280 310276
rect 288624 310224 288676 310276
rect 256516 310156 256568 310208
rect 314752 310156 314804 310208
rect 256608 310088 256660 310140
rect 317236 310088 317288 310140
rect 256240 310020 256292 310072
rect 316132 310020 316184 310072
rect 215760 309952 215812 310004
rect 281724 309952 281776 310004
rect 285036 309952 285088 310004
rect 318248 309952 318300 310004
rect 214932 309884 214984 309936
rect 284392 309884 284444 309936
rect 286508 309884 286560 309936
rect 318892 309884 318944 309936
rect 218612 309816 218664 309868
rect 291108 309816 291160 309868
rect 214564 309748 214616 309800
rect 290188 309748 290240 309800
rect 315580 309748 315632 309800
rect 327356 309748 327408 309800
rect 565820 309748 565872 309800
rect 282276 309476 282328 309528
rect 282552 309476 282604 309528
rect 282000 309340 282052 309392
rect 282552 309340 282604 309392
rect 217416 309204 217468 309256
rect 287152 309204 287204 309256
rect 213276 309136 213328 309188
rect 285680 309136 285732 309188
rect 327724 309136 327776 309188
rect 558920 309136 558972 309188
rect 214656 308456 214708 308508
rect 288808 308456 288860 308508
rect 289452 308456 289504 308508
rect 324412 308456 324464 308508
rect 210976 308388 211028 308440
rect 285956 308388 286008 308440
rect 313924 308388 313976 308440
rect 314936 308388 314988 308440
rect 416780 308388 416832 308440
rect 327816 307776 327868 307828
rect 523040 307776 523092 307828
rect 287888 307572 287940 307624
rect 296996 307572 297048 307624
rect 275836 307504 275888 307556
rect 288716 307504 288768 307556
rect 290556 307504 290608 307556
rect 293408 307504 293460 307556
rect 288348 307436 288400 307488
rect 303896 307436 303948 307488
rect 285588 307368 285640 307420
rect 303804 307368 303856 307420
rect 217324 307300 217376 307352
rect 276020 307300 276072 307352
rect 284208 307300 284260 307352
rect 304264 307300 304316 307352
rect 222200 307232 222252 307284
rect 283196 307232 283248 307284
rect 290464 307232 290516 307284
rect 315672 307232 315724 307284
rect 214748 307164 214800 307216
rect 285128 307164 285180 307216
rect 289360 307164 289412 307216
rect 313280 307164 313332 307216
rect 215852 307096 215904 307148
rect 285864 307096 285916 307148
rect 286692 307096 286744 307148
rect 321560 307096 321612 307148
rect 220360 307028 220412 307080
rect 294880 307028 294932 307080
rect 287796 306960 287848 307012
rect 294420 306960 294472 307012
rect 280896 306348 280948 306400
rect 289636 306348 289688 306400
rect 282092 306280 282144 306332
rect 580448 306348 580500 306400
rect 260288 305668 260340 305720
rect 282092 305668 282144 305720
rect 283748 305668 283800 305720
rect 304172 305668 304224 305720
rect 268660 305600 268712 305652
rect 327632 305600 327684 305652
rect 540980 305600 541032 305652
rect 3240 304988 3292 305040
rect 253112 304988 253164 305040
rect 247132 304444 247184 304496
rect 275100 304444 275152 304496
rect 218704 304376 218756 304428
rect 280620 304376 280672 304428
rect 220268 304308 220320 304360
rect 296904 304308 296956 304360
rect 220176 304240 220228 304292
rect 297548 304240 297600 304292
rect 314108 304240 314160 304292
rect 327540 304240 327592 304292
rect 563060 304240 563112 304292
rect 274456 302880 274508 302932
rect 318616 302880 318668 302932
rect 329656 302880 329708 302932
rect 245844 301928 245896 301980
rect 245752 301724 245804 301776
rect 253112 301724 253164 301776
rect 258816 301724 258868 301776
rect 240140 301520 240192 301572
rect 240324 301520 240376 301572
rect 221556 301452 221608 301504
rect 302516 301452 302568 301504
rect 329104 300840 329156 300892
rect 445760 300840 445812 300892
rect 258816 300772 258868 300824
rect 259092 300772 259144 300824
rect 275192 300772 275244 300824
rect 304264 300364 304316 300416
rect 305552 300364 305604 300416
rect 329656 300092 329708 300144
rect 452660 300092 452712 300144
rect 256792 299480 256844 299532
rect 257620 299480 257672 299532
rect 253940 298868 253992 298920
rect 254676 298868 254728 298920
rect 229468 298800 229520 298852
rect 242164 298800 242216 298852
rect 221464 298732 221516 298784
rect 302424 298732 302476 298784
rect 332048 298732 332100 298784
rect 572812 298732 572864 298784
rect 256700 297440 256752 297492
rect 257252 297440 257304 297492
rect 232964 297372 233016 297424
rect 277860 297372 277912 297424
rect 316684 297372 316736 297424
rect 330576 297372 330628 297424
rect 456800 297372 456852 297424
rect 255412 297304 255464 297356
rect 256332 297304 256384 297356
rect 256884 297304 256936 297356
rect 257068 297304 257120 297356
rect 226892 296692 226944 296744
rect 231124 296692 231176 296744
rect 244556 296012 244608 296064
rect 277952 296012 278004 296064
rect 222292 295944 222344 295996
rect 283380 295944 283432 295996
rect 258172 294652 258224 294704
rect 258540 294652 258592 294704
rect 235724 294584 235776 294636
rect 278596 294584 278648 294636
rect 318064 294584 318116 294636
rect 329196 294584 329248 294636
rect 463700 294584 463752 294636
rect 312176 293972 312228 294024
rect 312728 293972 312780 294024
rect 382280 293972 382332 294024
rect 248236 293904 248288 293956
rect 250444 293904 250496 293956
rect 233884 293564 233936 293616
rect 247592 293564 247644 293616
rect 231676 293496 231728 293548
rect 245016 293496 245068 293548
rect 228364 293428 228416 293480
rect 243544 293428 243596 293480
rect 236092 293360 236144 293412
rect 278504 293360 278556 293412
rect 223948 293292 224000 293344
rect 280712 293292 280764 293344
rect 3424 293224 3476 293276
rect 258724 293224 258776 293276
rect 334716 293224 334768 293276
rect 466460 293224 466512 293276
rect 223764 293020 223816 293072
rect 224500 293020 224552 293072
rect 225052 293020 225104 293072
rect 225972 293020 226024 293072
rect 226340 293020 226392 293072
rect 227076 293020 227128 293072
rect 230480 293020 230532 293072
rect 231124 293020 231176 293072
rect 236000 293020 236052 293072
rect 237012 293020 237064 293072
rect 241520 293020 241572 293072
rect 242164 293020 242216 293072
rect 242900 293020 242952 293072
rect 243268 293020 243320 293072
rect 245752 293020 245804 293072
rect 246580 293020 246632 293072
rect 247040 293020 247092 293072
rect 247684 293020 247736 293072
rect 249800 293020 249852 293072
rect 250260 293020 250312 293072
rect 251272 293020 251324 293072
rect 252100 293020 252152 293072
rect 252652 293020 252704 293072
rect 253204 293020 253256 293072
rect 242992 292952 243044 293004
rect 244004 292952 244056 293004
rect 252560 292952 252612 293004
rect 253572 292952 253624 293004
rect 220084 292544 220136 292596
rect 223948 292544 224000 292596
rect 319444 292544 319496 292596
rect 481640 292544 481692 292596
rect 238300 292476 238352 292528
rect 239404 292476 239456 292528
rect 259644 292476 259696 292528
rect 260196 292476 260248 292528
rect 262128 292476 262180 292528
rect 262588 292476 262640 292528
rect 264244 292476 264296 292528
rect 264796 292476 264848 292528
rect 234988 292136 235040 292188
rect 236552 292136 236604 292188
rect 236368 292068 236420 292120
rect 244924 292136 244976 292188
rect 234252 292000 234304 292052
rect 253112 292068 253164 292120
rect 232044 291932 232096 291984
rect 260288 292000 260340 292052
rect 263692 292000 263744 292052
rect 275928 292000 275980 292052
rect 237564 291932 237616 291984
rect 281080 291932 281132 291984
rect 235356 291864 235408 291916
rect 281172 291864 281224 291916
rect 318248 291864 318300 291916
rect 331680 291864 331732 291916
rect 217232 291796 217284 291848
rect 262588 291796 262640 291848
rect 265900 291796 265952 291848
rect 329012 291796 329064 291848
rect 470600 291796 470652 291848
rect 262312 291728 262364 291780
rect 262772 291728 262824 291780
rect 198004 291660 198056 291712
rect 263692 291660 263744 291712
rect 195244 291592 195296 291644
rect 264796 291592 264848 291644
rect 225052 291524 225104 291576
rect 226984 291524 227036 291576
rect 232228 291524 232280 291576
rect 259644 291524 259696 291576
rect 226524 291456 226576 291508
rect 256148 291456 256200 291508
rect 220912 291388 220964 291440
rect 260104 291388 260156 291440
rect 219900 291320 219952 291372
rect 261484 291320 261536 291372
rect 222016 291252 222068 291304
rect 222108 291184 222160 291236
rect 224224 291184 224276 291236
rect 225420 291184 225472 291236
rect 225604 291184 225656 291236
rect 230940 291184 230992 291236
rect 281356 291116 281408 291168
rect 264888 290844 264940 290896
rect 265532 290844 265584 290896
rect 239772 290640 239824 290692
rect 255964 290640 256016 290692
rect 240876 290572 240928 290624
rect 257344 290572 257396 290624
rect 116584 290504 116636 290556
rect 264888 290504 264940 290556
rect 3516 290436 3568 290488
rect 232228 290436 232280 290488
rect 243820 290436 243872 290488
rect 275744 290436 275796 290488
rect 281356 290436 281408 290488
rect 580724 290436 580776 290488
rect 219992 290096 220044 290148
rect 259828 290096 259880 290148
rect 262496 290096 262548 290148
rect 263324 290096 263376 290148
rect 229284 290028 229336 290080
rect 229744 290028 229796 290080
rect 269948 290028 270000 290080
rect 213460 289960 213512 290012
rect 260932 289960 260984 290012
rect 203524 289892 203576 289944
rect 262128 289892 262180 289944
rect 192484 289824 192536 289876
rect 262496 289824 262548 289876
rect 256148 289756 256200 289808
rect 256516 289756 256568 289808
rect 259552 289756 259604 289808
rect 260564 289756 260616 289808
rect 261300 289756 261352 289808
rect 261668 289756 261720 289808
rect 249248 289620 249300 289672
rect 211804 289212 211856 289264
rect 249248 289484 249300 289536
rect 199384 289144 199436 289196
rect 222476 289144 222528 289196
rect 91744 289076 91796 289128
rect 259552 289484 259604 289536
rect 262772 289552 262824 289604
rect 261300 289484 261352 289536
rect 222476 288804 222528 288856
rect 3424 286288 3476 286340
rect 220912 286288 220964 286340
rect 270224 284928 270276 284980
rect 290924 284928 290976 284980
rect 271788 283568 271840 283620
rect 284576 283568 284628 283620
rect 271052 282140 271104 282192
rect 286048 282140 286100 282192
rect 270316 275272 270368 275324
rect 290740 275272 290792 275324
rect 270960 273912 271012 273964
rect 283472 273912 283524 273964
rect 330484 273164 330536 273216
rect 580172 273164 580224 273216
rect 320548 271804 320600 271856
rect 321100 271804 321152 271856
rect 321100 270512 321152 270564
rect 498200 270512 498252 270564
rect 313464 269016 313516 269068
rect 314200 269016 314252 269068
rect 314200 267724 314252 267776
rect 407212 267724 407264 267776
rect 319076 265820 319128 265872
rect 319628 265820 319680 265872
rect 319628 264936 319680 264988
rect 467840 264936 467892 264988
rect 270408 264188 270460 264240
rect 291568 264188 291620 264240
rect 312084 263576 312136 263628
rect 313464 263576 313516 263628
rect 386420 263576 386472 263628
rect 316316 262624 316368 262676
rect 316776 262624 316828 262676
rect 316776 262216 316828 262268
rect 438860 262216 438912 262268
rect 269672 260108 269724 260160
rect 290832 260108 290884 260160
rect 306840 260108 306892 260160
rect 320548 260108 320600 260160
rect 349160 259428 349212 259480
rect 308956 259360 309008 259412
rect 309508 259360 309560 259412
rect 313372 259360 313424 259412
rect 314384 259360 314436 259412
rect 320456 259360 320508 259412
rect 321008 259360 321060 259412
rect 363604 259360 363656 259412
rect 579804 259360 579856 259412
rect 314384 258136 314436 258188
rect 402980 258136 403032 258188
rect 321008 258068 321060 258120
rect 496820 258068 496872 258120
rect 319536 255280 319588 255332
rect 320088 255280 320140 255332
rect 481732 255280 481784 255332
rect 314568 253920 314620 253972
rect 314844 253920 314896 253972
rect 420920 253920 420972 253972
rect 3516 253172 3568 253224
rect 219900 253172 219952 253224
rect 321928 252560 321980 252612
rect 322296 252560 322348 252612
rect 510620 252560 510672 252612
rect 321836 252492 321888 252544
rect 322572 252492 322624 252544
rect 269580 251812 269632 251864
rect 291476 251812 291528 251864
rect 322572 251200 322624 251252
rect 506480 251200 506532 251252
rect 312912 250452 312964 250504
rect 326436 250452 326488 250504
rect 385040 250452 385092 250504
rect 314292 249024 314344 249076
rect 322388 249024 322440 249076
rect 398840 249024 398892 249076
rect 312820 248412 312872 248464
rect 389180 248412 389232 248464
rect 321744 247868 321796 247920
rect 322388 247868 322440 247920
rect 316224 247120 316276 247172
rect 443000 247120 443052 247172
rect 322388 247052 322440 247104
rect 506572 247052 506624 247104
rect 269120 246304 269172 246356
rect 324136 246304 324188 246356
rect 309048 245760 309100 245812
rect 346400 245760 346452 245812
rect 320364 245692 320416 245744
rect 321284 245692 321336 245744
rect 491300 245692 491352 245744
rect 321192 245624 321244 245676
rect 321468 245624 321520 245676
rect 499580 245624 499632 245676
rect 310796 245148 310848 245200
rect 311256 245148 311308 245200
rect 268936 244944 268988 244996
rect 284484 244944 284536 244996
rect 269212 244876 269264 244928
rect 323676 244876 323728 244928
rect 311256 244332 311308 244384
rect 371240 244332 371292 244384
rect 322480 244264 322532 244316
rect 503720 244264 503772 244316
rect 269028 243516 269080 243568
rect 325700 243516 325752 243568
rect 321376 242904 321428 242956
rect 492680 242904 492732 242956
rect 215760 241476 215812 241528
rect 221004 241476 221056 241528
rect 3424 241408 3476 241460
rect 219992 241408 220044 241460
rect 220360 241000 220412 241052
rect 218796 240932 218848 240984
rect 202880 240864 202932 240916
rect 220360 240864 220412 240916
rect 193220 240796 193272 240848
rect 220176 240796 220228 240848
rect 222292 240864 222344 240916
rect 161480 240728 161532 240780
rect 218796 240728 218848 240780
rect 219256 240592 219308 240644
rect 220820 240592 220872 240644
rect 221372 240728 221424 240780
rect 221832 240728 221884 240780
rect 221740 240660 221792 240712
rect 222292 240592 222344 240644
rect 214380 240456 214432 240508
rect 218704 240456 218756 240508
rect 219164 240456 219216 240508
rect 221188 240456 221240 240508
rect 214472 240388 214524 240440
rect 215576 240320 215628 240372
rect 217692 240252 217744 240304
rect 221096 240252 221148 240304
rect 222292 240252 222344 240304
rect 216220 240184 216272 240236
rect 221740 240184 221792 240236
rect 210424 240048 210476 240100
rect 219348 240048 219400 240100
rect 222200 240048 222252 240100
rect 222292 239980 222344 240032
rect 207020 239912 207072 239964
rect 213368 239912 213420 239964
rect 216312 239844 216364 239896
rect 216588 239844 216640 239896
rect 219164 239844 219216 239896
rect 219348 239844 219400 239896
rect 197360 239776 197412 239828
rect 220268 239776 220320 239828
rect 221924 239912 221976 239964
rect 222384 239912 222436 239964
rect 222890 239912 222942 239964
rect 223350 239912 223402 239964
rect 223442 239912 223494 239964
rect 221004 239844 221056 239896
rect 221280 239776 221332 239828
rect 222706 239844 222758 239896
rect 222798 239844 222850 239896
rect 223166 239844 223218 239896
rect 182180 239708 182232 239760
rect 219164 239708 219216 239760
rect 219256 239708 219308 239760
rect 222200 239708 222252 239760
rect 222752 239708 222804 239760
rect 175280 239640 175332 239692
rect 218980 239640 219032 239692
rect 219348 239640 219400 239692
rect 223120 239640 223172 239692
rect 139400 239572 139452 239624
rect 125600 239504 125652 239556
rect 214380 239504 214432 239556
rect 103520 239436 103572 239488
rect 214564 239436 214616 239488
rect 215576 239436 215628 239488
rect 217968 239572 218020 239624
rect 222292 239572 222344 239624
rect 223718 239912 223770 239964
rect 223534 239776 223586 239828
rect 223396 239640 223448 239692
rect 223580 239640 223632 239692
rect 223902 239844 223954 239896
rect 223994 239844 224046 239896
rect 223856 239640 223908 239692
rect 223488 239572 223540 239624
rect 224546 239912 224598 239964
rect 224638 239912 224690 239964
rect 224730 239912 224782 239964
rect 224822 239912 224874 239964
rect 225006 239912 225058 239964
rect 224270 239844 224322 239896
rect 224362 239844 224414 239896
rect 224316 239708 224368 239760
rect 224592 239776 224644 239828
rect 224730 239776 224782 239828
rect 225282 239912 225334 239964
rect 225374 239912 225426 239964
rect 225558 239912 225610 239964
rect 225650 239912 225702 239964
rect 226202 239912 226254 239964
rect 226938 239912 226990 239964
rect 227030 239912 227082 239964
rect 225144 239708 225196 239760
rect 225236 239640 225288 239692
rect 226110 239844 226162 239896
rect 226570 239844 226622 239896
rect 226662 239844 226714 239896
rect 226754 239844 226806 239896
rect 225604 239776 225656 239828
rect 224224 239572 224276 239624
rect 224500 239572 224552 239624
rect 224776 239572 224828 239624
rect 225328 239572 225380 239624
rect 225512 239572 225564 239624
rect 226064 239572 226116 239624
rect 226616 239640 226668 239692
rect 226892 239708 226944 239760
rect 226800 239640 226852 239692
rect 226708 239572 226760 239624
rect 226892 239572 226944 239624
rect 227214 239844 227266 239896
rect 227122 239708 227174 239760
rect 227398 239912 227450 239964
rect 227766 239912 227818 239964
rect 228134 239912 228186 239964
rect 227490 239844 227542 239896
rect 227582 239844 227634 239896
rect 227536 239708 227588 239760
rect 227352 239640 227404 239692
rect 215944 239504 215996 239556
rect 227076 239504 227128 239556
rect 227168 239504 227220 239556
rect 227260 239504 227312 239556
rect 228042 239844 228094 239896
rect 227720 239572 227772 239624
rect 228226 239844 228278 239896
rect 228180 239640 228232 239692
rect 228686 239912 228738 239964
rect 228870 239912 228922 239964
rect 228962 239912 229014 239964
rect 229974 239912 230026 239964
rect 230250 239912 230302 239964
rect 230526 239912 230578 239964
rect 228594 239844 228646 239896
rect 228548 239708 228600 239760
rect 228824 239708 228876 239760
rect 229054 239844 229106 239896
rect 229606 239844 229658 239896
rect 229008 239708 229060 239760
rect 228640 239572 228692 239624
rect 228732 239572 228784 239624
rect 229192 239572 229244 239624
rect 230066 239844 230118 239896
rect 230342 239844 230394 239896
rect 230020 239708 230072 239760
rect 230112 239708 230164 239760
rect 230296 239708 230348 239760
rect 230388 239708 230440 239760
rect 230388 239572 230440 239624
rect 230802 239912 230854 239964
rect 230894 239844 230946 239896
rect 230756 239572 230808 239624
rect 231262 239912 231314 239964
rect 231354 239912 231406 239964
rect 231446 239912 231498 239964
rect 231630 239912 231682 239964
rect 232458 239912 232510 239964
rect 231814 239844 231866 239896
rect 231906 239844 231958 239896
rect 232090 239844 232142 239896
rect 231492 239708 231544 239760
rect 231584 239708 231636 239760
rect 231768 239708 231820 239760
rect 231032 239572 231084 239624
rect 231308 239572 231360 239624
rect 231952 239572 232004 239624
rect 228180 239504 228232 239556
rect 228364 239504 228416 239556
rect 230572 239504 230624 239556
rect 232734 239912 232786 239964
rect 232826 239912 232878 239964
rect 233010 239912 233062 239964
rect 233194 239912 233246 239964
rect 233286 239912 233338 239964
rect 233470 239912 233522 239964
rect 233838 239912 233890 239964
rect 234022 239912 234074 239964
rect 234390 239912 234442 239964
rect 232596 239640 232648 239692
rect 232780 239776 232832 239828
rect 232964 239708 233016 239760
rect 233148 239640 233200 239692
rect 232136 239572 232188 239624
rect 232688 239572 232740 239624
rect 232228 239504 232280 239556
rect 220636 239436 220688 239488
rect 233746 239844 233798 239896
rect 233700 239708 233752 239760
rect 233516 239572 233568 239624
rect 233792 239572 233844 239624
rect 234344 239640 234396 239692
rect 234850 239912 234902 239964
rect 235034 239912 235086 239964
rect 235310 239912 235362 239964
rect 235494 239912 235546 239964
rect 235862 239912 235914 239964
rect 236046 239912 236098 239964
rect 235218 239844 235270 239896
rect 234896 239708 234948 239760
rect 235172 239708 235224 239760
rect 235264 239640 235316 239692
rect 234620 239572 234672 239624
rect 235770 239844 235822 239896
rect 235908 239708 235960 239760
rect 235816 239640 235868 239692
rect 233976 239504 234028 239556
rect 235448 239504 235500 239556
rect 3424 239368 3476 239420
rect 217232 239368 217284 239420
rect 218704 239368 218756 239420
rect 219072 239368 219124 239420
rect 219348 239368 219400 239420
rect 236230 239912 236282 239964
rect 236322 239912 236374 239964
rect 236690 239912 236742 239964
rect 236782 239912 236834 239964
rect 237242 239912 237294 239964
rect 237518 239912 237570 239964
rect 237794 239912 237846 239964
rect 237978 239912 238030 239964
rect 238070 239912 238122 239964
rect 238254 239912 238306 239964
rect 239082 239912 239134 239964
rect 236184 239504 236236 239556
rect 178040 239300 178092 239352
rect 236506 239844 236558 239896
rect 236552 239708 236604 239760
rect 236552 239572 236604 239624
rect 237058 239844 237110 239896
rect 237012 239708 237064 239760
rect 237748 239776 237800 239828
rect 237656 239640 237708 239692
rect 237748 239640 237800 239692
rect 238806 239844 238858 239896
rect 238898 239844 238950 239896
rect 238530 239776 238582 239828
rect 237288 239572 237340 239624
rect 238024 239572 238076 239624
rect 236736 239504 236788 239556
rect 238944 239640 238996 239692
rect 238760 239572 238812 239624
rect 238392 239504 238444 239556
rect 238484 239504 238536 239556
rect 238852 239504 238904 239556
rect 239174 239844 239226 239896
rect 239450 239912 239502 239964
rect 239542 239912 239594 239964
rect 239726 239912 239778 239964
rect 239818 239912 239870 239964
rect 240002 239912 240054 239964
rect 240186 239912 240238 239964
rect 240738 239912 240790 239964
rect 240922 239912 240974 239964
rect 239358 239844 239410 239896
rect 239128 239708 239180 239760
rect 239220 239708 239272 239760
rect 239496 239776 239548 239828
rect 239772 239776 239824 239828
rect 240094 239844 240146 239896
rect 239956 239708 240008 239760
rect 240278 239844 240330 239896
rect 240140 239708 240192 239760
rect 240692 239708 240744 239760
rect 240048 239640 240100 239692
rect 240232 239640 240284 239692
rect 239496 239572 239548 239624
rect 239404 239504 239456 239556
rect 236460 239436 236512 239488
rect 241198 239912 241250 239964
rect 241290 239844 241342 239896
rect 241244 239708 241296 239760
rect 241152 239572 241204 239624
rect 241474 239912 241526 239964
rect 241934 239912 241986 239964
rect 242026 239912 242078 239964
rect 241336 239504 241388 239556
rect 241842 239844 241894 239896
rect 241888 239640 241940 239692
rect 242302 239912 242354 239964
rect 242394 239912 242446 239964
rect 242578 239912 242630 239964
rect 243406 239912 243458 239964
rect 243498 239912 243550 239964
rect 243958 239912 244010 239964
rect 244326 239912 244378 239964
rect 244510 239912 244562 239964
rect 244602 239912 244654 239964
rect 245062 239912 245114 239964
rect 242440 239708 242492 239760
rect 242532 239640 242584 239692
rect 242946 239844 242998 239896
rect 243222 239844 243274 239896
rect 242992 239708 243044 239760
rect 242164 239572 242216 239624
rect 242808 239572 242860 239624
rect 241612 239504 241664 239556
rect 242532 239436 242584 239488
rect 242716 239436 242768 239488
rect 242992 239436 243044 239488
rect 243452 239776 243504 239828
rect 244142 239844 244194 239896
rect 244372 239708 244424 239760
rect 244096 239640 244148 239692
rect 244188 239640 244240 239692
rect 243360 239572 243412 239624
rect 244694 239844 244746 239896
rect 244878 239844 244930 239896
rect 244924 239708 244976 239760
rect 245338 239912 245390 239964
rect 245430 239912 245482 239964
rect 245522 239912 245574 239964
rect 245706 239912 245758 239964
rect 245200 239640 245252 239692
rect 244740 239572 244792 239624
rect 245384 239776 245436 239828
rect 245568 239640 245620 239692
rect 245660 239640 245712 239692
rect 246166 239912 246218 239964
rect 246258 239912 246310 239964
rect 246350 239912 246402 239964
rect 246534 239912 246586 239964
rect 246810 239912 246862 239964
rect 246902 239912 246954 239964
rect 247178 239912 247230 239964
rect 247362 239912 247414 239964
rect 247546 239912 247598 239964
rect 248006 239912 248058 239964
rect 248098 239912 248150 239964
rect 248466 239912 248518 239964
rect 248650 239912 248702 239964
rect 245982 239844 246034 239896
rect 246212 239776 246264 239828
rect 246028 239640 246080 239692
rect 246212 239572 246264 239624
rect 245200 239504 245252 239556
rect 245936 239436 245988 239488
rect 244648 239368 244700 239420
rect 246488 239572 246540 239624
rect 246672 239572 246724 239624
rect 247040 239640 247092 239692
rect 247868 239708 247920 239760
rect 247960 239708 248012 239760
rect 247408 239572 247460 239624
rect 248052 239572 248104 239624
rect 246856 239504 246908 239556
rect 248328 239436 248380 239488
rect 248604 239708 248656 239760
rect 248926 239912 248978 239964
rect 249018 239912 249070 239964
rect 248972 239776 249024 239828
rect 248880 239572 248932 239624
rect 267464 241272 267516 241324
rect 268108 241272 268160 241324
rect 267648 241204 267700 241256
rect 268200 241204 268252 241256
rect 267740 241136 267792 241188
rect 249294 239912 249346 239964
rect 249386 239912 249438 239964
rect 250122 239912 250174 239964
rect 250306 239912 250358 239964
rect 250398 239912 250450 239964
rect 250582 239912 250634 239964
rect 250674 239912 250726 239964
rect 249662 239844 249714 239896
rect 249248 239504 249300 239556
rect 249800 239572 249852 239624
rect 250352 239640 250404 239692
rect 250260 239572 250312 239624
rect 250628 239776 250680 239828
rect 267556 241068 267608 241120
rect 267648 241068 267700 241120
rect 251134 239912 251186 239964
rect 251226 239912 251278 239964
rect 251778 239912 251830 239964
rect 252238 239912 252290 239964
rect 252330 239912 252382 239964
rect 250950 239844 251002 239896
rect 250904 239708 250956 239760
rect 251318 239844 251370 239896
rect 251594 239844 251646 239896
rect 251686 239844 251738 239896
rect 251180 239708 251232 239760
rect 252054 239844 252106 239896
rect 252146 239844 252198 239896
rect 250536 239572 250588 239624
rect 250720 239572 250772 239624
rect 251088 239572 251140 239624
rect 251364 239572 251416 239624
rect 251640 239640 251692 239692
rect 252008 239708 252060 239760
rect 313924 241000 313976 241052
rect 267740 240932 267792 240984
rect 309048 240932 309100 240984
rect 268108 240864 268160 240916
rect 300400 240864 300452 240916
rect 267740 240796 267792 240848
rect 316224 240796 316276 240848
rect 329104 240728 329156 240780
rect 267556 240660 267608 240712
rect 267740 240592 267792 240644
rect 252606 239912 252658 239964
rect 252698 239912 252750 239964
rect 253250 239912 253302 239964
rect 252422 239776 252474 239828
rect 252284 239640 252336 239692
rect 252376 239640 252428 239692
rect 252790 239844 252842 239896
rect 252744 239708 252796 239760
rect 252652 239640 252704 239692
rect 252192 239572 252244 239624
rect 253066 239844 253118 239896
rect 253112 239708 253164 239760
rect 253526 239912 253578 239964
rect 253618 239912 253670 239964
rect 253802 239912 253854 239964
rect 253894 239912 253946 239964
rect 253112 239572 253164 239624
rect 253388 239640 253440 239692
rect 253664 239640 253716 239692
rect 253756 239640 253808 239692
rect 254078 239844 254130 239896
rect 254354 239912 254406 239964
rect 254814 239912 254866 239964
rect 254906 239912 254958 239964
rect 255274 239912 255326 239964
rect 255458 239912 255510 239964
rect 254124 239640 254176 239692
rect 254216 239640 254268 239692
rect 253480 239572 253532 239624
rect 254446 239844 254498 239896
rect 254630 239844 254682 239896
rect 254860 239776 254912 239828
rect 254492 239640 254544 239692
rect 254768 239572 254820 239624
rect 251272 239504 251324 239556
rect 251548 239504 251600 239556
rect 251916 239504 251968 239556
rect 255044 239572 255096 239624
rect 255366 239844 255418 239896
rect 255550 239844 255602 239896
rect 255320 239504 255372 239556
rect 248880 239436 248932 239488
rect 249064 239436 249116 239488
rect 253204 239436 253256 239488
rect 255826 239912 255878 239964
rect 255918 239912 255970 239964
rect 256010 239912 256062 239964
rect 256102 239912 256154 239964
rect 255734 239844 255786 239896
rect 255504 239572 255556 239624
rect 255596 239572 255648 239624
rect 255964 239640 256016 239692
rect 256056 239572 256108 239624
rect 256378 239912 256430 239964
rect 256332 239572 256384 239624
rect 256562 239844 256614 239896
rect 268292 240524 268344 240576
rect 268752 240388 268804 240440
rect 267740 240320 267792 240372
rect 269304 240320 269356 240372
rect 256930 239912 256982 239964
rect 257022 239912 257074 239964
rect 257114 239844 257166 239896
rect 256976 239776 257028 239828
rect 257068 239708 257120 239760
rect 256516 239504 256568 239556
rect 256700 239436 256752 239488
rect 256976 239572 257028 239624
rect 257758 239912 257810 239964
rect 257850 239912 257902 239964
rect 257390 239844 257442 239896
rect 258034 239844 258086 239896
rect 258126 239844 258178 239896
rect 257804 239708 257856 239760
rect 257896 239640 257948 239692
rect 257988 239640 258040 239692
rect 257436 239572 257488 239624
rect 258678 239912 258730 239964
rect 258862 239912 258914 239964
rect 258310 239844 258362 239896
rect 258402 239844 258454 239896
rect 258356 239708 258408 239760
rect 258632 239640 258684 239692
rect 258540 239572 258592 239624
rect 258448 239504 258500 239556
rect 259414 239912 259466 239964
rect 259690 239912 259742 239964
rect 259874 239912 259926 239964
rect 259782 239844 259834 239896
rect 259368 239640 259420 239692
rect 259736 239640 259788 239692
rect 259092 239572 259144 239624
rect 259184 239572 259236 239624
rect 259966 239844 260018 239896
rect 259828 239572 259880 239624
rect 269212 240252 269264 240304
rect 268016 240184 268068 240236
rect 309784 240184 309836 240236
rect 260242 239912 260294 239964
rect 260334 239844 260386 239896
rect 260288 239640 260340 239692
rect 260380 239572 260432 239624
rect 259460 239504 259512 239556
rect 259920 239504 259972 239556
rect 260104 239504 260156 239556
rect 260610 239912 260662 239964
rect 260794 239912 260846 239964
rect 261070 239912 261122 239964
rect 261162 239912 261214 239964
rect 261254 239912 261306 239964
rect 261346 239912 261398 239964
rect 261438 239912 261490 239964
rect 261622 239912 261674 239964
rect 261714 239912 261766 239964
rect 261990 239912 262042 239964
rect 262358 239912 262410 239964
rect 262542 239912 262594 239964
rect 262634 239912 262686 239964
rect 263094 239912 263146 239964
rect 263186 239912 263238 239964
rect 263462 239912 263514 239964
rect 260656 239708 260708 239760
rect 260886 239844 260938 239896
rect 260978 239844 261030 239896
rect 261116 239776 261168 239828
rect 260840 239708 260892 239760
rect 261024 239708 261076 239760
rect 260932 239640 260984 239692
rect 257620 239436 257672 239488
rect 258816 239436 258868 239488
rect 260564 239436 260616 239488
rect 261346 239708 261398 239760
rect 261392 239504 261444 239556
rect 261576 239504 261628 239556
rect 261806 239844 261858 239896
rect 262266 239844 262318 239896
rect 262588 239776 262640 239828
rect 262404 239708 262456 239760
rect 261852 239640 261904 239692
rect 261944 239640 261996 239692
rect 262312 239640 262364 239692
rect 262910 239844 262962 239896
rect 263002 239844 263054 239896
rect 262496 239572 262548 239624
rect 262680 239572 262732 239624
rect 262772 239504 262824 239556
rect 263554 239844 263606 239896
rect 263140 239776 263192 239828
rect 263232 239776 263284 239828
rect 263508 239640 263560 239692
rect 263922 239912 263974 239964
rect 264106 239912 264158 239964
rect 264198 239912 264250 239964
rect 264290 239912 264342 239964
rect 263968 239708 264020 239760
rect 264060 239708 264112 239760
rect 264152 239708 264204 239760
rect 263876 239572 263928 239624
rect 263324 239504 263376 239556
rect 264658 239912 264710 239964
rect 264750 239912 264802 239964
rect 265026 239912 265078 239964
rect 265118 239912 265170 239964
rect 265302 239912 265354 239964
rect 265394 239912 265446 239964
rect 265670 239912 265722 239964
rect 265762 239912 265814 239964
rect 264566 239776 264618 239828
rect 264704 239776 264756 239828
rect 265072 239776 265124 239828
rect 264980 239708 265032 239760
rect 265256 239708 265308 239760
rect 265716 239776 265768 239828
rect 265348 239640 265400 239692
rect 264796 239572 264848 239624
rect 267924 240048 267976 240100
rect 268292 240116 268344 240168
rect 331588 240116 331640 240168
rect 269028 240048 269080 240100
rect 306748 240048 306800 240100
rect 314936 240048 314988 240100
rect 330392 240048 330444 240100
rect 331128 240048 331180 240100
rect 266130 239912 266182 239964
rect 266222 239912 266274 239964
rect 266406 239912 266458 239964
rect 266498 239912 266550 239964
rect 266314 239844 266366 239896
rect 266084 239572 266136 239624
rect 266452 239708 266504 239760
rect 267556 239980 267608 240032
rect 266866 239912 266918 239964
rect 267050 239912 267102 239964
rect 267142 239912 267194 239964
rect 267464 239912 267516 239964
rect 267832 239912 267884 239964
rect 266774 239844 266826 239896
rect 266820 239708 266872 239760
rect 267004 239708 267056 239760
rect 292948 239980 293000 240032
rect 267556 239776 267608 239828
rect 267648 239708 267700 239760
rect 269396 239640 269448 239692
rect 266360 239572 266412 239624
rect 266636 239572 266688 239624
rect 291752 239776 291804 239828
rect 264980 239504 265032 239556
rect 265348 239504 265400 239556
rect 267372 239504 267424 239556
rect 268200 239504 268252 239556
rect 269488 239504 269540 239556
rect 286784 239504 286836 239556
rect 321100 239436 321152 239488
rect 249616 239368 249668 239420
rect 251640 239368 251692 239420
rect 238116 239300 238168 239352
rect 247960 239300 248012 239352
rect 249156 239300 249208 239352
rect 252560 239300 252612 239352
rect 253388 239300 253440 239352
rect 257344 239368 257396 239420
rect 263508 239368 263560 239420
rect 266268 239368 266320 239420
rect 297180 239368 297232 239420
rect 265348 239300 265400 239352
rect 266544 239300 266596 239352
rect 267372 239300 267424 239352
rect 268200 239300 268252 239352
rect 274456 239300 274508 239352
rect 200120 239232 200172 239284
rect 216036 239232 216088 239284
rect 216588 239232 216640 239284
rect 220268 239232 220320 239284
rect 232044 239232 232096 239284
rect 232136 239232 232188 239284
rect 232780 239232 232832 239284
rect 233424 239232 233476 239284
rect 195980 239164 196032 239216
rect 219072 239164 219124 239216
rect 234988 239164 235040 239216
rect 247316 239232 247368 239284
rect 248144 239232 248196 239284
rect 248236 239232 248288 239284
rect 249340 239232 249392 239284
rect 250444 239232 250496 239284
rect 252100 239232 252152 239284
rect 255044 239232 255096 239284
rect 314200 239232 314252 239284
rect 252560 239164 252612 239216
rect 256424 239164 256476 239216
rect 294236 239164 294288 239216
rect 306656 239164 306708 239216
rect 321560 239164 321612 239216
rect 216128 239096 216180 239148
rect 215576 239028 215628 239080
rect 228364 239028 228416 239080
rect 229744 239096 229796 239148
rect 231860 239096 231912 239148
rect 232044 239096 232096 239148
rect 237748 239096 237800 239148
rect 237932 239096 237984 239148
rect 238392 239096 238444 239148
rect 253940 239096 253992 239148
rect 237656 239028 237708 239080
rect 248880 239028 248932 239080
rect 250720 239028 250772 239080
rect 254216 239028 254268 239080
rect 216588 238960 216640 239012
rect 221648 238892 221700 238944
rect 225604 238892 225656 238944
rect 238024 238960 238076 239012
rect 250168 238960 250220 239012
rect 250444 238960 250496 239012
rect 257712 239028 257764 239080
rect 260472 239028 260524 239080
rect 261852 239096 261904 239148
rect 322572 239096 322624 239148
rect 314384 239028 314436 239080
rect 232136 238892 232188 238944
rect 239588 238892 239640 238944
rect 217784 238824 217836 238876
rect 226340 238824 226392 238876
rect 227168 238824 227220 238876
rect 233700 238824 233752 238876
rect 234620 238824 234672 238876
rect 256424 238892 256476 238944
rect 313464 238960 313516 239012
rect 247408 238824 247460 238876
rect 248052 238824 248104 238876
rect 220360 238756 220412 238808
rect 235172 238756 235224 238808
rect 236460 238756 236512 238808
rect 236644 238756 236696 238808
rect 237932 238756 237984 238808
rect 238668 238756 238720 238808
rect 239588 238756 239640 238808
rect 251640 238824 251692 238876
rect 253388 238824 253440 238876
rect 258816 238824 258868 238876
rect 267556 238892 267608 238944
rect 267924 238892 267976 238944
rect 331128 238892 331180 238944
rect 260472 238824 260524 238876
rect 268200 238824 268252 238876
rect 250352 238756 250404 238808
rect 250904 238756 250956 238808
rect 251272 238756 251324 238808
rect 254492 238756 254544 238808
rect 206376 238688 206428 238740
rect 212080 238688 212132 238740
rect 225696 238688 225748 238740
rect 225972 238688 226024 238740
rect 233148 238688 233200 238740
rect 234252 238688 234304 238740
rect 239220 238688 239272 238740
rect 240876 238688 240928 238740
rect 241428 238688 241480 238740
rect 241980 238688 242032 238740
rect 242256 238688 242308 238740
rect 244556 238688 244608 238740
rect 244740 238688 244792 238740
rect 245016 238688 245068 238740
rect 245200 238688 245252 238740
rect 246028 238688 246080 238740
rect 246488 238688 246540 238740
rect 246580 238688 246632 238740
rect 246764 238688 246816 238740
rect 247408 238688 247460 238740
rect 247592 238688 247644 238740
rect 250628 238688 250680 238740
rect 250812 238688 250864 238740
rect 251732 238688 251784 238740
rect 251916 238688 251968 238740
rect 259184 238756 259236 238808
rect 260288 238756 260340 238808
rect 267924 238756 267976 238808
rect 221556 238620 221608 238672
rect 242992 238620 243044 238672
rect 250444 238620 250496 238672
rect 250904 238620 250956 238672
rect 253204 238620 253256 238672
rect 263508 238688 263560 238740
rect 266268 238688 266320 238740
rect 267280 238688 267332 238740
rect 267740 238688 267792 238740
rect 260840 238620 260892 238672
rect 332968 238824 333020 238876
rect 221372 238552 221424 238604
rect 226616 238552 226668 238604
rect 229008 238552 229060 238604
rect 239496 238552 239548 238604
rect 245752 238552 245804 238604
rect 249064 238552 249116 238604
rect 249616 238552 249668 238604
rect 253388 238552 253440 238604
rect 264244 238552 264296 238604
rect 264520 238552 264572 238604
rect 212264 238484 212316 238536
rect 225236 238484 225288 238536
rect 226248 238484 226300 238536
rect 227076 238484 227128 238536
rect 231860 238484 231912 238536
rect 232044 238484 232096 238536
rect 232872 238484 232924 238536
rect 233148 238484 233200 238536
rect 238484 238484 238536 238536
rect 241520 238484 241572 238536
rect 246396 238484 246448 238536
rect 248512 238484 248564 238536
rect 250444 238484 250496 238536
rect 256240 238484 256292 238536
rect 259000 238484 259052 238536
rect 261668 238484 261720 238536
rect 296628 238756 296680 238808
rect 489920 238756 489972 238808
rect 221188 238416 221240 238468
rect 224316 238416 224368 238468
rect 224592 238416 224644 238468
rect 229468 238416 229520 238468
rect 229928 238416 229980 238468
rect 270316 238416 270368 238468
rect 221740 238348 221792 238400
rect 230388 238348 230440 238400
rect 230480 238348 230532 238400
rect 270224 238348 270276 238400
rect 220268 238280 220320 238332
rect 228916 238280 228968 238332
rect 231768 238280 231820 238332
rect 270408 238280 270460 238332
rect 214564 238212 214616 238264
rect 221188 238212 221240 238264
rect 221280 238212 221332 238264
rect 225972 238212 226024 238264
rect 226616 238212 226668 238264
rect 227536 238212 227588 238264
rect 230940 238212 230992 238264
rect 269672 238212 269724 238264
rect 213368 238144 213420 238196
rect 223948 238144 224000 238196
rect 227260 238144 227312 238196
rect 232596 238144 232648 238196
rect 232780 238144 232832 238196
rect 269580 238144 269632 238196
rect 194600 238076 194652 238128
rect 85580 238008 85632 238060
rect 214656 238008 214708 238060
rect 221648 238076 221700 238128
rect 227628 238076 227680 238128
rect 231860 238076 231912 238128
rect 235816 238076 235868 238128
rect 238116 238076 238168 238128
rect 239220 238076 239272 238128
rect 243820 238076 243872 238128
rect 244832 238076 244884 238128
rect 245752 238076 245804 238128
rect 246304 238076 246356 238128
rect 255228 238076 255280 238128
rect 260472 238076 260524 238128
rect 262956 238076 263008 238128
rect 264888 238076 264940 238128
rect 217416 238008 217468 238060
rect 230204 238008 230256 238060
rect 230480 238008 230532 238060
rect 231032 238008 231084 238060
rect 236184 238008 236236 238060
rect 237196 238008 237248 238060
rect 240232 238008 240284 238060
rect 240416 238008 240468 238060
rect 242808 238008 242860 238060
rect 246948 238008 247000 238060
rect 249708 238008 249760 238060
rect 250168 238008 250220 238060
rect 255964 238008 256016 238060
rect 256424 238008 256476 238060
rect 256516 238008 256568 238060
rect 257068 238008 257120 238060
rect 267832 238008 267884 238060
rect 302700 238076 302752 238128
rect 268660 238008 268712 238060
rect 308404 238008 308456 238060
rect 216404 237940 216456 237992
rect 237564 237940 237616 237992
rect 253940 237940 253992 237992
rect 257344 237940 257396 237992
rect 214656 237872 214708 237924
rect 229100 237872 229152 237924
rect 231032 237872 231084 237924
rect 231768 237872 231820 237924
rect 234712 237872 234764 237924
rect 242164 237872 242216 237924
rect 245568 237872 245620 237924
rect 257068 237872 257120 237924
rect 260564 237872 260616 237924
rect 270132 237872 270184 237924
rect 221464 237804 221516 237856
rect 242808 237804 242860 237856
rect 252560 237804 252612 237856
rect 258724 237804 258776 237856
rect 221096 237736 221148 237788
rect 222752 237736 222804 237788
rect 224408 237736 224460 237788
rect 224868 237736 224920 237788
rect 226064 237736 226116 237788
rect 226984 237736 227036 237788
rect 246120 237736 246172 237788
rect 251916 237736 251968 237788
rect 256884 237736 256936 237788
rect 315488 237804 315540 237856
rect 261484 237736 261536 237788
rect 269120 237736 269172 237788
rect 220176 237668 220228 237720
rect 228732 237668 228784 237720
rect 218980 237600 219032 237652
rect 223304 237600 223356 237652
rect 224960 237600 225012 237652
rect 225144 237600 225196 237652
rect 226156 237600 226208 237652
rect 271052 237668 271104 237720
rect 243084 237600 243136 237652
rect 249708 237600 249760 237652
rect 254768 237600 254820 237652
rect 256884 237600 256936 237652
rect 220820 237532 220872 237584
rect 224132 237532 224184 237584
rect 224868 237532 224920 237584
rect 225420 237532 225472 237584
rect 231400 237532 231452 237584
rect 290648 237532 290700 237584
rect 213184 237464 213236 237516
rect 235724 237464 235776 237516
rect 236828 237464 236880 237516
rect 249064 237464 249116 237516
rect 254768 237464 254820 237516
rect 256056 237464 256108 237516
rect 315396 237464 315448 237516
rect 157340 237396 157392 237448
rect 233700 237396 233752 237448
rect 267740 237396 267792 237448
rect 336004 237396 336056 237448
rect 212356 237328 212408 237380
rect 215300 237328 215352 237380
rect 216588 237328 216640 237380
rect 222568 237328 222620 237380
rect 223120 237328 223172 237380
rect 234620 237328 234672 237380
rect 239496 237328 239548 237380
rect 249984 237328 250036 237380
rect 250720 237328 250772 237380
rect 265072 237328 265124 237380
rect 333980 237328 334032 237380
rect 334440 237328 334492 237380
rect 221004 237260 221056 237312
rect 223028 237260 223080 237312
rect 224776 237260 224828 237312
rect 225144 237260 225196 237312
rect 226248 237260 226300 237312
rect 232412 237260 232464 237312
rect 246948 237260 247000 237312
rect 222660 237192 222712 237244
rect 223396 237192 223448 237244
rect 265624 237260 265676 237312
rect 330208 237260 330260 237312
rect 260380 237192 260432 237244
rect 260748 237192 260800 237244
rect 321284 237192 321336 237244
rect 215116 237124 215168 237176
rect 230020 237124 230072 237176
rect 237564 237124 237616 237176
rect 240140 237124 240192 237176
rect 298100 237124 298152 237176
rect 214932 237056 214984 237108
rect 225420 237056 225472 237108
rect 249340 237056 249392 237108
rect 307576 237056 307628 237108
rect 215024 236988 215076 237040
rect 224960 236988 225012 237040
rect 250996 236988 251048 237040
rect 259000 236988 259052 237040
rect 259828 236988 259880 237040
rect 319444 236988 319496 237040
rect 215852 236920 215904 236972
rect 224592 236920 224644 236972
rect 232320 236920 232372 236972
rect 281264 236920 281316 236972
rect 217876 236852 217928 236904
rect 225972 236852 226024 236904
rect 228732 236852 228784 236904
rect 231124 236852 231176 236904
rect 239220 236852 239272 236904
rect 275652 236852 275704 236904
rect 331128 236852 331180 236904
rect 487160 236852 487212 236904
rect 191840 236716 191892 236768
rect 216312 236784 216364 236836
rect 236000 236784 236052 236836
rect 243084 236784 243136 236836
rect 244188 236784 244240 236836
rect 244924 236784 244976 236836
rect 279424 236784 279476 236836
rect 332968 236784 333020 236836
rect 494060 236784 494112 236836
rect 231124 236716 231176 236768
rect 231400 236716 231452 236768
rect 243452 236716 243504 236768
rect 246948 236716 247000 236768
rect 278688 236716 278740 236768
rect 330208 236716 330260 236768
rect 529204 236716 529256 236768
rect 126980 236648 127032 236700
rect 220544 236648 220596 236700
rect 226248 236648 226300 236700
rect 231860 236648 231912 236700
rect 232136 236648 232188 236700
rect 237472 236648 237524 236700
rect 238116 236648 238168 236700
rect 241336 236648 241388 236700
rect 244280 236648 244332 236700
rect 245936 236648 245988 236700
rect 210976 236580 211028 236632
rect 226892 236580 226944 236632
rect 256700 236580 256752 236632
rect 265256 236580 265308 236632
rect 266452 236648 266504 236700
rect 267188 236648 267240 236700
rect 271144 236648 271196 236700
rect 271696 236648 271748 236700
rect 307576 236648 307628 236700
rect 332600 236648 332652 236700
rect 333980 236648 334032 236700
rect 540244 236648 540296 236700
rect 214748 236512 214800 236564
rect 220912 236512 220964 236564
rect 223672 236512 223724 236564
rect 246764 236512 246816 236564
rect 255964 236512 256016 236564
rect 256792 236512 256844 236564
rect 257988 236512 258040 236564
rect 213552 236444 213604 236496
rect 229376 236444 229428 236496
rect 253664 236444 253716 236496
rect 261668 236444 261720 236496
rect 253020 236376 253072 236428
rect 256792 236376 256844 236428
rect 258724 236376 258776 236428
rect 269764 236376 269816 236428
rect 213920 236308 213972 236360
rect 214472 236308 214524 236360
rect 224224 236308 224276 236360
rect 224500 236308 224552 236360
rect 235172 236308 235224 236360
rect 282736 236308 282788 236360
rect 220728 236240 220780 236292
rect 223580 236240 223632 236292
rect 228364 236240 228416 236292
rect 235448 236240 235500 236292
rect 278136 236240 278188 236292
rect 244832 236172 244884 236224
rect 258724 236172 258776 236224
rect 249892 236104 249944 236156
rect 250352 236104 250404 236156
rect 252376 236104 252428 236156
rect 260748 236104 260800 236156
rect 266176 236036 266228 236088
rect 269028 236036 269080 236088
rect 214656 235968 214708 236020
rect 215116 235968 215168 236020
rect 252928 235968 252980 236020
rect 256148 235968 256200 236020
rect 263784 235968 263836 236020
rect 264152 235968 264204 236020
rect 212448 235900 212500 235952
rect 229192 235900 229244 235952
rect 251548 235900 251600 235952
rect 253204 235900 253256 235952
rect 253940 235900 253992 235952
rect 337016 235900 337068 235952
rect 338028 235900 338080 235952
rect 256516 235832 256568 235884
rect 263140 235832 263192 235884
rect 265440 235832 265492 235884
rect 331496 235832 331548 235884
rect 220820 235764 220872 235816
rect 237656 235764 237708 235816
rect 250904 235764 250956 235816
rect 267740 235764 267792 235816
rect 218612 235696 218664 235748
rect 230480 235696 230532 235748
rect 209780 235628 209832 235680
rect 238760 235628 238812 235680
rect 294604 235696 294656 235748
rect 246580 235628 246632 235680
rect 298744 235628 298796 235680
rect 211160 235560 211212 235612
rect 238944 235560 238996 235612
rect 286876 235560 286928 235612
rect 175924 235492 175976 235544
rect 226156 235492 226208 235544
rect 236000 235492 236052 235544
rect 236184 235492 236236 235544
rect 282644 235492 282696 235544
rect 115204 235424 115256 235476
rect 230572 235424 230624 235476
rect 235724 235424 235776 235476
rect 275284 235424 275336 235476
rect 95884 235356 95936 235408
rect 212448 235356 212500 235408
rect 213276 235356 213328 235408
rect 237380 235356 237432 235408
rect 106280 235288 106332 235340
rect 230848 235288 230900 235340
rect 232504 235288 232556 235340
rect 232872 235288 232924 235340
rect 60740 235220 60792 235272
rect 226800 235220 226852 235272
rect 228732 235220 228784 235272
rect 237564 235220 237616 235272
rect 224040 235152 224092 235204
rect 224684 235152 224736 235204
rect 244372 235356 244424 235408
rect 281540 235356 281592 235408
rect 282828 235356 282880 235408
rect 338028 235356 338080 235408
rect 369860 235356 369912 235408
rect 243268 235288 243320 235340
rect 262956 235288 263008 235340
rect 244004 235220 244056 235272
rect 266360 235220 266412 235272
rect 266820 235220 266872 235272
rect 331588 235288 331640 235340
rect 498292 235288 498344 235340
rect 275928 235220 275980 235272
rect 294696 235220 294748 235272
rect 331496 235220 331548 235272
rect 550640 235220 550692 235272
rect 258172 235152 258224 235204
rect 258448 235152 258500 235204
rect 262220 235152 262272 235204
rect 262864 235152 262916 235204
rect 262956 235152 263008 235204
rect 267832 235152 267884 235204
rect 272984 235084 273036 235136
rect 237656 235016 237708 235068
rect 239680 235016 239732 235068
rect 296260 235016 296312 235068
rect 235816 234948 235868 235000
rect 279884 234948 279936 235000
rect 251180 234880 251232 234932
rect 253940 234880 253992 234932
rect 257436 234880 257488 234932
rect 260196 234880 260248 234932
rect 262312 234880 262364 234932
rect 263416 234880 263468 234932
rect 236092 234608 236144 234660
rect 236460 234608 236512 234660
rect 331496 234608 331548 234660
rect 331956 234608 332008 234660
rect 512644 234608 512696 234660
rect 234252 234540 234304 234592
rect 294144 234540 294196 234592
rect 234344 234472 234396 234524
rect 292764 234472 292816 234524
rect 234804 234404 234856 234456
rect 235356 234404 235408 234456
rect 236552 234404 236604 234456
rect 239404 234404 239456 234456
rect 299204 234404 299256 234456
rect 247500 234336 247552 234388
rect 306656 234336 306708 234388
rect 233976 234268 234028 234320
rect 292856 234268 292908 234320
rect 231768 234200 231820 234252
rect 240508 234200 240560 234252
rect 298836 234200 298888 234252
rect 254032 234132 254084 234184
rect 311808 234132 311860 234184
rect 229560 234064 229612 234116
rect 230204 234064 230256 234116
rect 235724 234064 235776 234116
rect 236736 234064 236788 234116
rect 293224 234064 293276 234116
rect 218060 233996 218112 234048
rect 236552 233996 236604 234048
rect 241520 233996 241572 234048
rect 242256 233996 242308 234048
rect 243176 233996 243228 234048
rect 244188 233996 244240 234048
rect 247132 233996 247184 234048
rect 228272 233928 228324 233980
rect 228824 233928 228876 233980
rect 232964 233928 233016 233980
rect 282460 233928 282512 233980
rect 300952 233928 301004 233980
rect 313924 233928 313976 233980
rect 143540 233860 143592 233912
rect 233608 233860 233660 233912
rect 234344 233860 234396 233912
rect 237564 233860 237616 233912
rect 238392 233860 238444 233912
rect 241520 233860 241572 233912
rect 241888 233860 241940 233912
rect 245384 233860 245436 233912
rect 277216 233860 277268 233912
rect 278044 233860 278096 233912
rect 405740 233860 405792 233912
rect 227904 233792 227956 233844
rect 228548 233792 228600 233844
rect 229744 233792 229796 233844
rect 230388 233792 230440 233844
rect 245108 233792 245160 233844
rect 274548 233792 274600 233844
rect 275284 233792 275336 233844
rect 243544 233656 243596 233708
rect 271236 233724 271288 233776
rect 226616 233588 226668 233640
rect 227352 233588 227404 233640
rect 227996 233588 228048 233640
rect 228456 233588 228508 233640
rect 233608 233452 233660 233504
rect 234160 233452 234212 233504
rect 227812 233384 227864 233436
rect 249708 233384 249760 233436
rect 272616 233656 272668 233708
rect 256792 233316 256844 233368
rect 257436 233316 257488 233368
rect 234068 233180 234120 233232
rect 294512 233180 294564 233232
rect 345664 233180 345716 233232
rect 579988 233180 580040 233232
rect 241980 233112 242032 233164
rect 242716 233112 242768 233164
rect 249800 233112 249852 233164
rect 310152 233112 310204 233164
rect 310428 233112 310480 233164
rect 227812 233044 227864 233096
rect 247408 233044 247460 233096
rect 303712 233044 303764 233096
rect 242164 232976 242216 233028
rect 251180 232976 251232 233028
rect 254492 232976 254544 233028
rect 309508 232976 309560 233028
rect 239588 232908 239640 232960
rect 239864 232908 239916 232960
rect 292028 232908 292080 232960
rect 191104 232840 191156 232892
rect 236000 232840 236052 232892
rect 245660 232840 245712 232892
rect 295984 232840 296036 232892
rect 183560 232772 183612 232824
rect 235724 232772 235776 232824
rect 238760 232772 238812 232824
rect 240968 232772 241020 232824
rect 279608 232772 279660 232824
rect 132500 232704 132552 232756
rect 220084 232704 220136 232756
rect 238484 232704 238536 232756
rect 240692 232704 240744 232756
rect 241244 232704 241296 232756
rect 241428 232704 241480 232756
rect 272800 232704 272852 232756
rect 111800 232636 111852 232688
rect 231308 232636 231360 232688
rect 246396 232636 246448 232688
rect 276940 232636 276992 232688
rect 89720 232568 89772 232620
rect 213552 232568 213604 232620
rect 243912 232568 243964 232620
rect 271880 232568 271932 232620
rect 62764 232500 62816 232552
rect 210976 232500 211028 232552
rect 242532 232500 242584 232552
rect 251088 232500 251140 232552
rect 300308 232500 300360 232552
rect 310428 232500 310480 232552
rect 356060 232500 356112 232552
rect 251180 232432 251232 232484
rect 252376 232432 252428 232484
rect 279792 232432 279844 232484
rect 242716 232364 242768 232416
rect 268384 232364 268436 232416
rect 242256 232296 242308 232348
rect 248328 232296 248380 232348
rect 272892 232296 272944 232348
rect 266084 232228 266136 232280
rect 269396 232228 269448 232280
rect 227720 232160 227772 232212
rect 228732 232160 228784 232212
rect 252192 232160 252244 232212
rect 255320 232160 255372 232212
rect 271880 232160 271932 232212
rect 273168 232160 273220 232212
rect 273904 232160 273956 232212
rect 240324 231888 240376 231940
rect 240876 231888 240928 231940
rect 245660 231820 245712 231872
rect 246396 231820 246448 231872
rect 303712 231820 303764 231872
rect 324596 231820 324648 231872
rect 241796 231752 241848 231804
rect 243636 231752 243688 231804
rect 250168 231752 250220 231804
rect 335820 231752 335872 231804
rect 336648 231752 336700 231804
rect 248880 231684 248932 231736
rect 328828 231684 328880 231736
rect 329196 231684 329248 231736
rect 251364 231616 251416 231668
rect 311256 231616 311308 231668
rect 248052 231548 248104 231600
rect 306564 231548 306616 231600
rect 307576 231548 307628 231600
rect 225236 231480 225288 231532
rect 226064 231480 226116 231532
rect 236552 231480 236604 231532
rect 239312 231480 239364 231532
rect 299020 231480 299072 231532
rect 240416 231412 240468 231464
rect 240784 231412 240836 231464
rect 299848 231412 299900 231464
rect 265256 231344 265308 231396
rect 233240 231276 233292 231328
rect 240600 231276 240652 231328
rect 282552 231276 282604 231328
rect 244832 231208 244884 231260
rect 284208 231208 284260 231260
rect 236000 231140 236052 231192
rect 240876 231140 240928 231192
rect 279700 231140 279752 231192
rect 74540 231072 74592 231124
rect 228916 231072 228968 231124
rect 257068 231072 257120 231124
rect 296720 231072 296772 231124
rect 298008 231072 298060 231124
rect 307576 231140 307628 231192
rect 320180 231140 320232 231192
rect 336648 231140 336700 231192
rect 351184 231140 351236 231192
rect 315764 231072 315816 231124
rect 421564 231072 421616 231124
rect 275560 231004 275612 231056
rect 233884 230936 233936 230988
rect 234068 230936 234120 230988
rect 237656 230936 237708 230988
rect 238300 230936 238352 230988
rect 239956 230936 240008 230988
rect 274364 230936 274416 230988
rect 239404 230868 239456 230920
rect 271604 230868 271656 230920
rect 233700 230732 233752 230784
rect 234528 230732 234580 230784
rect 264060 230732 264112 230784
rect 264888 230732 264940 230784
rect 226432 230596 226484 230648
rect 227260 230596 227312 230648
rect 239496 230460 239548 230512
rect 239956 230460 240008 230512
rect 254308 230460 254360 230512
rect 254768 230460 254820 230512
rect 236736 230392 236788 230444
rect 237288 230392 237340 230444
rect 298008 230392 298060 230444
rect 305368 230392 305420 230444
rect 232688 230324 232740 230376
rect 292672 230324 292724 230376
rect 251456 230256 251508 230308
rect 311256 230256 311308 230308
rect 311624 230256 311676 230308
rect 232872 230188 232924 230240
rect 291660 230188 291712 230240
rect 248420 230120 248472 230172
rect 306104 230120 306156 230172
rect 237288 230052 237340 230104
rect 289268 230052 289320 230104
rect 218152 229984 218204 230036
rect 236552 229984 236604 230036
rect 244464 229984 244516 230036
rect 245200 229984 245252 230036
rect 246120 229984 246172 230036
rect 291844 229984 291896 230036
rect 235540 229916 235592 229968
rect 278320 229916 278372 229968
rect 234988 229848 235040 229900
rect 276848 229848 276900 229900
rect 179420 229780 179472 229832
rect 236368 229780 236420 229832
rect 274180 229780 274232 229832
rect 10324 229712 10376 229764
rect 221924 229712 221976 229764
rect 232596 229712 232648 229764
rect 232964 229712 233016 229764
rect 236644 229712 236696 229764
rect 274272 229712 274324 229764
rect 311256 229712 311308 229764
rect 374092 229712 374144 229764
rect 243084 229644 243136 229696
rect 278780 229644 278832 229696
rect 235908 229576 235960 229628
rect 239128 229508 239180 229560
rect 236276 229440 236328 229492
rect 244372 229372 244424 229424
rect 245292 229372 245344 229424
rect 238024 229304 238076 229356
rect 239128 229304 239180 229356
rect 254124 229440 254176 229492
rect 254584 229440 254636 229492
rect 255780 229440 255832 229492
rect 256516 229440 256568 229492
rect 256700 229440 256752 229492
rect 257712 229440 257764 229492
rect 258264 229440 258316 229492
rect 258908 229440 258960 229492
rect 260840 229440 260892 229492
rect 261392 229440 261444 229492
rect 254032 229372 254084 229424
rect 254860 229372 254912 229424
rect 258080 229372 258132 229424
rect 258632 229372 258684 229424
rect 260932 229372 260984 229424
rect 261576 229372 261628 229424
rect 264428 229576 264480 229628
rect 264704 229576 264756 229628
rect 265532 229576 265584 229628
rect 265992 229576 266044 229628
rect 271420 229440 271472 229492
rect 272708 229372 272760 229424
rect 258172 229304 258224 229356
rect 259276 229304 259328 229356
rect 297088 229440 297140 229492
rect 235080 229168 235132 229220
rect 235908 229168 235960 229220
rect 253940 229168 253992 229220
rect 255136 229168 255188 229220
rect 230848 229100 230900 229152
rect 240048 229100 240100 229152
rect 306104 229100 306156 229152
rect 333980 229100 334032 229152
rect 256884 229032 256936 229084
rect 289360 229032 289412 229084
rect 249248 228964 249300 229016
rect 338580 228964 338632 229016
rect 345020 228964 345072 229016
rect 247684 228896 247736 228948
rect 320548 228896 320600 228948
rect 247040 228828 247092 228880
rect 314936 228828 314988 228880
rect 246856 228760 246908 228812
rect 309416 228760 309468 228812
rect 246028 228692 246080 228744
rect 306472 228692 306524 228744
rect 252836 228624 252888 228676
rect 313096 228624 313148 228676
rect 172520 228556 172572 228608
rect 235080 228556 235132 228608
rect 249156 228556 249208 228608
rect 305644 228556 305696 228608
rect 150440 228488 150492 228540
rect 233884 228488 233936 228540
rect 255964 228488 256016 228540
rect 310520 228488 310572 228540
rect 96620 228420 96672 228472
rect 214656 228420 214708 228472
rect 253296 228420 253348 228472
rect 307944 228420 307996 228472
rect 46940 228352 46992 228404
rect 217876 228352 217928 228404
rect 251916 228352 251968 228404
rect 303620 228352 303672 228404
rect 313096 228352 313148 228404
rect 390652 228352 390704 228404
rect 254676 228284 254728 228336
rect 299572 228284 299624 228336
rect 230756 228080 230808 228132
rect 231308 228080 231360 228132
rect 269856 228216 269908 228268
rect 278780 228216 278832 228268
rect 304080 228216 304132 228268
rect 250076 228148 250128 228200
rect 342260 228148 342312 228200
rect 303620 227944 303672 227996
rect 304264 227944 304316 227996
rect 299572 227740 299624 227792
rect 300216 227740 300268 227792
rect 306472 227740 306524 227792
rect 309140 227740 309192 227792
rect 309416 227740 309468 227792
rect 309876 227740 309928 227792
rect 320548 227740 320600 227792
rect 320824 227740 320876 227792
rect 342260 227740 342312 227792
rect 342904 227740 342956 227792
rect 251732 227672 251784 227724
rect 334164 227672 334216 227724
rect 334532 227672 334584 227724
rect 250444 227604 250496 227656
rect 329932 227604 329984 227656
rect 259184 227536 259236 227588
rect 331312 227536 331364 227588
rect 241336 227468 241388 227520
rect 303988 227468 304040 227520
rect 233056 227400 233108 227452
rect 293132 227400 293184 227452
rect 258540 227332 258592 227384
rect 318524 227332 318576 227384
rect 255320 227264 255372 227316
rect 312728 227264 312780 227316
rect 186320 227196 186372 227248
rect 236644 227196 236696 227248
rect 240324 227196 240376 227248
rect 241336 227196 241388 227248
rect 246764 227196 246816 227248
rect 303252 227196 303304 227248
rect 123484 227128 123536 227180
rect 226524 227128 226576 227180
rect 247316 227128 247368 227180
rect 302056 227128 302108 227180
rect 122104 227060 122156 227112
rect 231032 227060 231084 227112
rect 250812 227060 250864 227112
rect 250996 227060 251048 227112
rect 260656 227060 260708 227112
rect 312912 227060 312964 227112
rect 334164 227060 334216 227112
rect 376024 227060 376076 227112
rect 7656 226992 7708 227044
rect 222936 226992 222988 227044
rect 234160 226992 234212 227044
rect 244556 226992 244608 227044
rect 283012 226992 283064 227044
rect 318524 226992 318576 227044
rect 458180 226992 458232 227044
rect 271328 226924 271380 226976
rect 241060 226856 241112 226908
rect 276756 226856 276808 226908
rect 241704 226788 241756 226840
rect 247040 226788 247092 226840
rect 274088 226788 274140 226840
rect 233700 226652 233752 226704
rect 234160 226652 234212 226704
rect 283012 226380 283064 226432
rect 283748 226380 283800 226432
rect 240140 226312 240192 226364
rect 241060 226312 241112 226364
rect 302056 226312 302108 226364
rect 319444 226312 319496 226364
rect 329932 226312 329984 226364
rect 330576 226312 330628 226364
rect 331312 226312 331364 226364
rect 331956 226312 332008 226364
rect 260196 226244 260248 226296
rect 349252 226244 349304 226296
rect 258448 226176 258500 226228
rect 335544 226176 335596 226228
rect 336096 226176 336148 226228
rect 252744 226108 252796 226160
rect 312820 226108 312872 226160
rect 261208 226040 261260 226092
rect 321192 226040 321244 226092
rect 254216 225972 254268 226024
rect 314016 225972 314068 226024
rect 256976 225904 257028 225956
rect 317144 225904 317196 225956
rect 317328 225904 317380 225956
rect 248604 225836 248656 225888
rect 305276 225836 305328 225888
rect 256148 225768 256200 225820
rect 312544 225768 312596 225820
rect 229376 225700 229428 225752
rect 230020 225700 230072 225752
rect 240048 225700 240100 225752
rect 296168 225700 296220 225752
rect 146300 225632 146352 225684
rect 233976 225632 234028 225684
rect 309784 225632 309836 225684
rect 385684 225632 385736 225684
rect 136640 225564 136692 225616
rect 233056 225564 233108 225616
rect 260380 225564 260432 225616
rect 314844 225564 314896 225616
rect 317328 225564 317380 225616
rect 443644 225564 443696 225616
rect 264336 225496 264388 225548
rect 317972 225496 318024 225548
rect 318708 225496 318760 225548
rect 243544 225428 243596 225480
rect 273260 225428 273312 225480
rect 230020 225360 230072 225412
rect 275836 225360 275888 225412
rect 261668 225292 261720 225344
rect 314292 225292 314344 225344
rect 273260 224952 273312 225004
rect 273996 224952 274048 225004
rect 305276 224952 305328 225004
rect 338120 224952 338172 225004
rect 349252 224952 349304 225004
rect 349804 224952 349856 225004
rect 254768 224884 254820 224936
rect 332784 224884 332836 224936
rect 333060 224884 333112 224936
rect 263692 224816 263744 224868
rect 332876 224816 332928 224868
rect 260932 224748 260984 224800
rect 322480 224748 322532 224800
rect 261024 224680 261076 224732
rect 321008 224680 321060 224732
rect 259920 224612 259972 224664
rect 319536 224612 319588 224664
rect 249984 224544 250036 224596
rect 309324 224544 309376 224596
rect 234896 224476 234948 224528
rect 235632 224476 235684 224528
rect 290556 224476 290608 224528
rect 263140 224408 263192 224460
rect 316776 224408 316828 224460
rect 234804 224340 234856 224392
rect 235540 224340 235592 224392
rect 286600 224340 286652 224392
rect 358820 224340 358872 224392
rect 66904 224272 66956 224324
rect 226340 224272 226392 224324
rect 233516 224272 233568 224324
rect 275468 224272 275520 224324
rect 332784 224272 332836 224324
rect 406384 224272 406436 224324
rect 19984 224204 20036 224256
rect 223580 224204 223632 224256
rect 241520 224204 241572 224256
rect 249524 224204 249576 224256
rect 301412 224204 301464 224256
rect 332876 224204 332928 224256
rect 537484 224204 537536 224256
rect 255504 223524 255556 223576
rect 340972 223524 341024 223576
rect 341524 223524 341576 223576
rect 248512 223456 248564 223508
rect 331220 223456 331272 223508
rect 332048 223456 332100 223508
rect 251272 223388 251324 223440
rect 322940 223388 322992 223440
rect 264612 223320 264664 223372
rect 334256 223320 334308 223372
rect 334808 223320 334860 223372
rect 250996 223252 251048 223304
rect 311348 223252 311400 223304
rect 228364 223184 228416 223236
rect 228824 223184 228876 223236
rect 287612 223184 287664 223236
rect 257804 223116 257856 223168
rect 204260 223048 204312 223100
rect 237656 223048 237708 223100
rect 255136 223048 255188 223100
rect 302884 223048 302936 223100
rect 140780 222980 140832 223032
rect 233424 222980 233476 223032
rect 244096 222980 244148 223032
rect 273168 222980 273220 223032
rect 75920 222912 75972 222964
rect 228364 222912 228416 222964
rect 256884 222912 256936 222964
rect 313280 222912 313332 222964
rect 322940 222980 322992 223032
rect 323584 222980 323636 223032
rect 380900 222980 380952 223032
rect 317052 222912 317104 222964
rect 447784 222912 447836 222964
rect 33140 222844 33192 222896
rect 225052 222844 225104 222896
rect 226616 222844 226668 222896
rect 227076 222844 227128 222896
rect 287428 222844 287480 222896
rect 334808 222844 334860 222896
rect 543740 222844 543792 222896
rect 254400 222776 254452 222828
rect 255136 222776 255188 222828
rect 256884 222776 256936 222828
rect 229284 222096 229336 222148
rect 230112 222096 230164 222148
rect 241152 222096 241204 222148
rect 241520 222096 241572 222148
rect 249892 222096 249944 222148
rect 338488 222096 338540 222148
rect 339408 222096 339460 222148
rect 259644 222028 259696 222080
rect 329840 222028 329892 222080
rect 330300 222028 330352 222080
rect 236092 221960 236144 222012
rect 295708 221960 295760 222012
rect 254124 221892 254176 221944
rect 313280 221892 313332 221944
rect 237564 221824 237616 221876
rect 296076 221824 296128 221876
rect 223856 221756 223908 221808
rect 224132 221756 224184 221808
rect 282368 221756 282420 221808
rect 237196 221688 237248 221740
rect 287888 221688 287940 221740
rect 230112 221620 230164 221672
rect 278228 221620 278280 221672
rect 273168 221552 273220 221604
rect 305184 221552 305236 221604
rect 339408 221552 339460 221604
rect 362960 221552 363012 221604
rect 107660 221484 107712 221536
rect 230480 221484 230532 221536
rect 241520 221484 241572 221536
rect 297364 221484 297416 221536
rect 313280 221484 313332 221536
rect 314476 221484 314528 221536
rect 411904 221484 411956 221536
rect 17960 221416 18012 221468
rect 224132 221416 224184 221468
rect 264612 221416 264664 221468
rect 323768 221416 323820 221468
rect 330300 221416 330352 221468
rect 478144 221416 478196 221468
rect 222384 220736 222436 220788
rect 222936 220736 222988 220788
rect 226984 220736 227036 220788
rect 227260 220736 227312 220788
rect 228088 220736 228140 220788
rect 228548 220736 228600 220788
rect 249800 220736 249852 220788
rect 336832 220736 336884 220788
rect 338028 220736 338080 220788
rect 255412 220668 255464 220720
rect 340880 220668 340932 220720
rect 266544 220600 266596 220652
rect 338672 220600 338724 220652
rect 339408 220600 339460 220652
rect 228180 220532 228232 220584
rect 290280 220532 290332 220584
rect 180800 220464 180852 220516
rect 236092 220464 236144 220516
rect 256424 220464 256476 220516
rect 315856 220464 315908 220516
rect 340880 220464 340932 220516
rect 341616 220464 341668 220516
rect 226340 220396 226392 220448
rect 227168 220396 227220 220448
rect 286324 220396 286376 220448
rect 226984 220328 227036 220380
rect 284944 220328 284996 220380
rect 228548 220260 228600 220312
rect 286416 220260 286468 220312
rect 222936 220192 222988 220244
rect 282920 220192 282972 220244
rect 338028 220192 338080 220244
rect 353944 220192 353996 220244
rect 129740 220124 129792 220176
rect 232964 220124 233016 220176
rect 244556 220124 244608 220176
rect 285588 220124 285640 220176
rect 318708 220124 318760 220176
rect 426440 220124 426492 220176
rect 64880 220056 64932 220108
rect 226340 220056 226392 220108
rect 339408 220056 339460 220108
rect 568580 220056 568632 220108
rect 260840 219376 260892 219428
rect 332692 219376 332744 219428
rect 258356 219308 258408 219360
rect 323400 219308 323452 219360
rect 224316 219240 224368 219292
rect 283564 219240 283616 219292
rect 230296 219172 230348 219224
rect 287704 219172 287756 219224
rect 260748 219104 260800 219156
rect 319996 219104 320048 219156
rect 231584 219036 231636 219088
rect 283656 219036 283708 219088
rect 230204 218968 230256 219020
rect 280896 218968 280948 219020
rect 253480 218900 253532 218952
rect 303436 218900 303488 218952
rect 147680 218832 147732 218884
rect 233332 218832 233384 218884
rect 244464 218832 244516 218884
rect 288348 218832 288400 218884
rect 100760 218764 100812 218816
rect 230296 218764 230348 218816
rect 323400 218764 323452 218816
rect 462320 218764 462372 218816
rect 35900 218696 35952 218748
rect 225420 218696 225472 218748
rect 332692 218696 332744 218748
rect 500960 218696 501012 218748
rect 288348 218016 288400 218068
rect 289084 218016 289136 218068
rect 303436 218016 303488 218068
rect 394700 218016 394752 218068
rect 254032 217948 254084 218000
rect 338304 217948 338356 218000
rect 266820 217880 266872 217932
rect 338396 217880 338448 217932
rect 245844 217812 245896 217864
rect 300124 217812 300176 217864
rect 187700 217472 187752 217524
rect 237196 217472 237248 217524
rect 151820 217404 151872 217456
rect 233976 217404 234028 217456
rect 78680 217336 78732 217388
rect 227996 217336 228048 217388
rect 338304 217336 338356 217388
rect 415400 217336 415452 217388
rect 26240 217268 26292 217320
rect 224316 217268 224368 217320
rect 248236 217268 248288 217320
rect 322940 217268 322992 217320
rect 338396 217268 338448 217320
rect 565084 217268 565136 217320
rect 249340 216588 249392 216640
rect 338212 216588 338264 216640
rect 339408 216588 339460 216640
rect 266452 216520 266504 216572
rect 327172 216520 327224 216572
rect 328368 216520 328420 216572
rect 224868 216452 224920 216504
rect 282184 216452 282236 216504
rect 225052 216112 225104 216164
rect 239588 216112 239640 216164
rect 118700 216044 118752 216096
rect 231584 216044 231636 216096
rect 339408 216044 339460 216096
rect 349252 216044 349304 216096
rect 46204 215976 46256 216028
rect 224960 215976 225012 216028
rect 315856 215976 315908 216028
rect 430580 215976 430632 216028
rect 11060 215908 11112 215960
rect 222200 215908 222252 215960
rect 244188 215908 244240 215960
rect 266360 215908 266412 215960
rect 328368 215908 328420 215960
rect 575480 215908 575532 215960
rect 224316 215296 224368 215348
rect 224868 215296 224920 215348
rect 3332 215228 3384 215280
rect 91744 215228 91796 215280
rect 256792 215228 256844 215280
rect 334072 215228 334124 215280
rect 252192 215160 252244 215212
rect 328092 215160 328144 215212
rect 328368 215160 328420 215212
rect 264980 215092 265032 215144
rect 324320 215092 324372 215144
rect 168380 214684 168432 214736
rect 235448 214684 235500 214736
rect 328368 214684 328420 214736
rect 378784 214684 378836 214736
rect 91100 214616 91152 214668
rect 230204 214616 230256 214668
rect 334072 214616 334124 214668
rect 451280 214616 451332 214668
rect 50344 214548 50396 214600
rect 225236 214548 225288 214600
rect 242716 214548 242768 214600
rect 253204 214548 253256 214600
rect 324320 214548 324372 214600
rect 547144 214548 547196 214600
rect 253572 213868 253624 213920
rect 320732 213868 320784 213920
rect 256700 213800 256752 213852
rect 307668 213800 307720 213852
rect 205640 213256 205692 213308
rect 237564 213256 237616 213308
rect 320732 213256 320784 213308
rect 398932 213256 398984 213308
rect 29000 213188 29052 213240
rect 224040 213188 224092 213240
rect 307668 213188 307720 213240
rect 454684 213188 454736 213240
rect 262220 212440 262272 212492
rect 328552 212440 328604 212492
rect 329748 212440 329800 212492
rect 258080 212372 258132 212424
rect 318432 212372 318484 212424
rect 318708 212372 318760 212424
rect 162860 211896 162912 211948
rect 235632 211896 235684 211948
rect 55864 211828 55916 211880
rect 226984 211828 227036 211880
rect 318708 211828 318760 211880
rect 465080 211828 465132 211880
rect 40040 211760 40092 211812
rect 225512 211760 225564 211812
rect 329748 211760 329800 211812
rect 518900 211760 518952 211812
rect 253940 211080 253992 211132
rect 336740 211080 336792 211132
rect 338028 211080 338080 211132
rect 248144 211012 248196 211064
rect 307208 211012 307260 211064
rect 307668 211012 307720 211064
rect 259552 210944 259604 210996
rect 318800 210944 318852 210996
rect 320088 210944 320140 210996
rect 167000 210536 167052 210588
rect 235540 210536 235592 210588
rect 86960 210468 87012 210520
rect 230112 210468 230164 210520
rect 338028 210468 338080 210520
rect 417424 210468 417476 210520
rect 2780 210400 2832 210452
rect 223028 210400 223080 210452
rect 307668 210400 307720 210452
rect 318064 210400 318116 210452
rect 320088 210400 320140 210452
rect 476120 210400 476172 210452
rect 138664 209108 138716 209160
rect 232872 209108 232924 209160
rect 244372 209108 244424 209160
rect 292580 209108 292632 209160
rect 341616 209108 341668 209160
rect 425704 209108 425756 209160
rect 22100 209040 22152 209092
rect 224500 209040 224552 209092
rect 264520 209040 264572 209092
rect 530584 209040 530636 209092
rect 245752 208292 245804 208344
rect 305092 208292 305144 208344
rect 305092 207884 305144 207936
rect 306288 207884 306340 207936
rect 307024 207884 307076 207936
rect 190460 207680 190512 207732
rect 236736 207680 236788 207732
rect 67640 207612 67692 207664
rect 221648 207612 221700 207664
rect 341524 207612 341576 207664
rect 436744 207612 436796 207664
rect 233976 207544 234028 207596
rect 239496 207544 239548 207596
rect 269948 206932 270000 206984
rect 580172 206932 580224 206984
rect 201592 206388 201644 206440
rect 237472 206388 237524 206440
rect 155960 206320 156012 206372
rect 234160 206320 234212 206372
rect 55220 206252 55272 206304
rect 226892 206252 226944 206304
rect 258264 205572 258316 205624
rect 328460 205572 328512 205624
rect 329748 205572 329800 205624
rect 265992 205504 266044 205556
rect 324872 205504 324924 205556
rect 325332 205504 325384 205556
rect 121460 204960 121512 205012
rect 231952 204960 232004 205012
rect 329748 204960 329800 205012
rect 461584 204960 461636 205012
rect 80060 204892 80112 204944
rect 228732 204892 228784 204944
rect 324872 204892 324924 204944
rect 553400 204892 553452 204944
rect 258172 204212 258224 204264
rect 335360 204212 335412 204264
rect 336648 204212 336700 204264
rect 8300 203532 8352 203584
rect 222936 203532 222988 203584
rect 336648 203532 336700 203584
rect 472624 203532 472676 203584
rect 21364 202104 21416 202156
rect 222752 202104 222804 202156
rect 126244 200744 126296 200796
rect 232780 200744 232832 200796
rect 31024 199384 31076 199436
rect 223948 199384 224000 199436
rect 165620 198024 165672 198076
rect 235356 198024 235408 198076
rect 65524 197956 65576 198008
rect 227076 197956 227128 198008
rect 176752 196596 176804 196648
rect 236644 196596 236696 196648
rect 249432 196596 249484 196648
rect 340972 196596 341024 196648
rect 75184 195236 75236 195288
rect 228548 195236 228600 195288
rect 250812 195236 250864 195288
rect 357532 195236 357584 195288
rect 39304 193808 39356 193860
rect 225144 193808 225196 193860
rect 577596 193128 577648 193180
rect 579620 193128 579672 193180
rect 133880 192516 133932 192568
rect 232688 192516 232740 192568
rect 46296 192448 46348 192500
rect 225788 192448 225840 192500
rect 93952 191088 94004 191140
rect 230020 191088 230072 191140
rect 14464 189728 14516 189780
rect 222660 189728 222712 189780
rect 255044 189728 255096 189780
rect 415492 189728 415544 189780
rect 3516 188980 3568 189032
rect 213460 188980 213512 189032
rect 112444 186940 112496 186992
rect 231308 186940 231360 186992
rect 263324 186940 263376 186992
rect 521660 186940 521712 186992
rect 115940 185580 115992 185632
rect 231492 185580 231544 185632
rect 264612 185580 264664 185632
rect 535460 185580 535512 185632
rect 32404 184152 32456 184204
rect 223672 184152 223724 184204
rect 264704 184152 264756 184204
rect 539692 184152 539744 184204
rect 222200 181500 222252 181552
rect 239404 181500 239456 181552
rect 9680 181432 9732 181484
rect 222568 181432 222620 181484
rect 264796 181432 264848 181484
rect 542360 181432 542412 181484
rect 49700 180072 49752 180124
rect 225328 180072 225380 180124
rect 265716 180072 265768 180124
rect 559564 180072 559616 180124
rect 577504 179324 577556 179376
rect 579712 179324 579764 179376
rect 70400 178644 70452 178696
rect 228456 178644 228508 178696
rect 54484 177284 54536 177336
rect 226800 177284 226852 177336
rect 266176 177284 266228 177336
rect 564532 177284 564584 177336
rect 81440 175924 81492 175976
rect 220268 175924 220320 175976
rect 267372 175924 267424 175976
rect 563704 175924 563756 175976
rect 15844 174496 15896 174548
rect 222476 174496 222528 174548
rect 267556 174496 267608 174548
rect 571340 174496 571392 174548
rect 90364 173136 90416 173188
rect 229928 173136 229980 173188
rect 267280 173136 267332 173188
rect 578240 173136 578292 173188
rect 85672 171776 85724 171828
rect 220176 171776 220228 171828
rect 255136 171776 255188 171828
rect 411260 171776 411312 171828
rect 97264 170348 97316 170400
rect 229836 170348 229888 170400
rect 267648 170348 267700 170400
rect 574100 170348 574152 170400
rect 19340 168988 19392 169040
rect 218980 168988 219032 169040
rect 31760 167628 31812 167680
rect 224408 167628 224460 167680
rect 137284 166268 137336 166320
rect 232596 166268 232648 166320
rect 35992 164840 36044 164892
rect 215300 164840 215352 164892
rect 250904 164840 250956 164892
rect 361580 164840 361632 164892
rect 3240 164160 3292 164212
rect 199384 164160 199436 164212
rect 155316 162120 155368 162172
rect 234068 162120 234120 162172
rect 241612 162120 241664 162172
rect 251272 162120 251324 162172
rect 42800 160692 42852 160744
rect 206376 160692 206428 160744
rect 79324 159332 79376 159384
rect 228364 159332 228416 159384
rect 127072 157972 127124 158024
rect 232504 157972 232556 158024
rect 53840 155184 53892 155236
rect 227352 155184 227404 155236
rect 334624 153144 334676 153196
rect 580172 153144 580224 153196
rect 257988 149676 258040 149728
rect 454040 149676 454092 149728
rect 260748 145528 260800 145580
rect 478880 145528 478932 145580
rect 263416 144168 263468 144220
rect 512000 144168 512052 144220
rect 263508 141380 263560 141432
rect 519544 141380 519596 141432
rect 2872 137912 2924 137964
rect 203524 137912 203576 137964
rect 266268 137232 266320 137284
rect 555516 137232 555568 137284
rect 222016 126216 222068 126268
rect 580356 126216 580408 126268
rect 3424 111732 3476 111784
rect 211804 111732 211856 111784
rect 280068 100648 280120 100700
rect 579620 100648 579672 100700
rect 3424 97928 3476 97980
rect 198004 97928 198056 97980
rect 11152 90312 11204 90364
rect 209044 90312 209096 90364
rect 222108 87592 222160 87644
rect 580264 87592 580316 87644
rect 3148 85484 3200 85536
rect 192484 85484 192536 85536
rect 331864 73108 331916 73160
rect 580172 73108 580224 73160
rect 3424 71680 3476 71732
rect 186964 71680 187016 71732
rect 280804 60664 280856 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 195244 59304 195296 59356
rect 3424 45500 3476 45552
rect 206284 45500 206336 45552
rect 242808 33736 242860 33788
rect 255320 33736 255372 33788
rect 3424 32988 3476 33040
rect 7564 32988 7616 33040
rect 264888 29588 264940 29640
rect 527824 29588 527876 29640
rect 19432 24080 19484 24132
rect 188344 24080 188396 24132
rect 15200 22720 15252 22772
rect 222844 22720 222896 22772
rect 27620 21360 27672 21412
rect 213368 21360 213420 21412
rect 3424 20612 3476 20664
rect 43444 20612 43496 20664
rect 418804 20612 418856 20664
rect 580172 20612 580224 20664
rect 23480 18572 23532 18624
rect 214564 18572 214616 18624
rect 99380 17212 99432 17264
rect 217416 17212 217468 17264
rect 149520 14424 149572 14476
rect 233884 14424 233936 14476
rect 255228 14424 255280 14476
rect 422576 14424 422628 14476
rect 25320 13064 25372 13116
rect 224132 13064 224184 13116
rect 126980 11772 127032 11824
rect 128176 11772 128228 11824
rect 176660 11772 176712 11824
rect 177856 11772 177908 11824
rect 201500 11772 201552 11824
rect 202696 11772 202748 11824
rect 39120 11704 39172 11756
rect 224316 11704 224368 11756
rect 110512 10276 110564 10328
rect 230940 10276 230992 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 84476 8916 84528 8968
rect 227812 8916 227864 8968
rect 250996 8916 251048 8968
rect 369400 8916 369452 8968
rect 103336 7556 103388 7608
rect 229744 7556 229796 7608
rect 249616 7556 249668 7608
rect 344560 7556 344612 7608
rect 355324 7556 355376 7608
rect 474556 7556 474608 7608
rect 3424 6808 3476 6860
rect 116584 6808 116636 6860
rect 336096 6468 336148 6520
rect 460388 6468 460440 6520
rect 252652 6400 252704 6452
rect 394240 6400 394292 6452
rect 253848 6332 253900 6384
rect 397736 6332 397788 6384
rect 256516 6264 256568 6316
rect 429660 6264 429712 6316
rect 256608 6196 256660 6248
rect 433248 6196 433300 6248
rect 117596 6128 117648 6180
rect 231124 6128 231176 6180
rect 259368 6128 259420 6180
rect 461584 6128 461636 6180
rect 475384 5516 475436 5568
rect 478052 5516 478104 5568
rect 78588 4768 78640 4820
rect 227904 4768 227956 4820
rect 349804 4768 349856 4820
rect 449808 4768 449860 4820
rect 45468 4088 45520 4140
rect 46204 4088 46256 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 199108 4088 199160 4140
rect 216128 4088 216180 4140
rect 248328 4088 248380 4140
rect 249984 4088 250036 4140
rect 315304 4088 315356 4140
rect 318524 4088 318576 4140
rect 330576 4088 330628 4140
rect 336280 4088 336332 4140
rect 353944 4088 353996 4140
rect 193312 4020 193364 4072
rect 213276 4020 213328 4072
rect 251088 4020 251140 4072
rect 260656 4020 260708 4072
rect 275928 4020 275980 4072
rect 278320 4020 278372 4072
rect 329196 4020 329248 4072
rect 2872 3952 2924 4004
rect 7656 3952 7708 4004
rect 92756 3952 92808 4004
rect 95884 3952 95936 4004
rect 171968 3952 172020 4004
rect 215944 3952 215996 4004
rect 244924 3952 244976 4004
rect 257068 3952 257120 4004
rect 279424 3952 279476 4004
rect 288992 3952 289044 4004
rect 319444 3952 319496 4004
rect 331588 3952 331640 4004
rect 331956 4020 332008 4072
rect 335912 4020 335964 4072
rect 336004 4020 336056 4072
rect 339868 3952 339920 4004
rect 342904 4020 342956 4072
rect 354036 4020 354088 4072
rect 378784 4088 378836 4140
rect 384764 4088 384816 4140
rect 411996 4088 412048 4140
rect 413100 4088 413152 4140
rect 425704 4088 425756 4140
rect 434444 4088 434496 4140
rect 478144 4088 478196 4140
rect 480536 4088 480588 4140
rect 508504 4088 508556 4140
rect 510068 4088 510120 4140
rect 527824 4088 527876 4140
rect 530124 4088 530176 4140
rect 367008 4020 367060 4072
rect 357440 3952 357492 4004
rect 547144 3952 547196 4004
rect 550272 3952 550324 4004
rect 563704 3952 563756 4004
rect 568028 3952 568080 4004
rect 168472 3884 168524 3936
rect 215576 3884 215628 3936
rect 252284 3884 252336 3936
rect 372896 3884 372948 3936
rect 52552 3816 52604 3868
rect 55864 3816 55916 3868
rect 62028 3816 62080 3868
rect 66904 3816 66956 3868
rect 164884 3816 164936 3868
rect 220360 3816 220412 3868
rect 252468 3816 252520 3868
rect 376484 3816 376536 3868
rect 161296 3748 161348 3800
rect 218704 3748 218756 3800
rect 249708 3748 249760 3800
rect 259368 3748 259420 3800
rect 41880 3680 41932 3732
rect 46296 3680 46348 3732
rect 135260 3680 135312 3732
rect 138664 3680 138716 3732
rect 155408 3680 155460 3732
rect 218796 3680 218848 3732
rect 252376 3680 252428 3732
rect 253480 3680 253532 3732
rect 253664 3680 253716 3732
rect 259828 3680 259880 3732
rect 57244 3612 57296 3664
rect 1676 3544 1728 3596
rect 10324 3544 10376 3596
rect 7656 3476 7708 3528
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 14740 3544 14792 3596
rect 15844 3544 15896 3596
rect 46664 3544 46716 3596
rect 21364 3476 21416 3528
rect 21824 3476 21876 3528
rect 25504 3476 25556 3528
rect 31300 3476 31352 3528
rect 32404 3476 32456 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 38384 3476 38436 3528
rect 39304 3476 39356 3528
rect 48964 3476 49016 3528
rect 50344 3476 50396 3528
rect 53748 3544 53800 3596
rect 54484 3544 54536 3596
rect 59636 3544 59688 3596
rect 62764 3544 62816 3596
rect 69112 3612 69164 3664
rect 71044 3612 71096 3664
rect 96252 3612 96304 3664
rect 97264 3612 97316 3664
rect 109316 3612 109368 3664
rect 112444 3612 112496 3664
rect 121092 3612 121144 3664
rect 122104 3612 122156 3664
rect 123484 3612 123536 3664
rect 152464 3612 152516 3664
rect 160100 3612 160152 3664
rect 235264 3612 235316 3664
rect 246856 3612 246908 3664
rect 265348 3748 265400 3800
rect 278136 3748 278188 3800
rect 402520 3884 402572 3936
rect 537484 3884 537536 3936
rect 540796 3884 540848 3936
rect 260012 3680 260064 3732
rect 390560 3816 390612 3868
rect 574744 3816 574796 3868
rect 577412 3816 577464 3868
rect 385684 3680 385736 3732
rect 388260 3680 388312 3732
rect 400864 3680 400916 3732
rect 531320 3680 531372 3732
rect 260104 3612 260156 3664
rect 261760 3612 261812 3664
rect 269764 3612 269816 3664
rect 274824 3612 274876 3664
rect 123392 3544 123444 3596
rect 129372 3544 129424 3596
rect 210424 3544 210476 3596
rect 213184 3544 213236 3596
rect 226432 3544 226484 3596
rect 233976 3544 234028 3596
rect 242992 3544 243044 3596
rect 175924 3476 175976 3528
rect 186136 3476 186188 3528
rect 215668 3476 215720 3528
rect 238024 3476 238076 3528
rect 241336 3476 241388 3528
rect 244096 3476 244148 3528
rect 246948 3544 247000 3596
rect 270868 3544 270920 3596
rect 271144 3544 271196 3596
rect 285404 3612 285456 3664
rect 291844 3612 291896 3664
rect 306748 3612 306800 3664
rect 313924 3612 313976 3664
rect 317328 3612 317380 3664
rect 330484 3612 330536 3664
rect 485228 3612 485280 3664
rect 493324 3612 493376 3664
rect 552664 3612 552716 3664
rect 275284 3544 275336 3596
rect 267740 3476 267792 3528
rect 271236 3476 271288 3528
rect 272432 3476 272484 3528
rect 273904 3476 273956 3528
rect 276020 3476 276072 3528
rect 278044 3544 278096 3596
rect 296076 3544 296128 3596
rect 298744 3544 298796 3596
rect 6460 3408 6512 3460
rect 217324 3408 217376 3460
rect 226340 3408 226392 3460
rect 227536 3408 227588 3460
rect 229836 3408 229888 3460
rect 240784 3408 240836 3460
rect 241428 3408 241480 3460
rect 242900 3408 242952 3460
rect 245568 3408 245620 3460
rect 287796 3408 287848 3460
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 89168 3340 89220 3392
rect 90364 3340 90416 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 114008 3340 114060 3392
rect 115204 3340 115256 3392
rect 136456 3340 136508 3392
rect 137284 3340 137336 3392
rect 153016 3340 153068 3392
rect 155224 3340 155276 3392
rect 168380 3340 168432 3392
rect 169576 3340 169628 3392
rect 193220 3340 193272 3392
rect 194416 3340 194468 3392
rect 249524 3340 249576 3392
rect 251180 3340 251232 3392
rect 253204 3340 253256 3392
rect 254676 3340 254728 3392
rect 259368 3340 259420 3392
rect 264152 3340 264204 3392
rect 289084 3476 289136 3528
rect 290188 3476 290240 3528
rect 300124 3476 300176 3528
rect 301964 3476 302016 3528
rect 307024 3476 307076 3528
rect 309048 3476 309100 3528
rect 311164 3544 311216 3596
rect 312636 3544 312688 3596
rect 327724 3544 327776 3596
rect 329104 3544 329156 3596
rect 495900 3544 495952 3596
rect 498200 3544 498252 3596
rect 499028 3544 499080 3596
rect 500224 3544 500276 3596
rect 502892 3544 502944 3596
rect 502984 3544 503036 3596
rect 505376 3544 505428 3596
rect 554044 3544 554096 3596
rect 556160 3544 556212 3596
rect 313832 3476 313884 3528
rect 318064 3476 318116 3528
rect 319720 3476 319772 3528
rect 320824 3476 320876 3528
rect 325608 3476 325660 3528
rect 517152 3476 517204 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 526444 3476 526496 3528
rect 527824 3476 527876 3528
rect 536196 3476 536248 3528
rect 537208 3476 537260 3528
rect 540244 3476 540296 3528
rect 547880 3476 547932 3528
rect 555516 3476 555568 3528
rect 557356 3476 557408 3528
rect 559564 3476 559616 3528
rect 560852 3476 560904 3528
rect 289176 3408 289228 3460
rect 291384 3408 291436 3460
rect 295984 3408 296036 3460
rect 292580 3340 292632 3392
rect 299572 3408 299624 3460
rect 300768 3408 300820 3460
rect 305644 3408 305696 3460
rect 329196 3408 329248 3460
rect 329288 3408 329340 3460
rect 520740 3408 520792 3460
rect 529204 3408 529256 3460
rect 554964 3408 555016 3460
rect 555424 3408 555476 3460
rect 562048 3408 562100 3460
rect 565084 3408 565136 3460
rect 572720 3408 572772 3460
rect 299664 3340 299716 3392
rect 324964 3340 325016 3392
rect 326804 3340 326856 3392
rect 332048 3340 332100 3392
rect 342168 3340 342220 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 357532 3340 357584 3392
rect 358728 3340 358780 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 376024 3340 376076 3392
rect 377680 3340 377732 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 422944 3340 422996 3392
rect 424968 3340 425020 3392
rect 436744 3340 436796 3392
rect 437940 3340 437992 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 443644 3340 443696 3392
rect 445024 3340 445076 3392
rect 456892 3340 456944 3392
rect 458088 3340 458140 3392
rect 461676 3340 461728 3392
rect 469864 3340 469916 3392
rect 77392 3272 77444 3324
rect 79324 3272 79376 3324
rect 335912 3272 335964 3324
rect 343364 3272 343416 3324
rect 417516 3272 417568 3324
rect 420184 3272 420236 3324
rect 421564 3272 421616 3324
rect 423772 3272 423824 3324
rect 454684 3272 454736 3324
rect 455696 3272 455748 3324
rect 562324 3272 562376 3324
rect 565636 3272 565688 3324
rect 27712 3204 27764 3256
rect 31024 3204 31076 3256
rect 243636 3204 243688 3256
rect 248788 3204 248840 3256
rect 519636 3204 519688 3256
rect 525432 3204 525484 3256
rect 64328 3136 64380 3188
rect 65524 3136 65576 3188
rect 124680 3136 124732 3188
rect 126244 3136 126296 3188
rect 309876 3136 309928 3188
rect 315028 3136 315080 3188
rect 512644 3136 512696 3188
rect 515956 3136 516008 3188
rect 223948 3068 224000 3120
rect 226984 3068 227036 3120
rect 273168 3068 273220 3120
rect 277124 3068 277176 3120
rect 406384 3068 406436 3120
rect 409604 3068 409656 3120
rect 543004 3068 543056 3120
rect 545488 3068 545540 3120
rect 17040 3000 17092 3052
rect 19984 3000 20036 3052
rect 154212 3000 154264 3052
rect 155316 3000 155368 3052
rect 351276 3000 351328 3052
rect 352840 3000 352892 3052
rect 447784 3000 447836 3052
rect 448612 3000 448664 3052
rect 472624 3000 472676 3052
rect 473452 3000 473504 3052
rect 530584 3000 530636 3052
rect 532516 3000 532568 3052
rect 189724 2932 189776 2984
rect 191104 2932 191156 2984
rect 358084 2864 358136 2916
rect 361120 2864 361172 2916
rect 511356 2864 511408 2916
rect 513564 2864 513616 2916
rect 398840 2592 398892 2644
rect 400128 2592 400180 2644
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 699718 8156 703520
rect 24320 699718 24348 703520
rect 8116 699712 8168 699718
rect 8116 699654 8168 699660
rect 10324 699712 10376 699718
rect 10324 699654 10376 699660
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 26884 699712 26936 699718
rect 26884 699654 26936 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2778 527912 2834 527921
rect 2778 527847 2834 527856
rect 2792 527202 2820 527847
rect 2780 527196 2832 527202
rect 2780 527138 2832 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3436 376038 3464 579935
rect 4804 527196 4856 527202
rect 4804 527138 4856 527144
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 4816 380225 4844 527138
rect 7564 474768 7616 474774
rect 7564 474710 7616 474716
rect 7576 381585 7604 474710
rect 10336 388482 10364 699654
rect 14464 501016 14516 501022
rect 14464 500958 14516 500964
rect 14476 395350 14504 500958
rect 15844 448588 15896 448594
rect 15844 448530 15896 448536
rect 14464 395344 14516 395350
rect 14464 395286 14516 395292
rect 15856 391270 15884 448530
rect 26896 407794 26924 699654
rect 26884 407788 26936 407794
rect 26884 407730 26936 407736
rect 15844 391264 15896 391270
rect 15844 391206 15896 391212
rect 10324 388476 10376 388482
rect 10324 388418 10376 388424
rect 7562 381576 7618 381585
rect 7562 381511 7618 381520
rect 4802 380216 4858 380225
rect 4802 380151 4858 380160
rect 40052 378729 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 46204 553444 46256 553450
rect 46204 553386 46256 553392
rect 46216 389881 46244 553386
rect 46202 389872 46258 389881
rect 46202 389807 46258 389816
rect 71792 382974 71820 702986
rect 89180 699718 89208 703520
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 90364 699712 90416 699718
rect 90364 699654 90416 699660
rect 90376 403617 90404 699654
rect 90362 403608 90418 403617
rect 90362 403543 90418 403552
rect 71780 382968 71832 382974
rect 71780 382910 71832 382916
rect 40038 378720 40094 378729
rect 40038 378655 40094 378664
rect 3424 376032 3476 376038
rect 3424 375974 3476 375980
rect 104912 374649 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 387122 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700126 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700120 154172 700126
rect 154120 700062 154172 700068
rect 155224 700120 155276 700126
rect 155224 700062 155276 700068
rect 151084 422340 151136 422346
rect 151084 422282 151136 422288
rect 136640 387116 136692 387122
rect 136640 387058 136692 387064
rect 151096 384402 151124 422282
rect 155236 392630 155264 700062
rect 155224 392624 155276 392630
rect 155224 392566 155276 392572
rect 151084 384396 151136 384402
rect 151084 384338 151136 384344
rect 169772 377369 169800 702406
rect 201512 394058 201540 702986
rect 218992 698970 219020 703520
rect 218980 698964 219032 698970
rect 218980 698906 219032 698912
rect 201500 394052 201552 394058
rect 201500 393994 201552 394000
rect 169758 377360 169814 377369
rect 169758 377295 169814 377304
rect 104898 374640 104954 374649
rect 104898 374575 104954 374584
rect 230480 373380 230532 373386
rect 230480 373322 230532 373328
rect 229100 373040 229152 373046
rect 229100 372982 229152 372988
rect 3424 372632 3476 372638
rect 3424 372574 3476 372580
rect 3436 371385 3464 372574
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 227718 367704 227774 367713
rect 227718 367639 227774 367648
rect 226982 367568 227038 367577
rect 226982 367503 227038 367512
rect 224222 363624 224278 363633
rect 224222 363559 224278 363568
rect 223764 360256 223816 360262
rect 223764 360198 223816 360204
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 358086 3464 358391
rect 3424 358080 3476 358086
rect 3424 358022 3476 358028
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 220726 322144 220782 322153
rect 220726 322079 220782 322088
rect 217966 322008 218022 322017
rect 217966 321943 218022 321952
rect 213734 321872 213790 321881
rect 213734 321807 213790 321816
rect 213642 321600 213698 321609
rect 213642 321535 213698 321544
rect 211068 320612 211120 320618
rect 211068 320554 211120 320560
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 209688 318368 209740 318374
rect 209688 318310 209740 318316
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3424 293276 3476 293282
rect 3424 293218 3476 293224
rect 3436 293185 3464 293218
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 198004 291712 198056 291718
rect 198004 291654 198056 291660
rect 195244 291644 195296 291650
rect 195244 291586 195296 291592
rect 43442 291272 43498 291281
rect 43442 291207 43498 291216
rect 3516 290488 3568 290494
rect 3516 290430 3568 290436
rect 3424 286340 3476 286346
rect 3424 286282 3476 286288
rect 3436 254153 3464 286282
rect 3528 267209 3556 290430
rect 7562 289096 7618 289105
rect 7562 289031 7618 289040
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3516 253224 3568 253230
rect 3516 253166 3568 253172
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3424 239420 3476 239426
rect 3424 239362 3476 239368
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 2780 210452 2832 210458
rect 2780 210394 2832 210400
rect 2792 16574 2820 210394
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 149841 3464 239362
rect 3528 201929 3556 253166
rect 4158 237552 4214 237561
rect 4158 237487 4214 237496
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 2872 137964 2924 137970
rect 2872 137906 2924 137912
rect 2884 136785 2912 137906
rect 2870 136776 2926 136785
rect 2870 136711 2926 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 33040 3476 33046
rect 3424 32982 3476 32988
rect 3436 32473 3464 32982
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 237487
rect 7576 33046 7604 289031
rect 34518 236600 34574 236609
rect 34518 236535 34574 236544
rect 10324 229764 10376 229770
rect 10324 229706 10376 229712
rect 7656 227044 7708 227050
rect 7656 226986 7708 226992
rect 7564 33040 7616 33046
rect 7564 32982 7616 32988
rect 2792 16546 3648 16574
rect 4172 16546 5304 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 480 1716 3538
rect 2884 480 2912 3946
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 7668 4010 7696 226986
rect 8300 203584 8352 203590
rect 8300 203526 8352 203532
rect 8312 16574 8340 203526
rect 9680 181484 9732 181490
rect 9680 181426 9732 181432
rect 8312 16546 8800 16574
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 3470
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 181426
rect 10336 3602 10364 229706
rect 25502 226944 25558 226953
rect 25502 226879 25558 226888
rect 19984 224256 20036 224262
rect 19984 224198 20036 224204
rect 17960 221468 18012 221474
rect 17960 221410 18012 221416
rect 11060 215960 11112 215966
rect 11060 215902 11112 215908
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11072 3534 11100 215902
rect 14464 189780 14516 189786
rect 14464 189722 14516 189728
rect 11152 90364 11204 90370
rect 11152 90306 11204 90312
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 90306
rect 14476 3534 14504 189722
rect 15844 174548 15896 174554
rect 15844 174490 15896 174496
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15212 16574 15240 22714
rect 15212 16546 15792 16574
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 3470
rect 14752 480 14780 3538
rect 15764 3482 15792 16546
rect 15856 3602 15884 174490
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15764 3454 15976 3482
rect 15948 480 15976 3454
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17052 480 17080 2994
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 221410
rect 19340 169040 19392 169046
rect 19340 168982 19392 168988
rect 19352 6914 19380 168982
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19444 16574 19472 24074
rect 19444 16546 19932 16574
rect 19352 6886 19472 6914
rect 19444 480 19472 6886
rect 19904 490 19932 16546
rect 19996 3058 20024 224198
rect 22100 209092 22152 209098
rect 22100 209034 22152 209040
rect 21364 202156 21416 202162
rect 21364 202098 21416 202104
rect 21376 3534 21404 202098
rect 22112 16574 22140 209034
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 16574 23520 18566
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 19904 462 20300 490
rect 21836 480 21864 3470
rect 20272 354 20300 462
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25320 13116 25372 13122
rect 25320 13058 25372 13064
rect 25332 480 25360 13058
rect 25516 3534 25544 226879
rect 33140 222896 33192 222902
rect 33140 222838 33192 222844
rect 26240 217320 26292 217326
rect 26240 217262 26292 217268
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 217262
rect 29000 213240 29052 213246
rect 29000 213182 29052 213188
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27632 16574 27660 21354
rect 29012 16574 29040 213182
rect 31024 199436 31076 199442
rect 31024 199378 31076 199384
rect 27632 16546 28488 16574
rect 29012 16546 30144 16574
rect 27712 3256 27764 3262
rect 27712 3198 27764 3204
rect 27724 480 27752 3198
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 31036 3262 31064 199378
rect 32404 184204 32456 184210
rect 32404 184146 32456 184152
rect 31760 167680 31812 167686
rect 31760 167622 31812 167628
rect 31772 16574 31800 167622
rect 31772 16546 31984 16574
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31024 3256 31076 3262
rect 31024 3198 31076 3204
rect 31312 480 31340 3470
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 32416 3534 32444 184146
rect 33152 16574 33180 222838
rect 33152 16546 33640 16574
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 236535
rect 35900 218748 35952 218754
rect 35900 218690 35952 218696
rect 35912 3534 35940 218690
rect 40040 211812 40092 211818
rect 40040 211754 40092 211760
rect 39304 193860 39356 193866
rect 39304 193802 39356 193808
rect 35992 164892 36044 164898
rect 35992 164834 36044 164840
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 164834
rect 39120 11756 39172 11762
rect 39120 11698 39172 11704
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 3470
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 11698
rect 39316 3534 39344 193802
rect 40052 16574 40080 211754
rect 42800 160744 42852 160750
rect 42800 160686 42852 160692
rect 40052 16546 40264 16574
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41892 480 41920 3674
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 160686
rect 43456 20670 43484 291207
rect 116584 290556 116636 290562
rect 116584 290498 116636 290504
rect 91744 289128 91796 289134
rect 91744 289070 91796 289076
rect 85580 238060 85632 238066
rect 85580 238002 85632 238008
rect 60740 235272 60792 235278
rect 60740 235214 60792 235220
rect 44178 233880 44234 233889
rect 44178 233815 44234 233824
rect 43444 20664 43496 20670
rect 43444 20606 43496 20612
rect 44192 16574 44220 233815
rect 51078 231160 51134 231169
rect 51078 231095 51134 231104
rect 46940 228404 46992 228410
rect 46940 228346 46992 228352
rect 46204 216028 46256 216034
rect 46204 215970 46256 215976
rect 44192 16546 44312 16574
rect 44284 480 44312 16546
rect 46216 4146 46244 215970
rect 46296 192500 46348 192506
rect 46296 192442 46348 192448
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 45480 480 45508 4082
rect 46308 3738 46336 192442
rect 46952 16574 46980 228346
rect 50344 214600 50396 214606
rect 50344 214542 50396 214548
rect 49700 180124 49752 180130
rect 49700 180066 49752 180072
rect 49712 16574 49740 180066
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 46296 3732 46348 3738
rect 46296 3674 46348 3680
rect 46664 3596 46716 3602
rect 46664 3538 46716 3544
rect 46676 480 46704 3538
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 48976 480 49004 3470
rect 50172 480 50200 16546
rect 50356 3534 50384 214542
rect 50344 3528 50396 3534
rect 50344 3470 50396 3476
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 231095
rect 57978 225584 58034 225593
rect 57978 225519 58034 225528
rect 55864 211880 55916 211886
rect 55864 211822 55916 211828
rect 55220 206304 55272 206310
rect 55220 206246 55272 206252
rect 54484 177336 54536 177342
rect 54484 177278 54536 177284
rect 53840 155236 53892 155242
rect 53840 155178 53892 155184
rect 53852 16574 53880 155178
rect 53852 16546 54432 16574
rect 52552 3868 52604 3874
rect 52552 3810 52604 3816
rect 52564 480 52592 3810
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 53760 480 53788 3538
rect 54404 3482 54432 16546
rect 54496 3602 54524 177278
rect 55232 16574 55260 206246
rect 55232 16546 55812 16574
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 55784 3482 55812 16546
rect 55876 3874 55904 211822
rect 57992 16574 58020 225519
rect 60752 16574 60780 235214
rect 62764 232552 62816 232558
rect 62764 232494 62816 232500
rect 62118 200696 62174 200705
rect 62118 200631 62174 200640
rect 62132 16574 62160 200631
rect 57992 16546 58480 16574
rect 60752 16546 60872 16574
rect 62132 16546 62712 16574
rect 55864 3868 55916 3874
rect 55864 3810 55916 3816
rect 57244 3664 57296 3670
rect 57244 3606 57296 3612
rect 54404 3454 54984 3482
rect 55784 3454 56088 3482
rect 54956 480 54984 3454
rect 56060 480 56088 3454
rect 57256 480 57284 3606
rect 58452 480 58480 16546
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59648 480 59676 3538
rect 60844 480 60872 16546
rect 62028 3868 62080 3874
rect 62028 3810 62080 3816
rect 62040 480 62068 3810
rect 62684 3482 62712 16546
rect 62776 3602 62804 232494
rect 74540 231124 74592 231130
rect 74540 231066 74592 231072
rect 71042 229800 71098 229809
rect 71042 229735 71098 229744
rect 66904 224324 66956 224330
rect 66904 224266 66956 224272
rect 64880 220108 64932 220114
rect 64880 220050 64932 220056
rect 64892 16574 64920 220050
rect 65524 198008 65576 198014
rect 65524 197950 65576 197956
rect 64892 16546 65104 16574
rect 62764 3596 62816 3602
rect 62764 3538 62816 3544
rect 62684 3454 63264 3482
rect 63236 480 63264 3454
rect 64328 3188 64380 3194
rect 64328 3130 64380 3136
rect 64340 480 64368 3130
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 65536 3194 65564 197950
rect 66258 196616 66314 196625
rect 66258 196551 66314 196560
rect 66272 16574 66300 196551
rect 66272 16546 66760 16574
rect 65524 3188 65576 3194
rect 65524 3130 65576 3136
rect 66732 480 66760 16546
rect 66916 3874 66944 224266
rect 69018 213208 69074 213217
rect 69018 213143 69074 213152
rect 67640 207664 67692 207670
rect 67640 207606 67692 207612
rect 66904 3868 66956 3874
rect 66904 3810 66956 3816
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 207606
rect 69032 16574 69060 213143
rect 70400 178696 70452 178702
rect 70400 178638 70452 178644
rect 70412 16574 70440 178638
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3664 69164 3670
rect 69112 3606 69164 3612
rect 69124 480 69152 3606
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3670 71084 229735
rect 71778 228304 71834 228313
rect 71778 228239 71834 228248
rect 71792 16574 71820 228239
rect 74552 16574 74580 231066
rect 75920 222964 75972 222970
rect 75920 222906 75972 222912
rect 75184 195288 75236 195294
rect 75184 195230 75236 195236
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 71044 3664 71096 3670
rect 71044 3606 71096 3612
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 195230
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 222906
rect 82818 222864 82874 222873
rect 82818 222799 82874 222808
rect 78680 217388 78732 217394
rect 78680 217330 78732 217336
rect 78692 16574 78720 217330
rect 80060 204944 80112 204950
rect 80060 204886 80112 204892
rect 79324 159384 79376 159390
rect 79324 159326 79376 159332
rect 78692 16546 79272 16574
rect 78588 4820 78640 4826
rect 78588 4762 78640 4768
rect 77392 3324 77444 3330
rect 77392 3266 77444 3272
rect 77404 480 77432 3266
rect 78600 480 78628 4762
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 79336 3330 79364 159326
rect 80072 16574 80100 204886
rect 81440 175976 81492 175982
rect 81440 175918 81492 175924
rect 81452 16574 81480 175918
rect 82832 16574 82860 222799
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 79324 3324 79376 3330
rect 79324 3266 79376 3272
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84476 8968 84528 8974
rect 84476 8910 84528 8916
rect 84488 480 84516 8910
rect 85592 3398 85620 238002
rect 89720 232620 89772 232626
rect 89720 232562 89772 232568
rect 86960 210520 87012 210526
rect 86960 210462 87012 210468
rect 85672 171828 85724 171834
rect 85672 171770 85724 171776
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 85684 480 85712 171770
rect 86972 16574 87000 210462
rect 89732 16574 89760 232562
rect 91756 215286 91784 289070
rect 103520 239488 103572 239494
rect 103520 239430 103572 239436
rect 95884 235408 95936 235414
rect 95884 235350 95936 235356
rect 93858 224224 93914 224233
rect 93858 224159 93914 224168
rect 91744 215280 91796 215286
rect 91744 215222 91796 215228
rect 91100 214668 91152 214674
rect 91100 214610 91152 214616
rect 90364 173188 90416 173194
rect 90364 173130 90416 173136
rect 86972 16546 87552 16574
rect 89732 16546 89944 16574
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89180 480 89208 3334
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 90376 3398 90404 173130
rect 91112 16574 91140 214610
rect 91112 16546 91600 16574
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91572 480 91600 16546
rect 93872 6914 93900 224159
rect 93952 191140 94004 191146
rect 93952 191082 94004 191088
rect 93964 16574 93992 191082
rect 93964 16546 94728 16574
rect 93872 6886 93992 6914
rect 92756 4004 92808 4010
rect 92756 3946 92808 3952
rect 92768 480 92796 3946
rect 93964 480 93992 6886
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95896 4010 95924 235350
rect 97998 234016 98054 234025
rect 97998 233951 98054 233960
rect 96620 228472 96672 228478
rect 96620 228414 96672 228420
rect 96632 16574 96660 228414
rect 97264 170400 97316 170406
rect 97264 170342 97316 170348
rect 96632 16546 97212 16574
rect 95884 4004 95936 4010
rect 95884 3946 95936 3952
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 96264 480 96292 3606
rect 97184 3482 97212 16546
rect 97276 3670 97304 170342
rect 98012 16574 98040 233951
rect 100760 218816 100812 218822
rect 100760 218758 100812 218764
rect 99380 17264 99432 17270
rect 99380 17206 99432 17212
rect 99392 16574 99420 17206
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 97264 3664 97316 3670
rect 97264 3606 97316 3612
rect 97184 3454 97488 3482
rect 97460 480 97488 3454
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 218758
rect 102138 199336 102194 199345
rect 102138 199271 102194 199280
rect 102152 16574 102180 199271
rect 103532 16574 103560 239430
rect 115204 235476 115256 235482
rect 115204 235418 115256 235424
rect 106280 235340 106332 235346
rect 106280 235282 106332 235288
rect 104898 203552 104954 203561
rect 104898 203487 104954 203496
rect 104912 16574 104940 203487
rect 106292 16574 106320 235282
rect 111800 232688 111852 232694
rect 111800 232630 111852 232636
rect 110418 229936 110474 229945
rect 110418 229871 110474 229880
rect 107660 221536 107712 221542
rect 107660 221478 107712 221484
rect 107672 16574 107700 221478
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 7608 103388 7614
rect 103336 7550 103388 7556
rect 103348 480 103376 7550
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109316 3664 109368 3670
rect 109316 3606 109368 3612
rect 109328 480 109356 3606
rect 110432 3398 110460 229871
rect 111812 16574 111840 232630
rect 114558 220280 114614 220289
rect 114558 220215 114614 220224
rect 112444 186992 112496 186998
rect 112444 186934 112496 186940
rect 111812 16546 112392 16574
rect 110512 10328 110564 10334
rect 110512 10270 110564 10276
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 10270
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 112456 3670 112484 186934
rect 114572 16574 114600 220215
rect 114572 16546 114784 16574
rect 112444 3664 112496 3670
rect 112444 3606 112496 3612
rect 114008 3392 114060 3398
rect 114008 3334 114060 3340
rect 114020 480 114048 3334
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 115216 3398 115244 235418
rect 115940 185632 115992 185638
rect 115940 185574 115992 185580
rect 115952 16574 115980 185574
rect 115952 16546 116440 16574
rect 115204 3392 115256 3398
rect 115204 3334 115256 3340
rect 116412 480 116440 16546
rect 116596 6866 116624 290498
rect 192484 289876 192536 289882
rect 192484 289818 192536 289824
rect 186962 289232 187018 289241
rect 186962 289167 187018 289176
rect 161480 240780 161532 240786
rect 161480 240722 161532 240728
rect 139400 239624 139452 239630
rect 139400 239566 139452 239572
rect 125600 239556 125652 239562
rect 125600 239498 125652 239504
rect 123484 227180 123536 227186
rect 123484 227122 123536 227128
rect 122104 227112 122156 227118
rect 122104 227054 122156 227060
rect 118700 216096 118752 216102
rect 118700 216038 118752 216044
rect 118712 6914 118740 216038
rect 121460 205012 121512 205018
rect 121460 204954 121512 204960
rect 118790 182880 118846 182889
rect 118790 182815 118846 182824
rect 118804 16574 118832 182815
rect 121472 16574 121500 204954
rect 118804 16546 119936 16574
rect 121472 16546 122052 16574
rect 118712 6886 118832 6914
rect 116584 6860 116636 6866
rect 116584 6802 116636 6808
rect 117596 6180 117648 6186
rect 117596 6122 117648 6128
rect 117608 480 117636 6122
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 121092 3664 121144 3670
rect 121092 3606 121144 3612
rect 121104 480 121132 3606
rect 122024 3482 122052 16546
rect 122116 3670 122144 227054
rect 123496 6914 123524 227122
rect 123404 6886 123524 6914
rect 122104 3664 122156 3670
rect 122104 3606 122156 3612
rect 123404 3602 123432 6886
rect 123484 3664 123536 3670
rect 123484 3606 123536 3612
rect 123392 3596 123444 3602
rect 123392 3538 123444 3544
rect 122024 3454 122328 3482
rect 122300 480 122328 3454
rect 123496 480 123524 3606
rect 124680 3188 124732 3194
rect 124680 3130 124732 3136
rect 124692 480 124720 3130
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 239498
rect 126980 236700 127032 236706
rect 126980 236642 127032 236648
rect 126244 200796 126296 200802
rect 126244 200738 126296 200744
rect 126256 3194 126284 200738
rect 126992 11830 127020 236642
rect 132500 232756 132552 232762
rect 132500 232698 132552 232704
rect 131118 221504 131174 221513
rect 131118 221439 131174 221448
rect 129740 220176 129792 220182
rect 129740 220118 129792 220124
rect 127072 158024 127124 158030
rect 127072 157966 127124 157972
rect 126980 11824 127032 11830
rect 126980 11766 127032 11772
rect 127084 6914 127112 157966
rect 129752 16574 129780 220118
rect 131132 16574 131160 221439
rect 132512 16574 132540 232698
rect 138018 232520 138074 232529
rect 138018 232455 138074 232464
rect 136640 225616 136692 225622
rect 136640 225558 136692 225564
rect 133880 192568 133932 192574
rect 133880 192510 133932 192516
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128176 11824 128228 11830
rect 128176 11766 128228 11772
rect 126992 6886 127112 6914
rect 126244 3188 126296 3194
rect 126244 3130 126296 3136
rect 126992 480 127020 6886
rect 128188 480 128216 11766
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 129384 480 129412 3538
rect 130580 480 130608 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 192510
rect 136652 16574 136680 225558
rect 137284 166320 137336 166326
rect 137284 166262 137336 166268
rect 136652 16546 137232 16574
rect 135260 3732 135312 3738
rect 135260 3674 135312 3680
rect 135272 480 135300 3674
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 136468 480 136496 3334
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 3398 137324 166262
rect 138032 16574 138060 232455
rect 138664 209160 138716 209166
rect 138664 209102 138716 209108
rect 138032 16546 138612 16574
rect 138584 3482 138612 16546
rect 138676 3738 138704 209102
rect 139412 16574 139440 239566
rect 157340 237448 157392 237454
rect 157340 237390 157392 237396
rect 152462 235240 152518 235249
rect 152462 235175 152518 235184
rect 143540 233912 143592 233918
rect 143540 233854 143592 233860
rect 140780 223032 140832 223038
rect 140780 222974 140832 222980
rect 140792 16574 140820 222974
rect 142158 207632 142214 207641
rect 142158 207567 142214 207576
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 138664 3732 138716 3738
rect 138664 3674 138716 3680
rect 138584 3454 138888 3482
rect 137284 3392 137336 3398
rect 137284 3334 137336 3340
rect 138860 480 138888 3454
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 207567
rect 143552 480 143580 233854
rect 150440 228540 150492 228546
rect 150440 228482 150492 228488
rect 146300 225684 146352 225690
rect 146300 225626 146352 225632
rect 143630 193896 143686 193905
rect 143630 193831 143686 193840
rect 143644 16574 143672 193831
rect 144918 188320 144974 188329
rect 144918 188255 144974 188264
rect 144932 16574 144960 188255
rect 146312 16574 146340 225626
rect 147680 218884 147732 218890
rect 147680 218826 147732 218832
rect 147692 16574 147720 218826
rect 150452 16574 150480 228482
rect 151820 217456 151872 217462
rect 151820 217398 151872 217404
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149520 14476 149572 14482
rect 149520 14418 149572 14424
rect 149532 480 149560 14418
rect 150636 480 150664 16546
rect 151832 480 151860 217398
rect 152476 3670 152504 235175
rect 155222 231432 155278 231441
rect 155222 231367 155278 231376
rect 152464 3664 152516 3670
rect 152464 3606 152516 3612
rect 155236 3398 155264 231367
rect 155960 206372 156012 206378
rect 155960 206314 156012 206320
rect 155316 162172 155368 162178
rect 155316 162114 155368 162120
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 155224 3392 155276 3398
rect 155224 3334 155276 3340
rect 153028 480 153056 3334
rect 155328 3058 155356 162114
rect 155972 16574 156000 206314
rect 157352 16574 157380 237390
rect 158718 224360 158774 224369
rect 158718 224295 158774 224304
rect 158732 16574 158760 224295
rect 161492 16574 161520 240722
rect 182180 239760 182232 239766
rect 182180 239702 182232 239708
rect 175280 239692 175332 239698
rect 175280 239634 175332 239640
rect 173898 236872 173954 236881
rect 173898 236807 173954 236816
rect 169758 236736 169814 236745
rect 169758 236671 169814 236680
rect 168380 214736 168432 214742
rect 168380 214678 168432 214684
rect 162860 211948 162912 211954
rect 162860 211890 162912 211896
rect 162872 16574 162900 211890
rect 167000 210588 167052 210594
rect 167000 210530 167052 210536
rect 165620 198076 165672 198082
rect 165620 198018 165672 198024
rect 165632 16574 165660 198018
rect 167012 16574 167040 210530
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 155408 3732 155460 3738
rect 155408 3674 155460 3680
rect 154212 3052 154264 3058
rect 154212 2994 154264 3000
rect 155316 3052 155368 3058
rect 155316 2994 155368 3000
rect 154224 480 154252 2994
rect 155420 480 155448 3674
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 161296 3800 161348 3806
rect 161296 3742 161348 3748
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 160112 480 160140 3606
rect 161308 480 161336 3742
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 164884 3868 164936 3874
rect 164884 3810 164936 3816
rect 164896 480 164924 3810
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 3398 168420 214678
rect 169772 16574 169800 236671
rect 172520 228608 172572 228614
rect 172520 228550 172572 228556
rect 172532 16574 172560 228550
rect 169772 16546 170352 16574
rect 172532 16546 172744 16574
rect 168472 3936 168524 3942
rect 168472 3878 168524 3884
rect 168380 3392 168432 3398
rect 168380 3334 168432 3340
rect 168484 1578 168512 3878
rect 169576 3392 169628 3398
rect 169576 3334 169628 3340
rect 168392 1550 168512 1578
rect 168392 480 168420 1550
rect 169588 480 169616 3334
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171968 4004 172020 4010
rect 171968 3946 172020 3952
rect 171980 480 172008 3946
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 236807
rect 175292 16574 175320 239634
rect 178040 239352 178092 239358
rect 178040 239294 178092 239300
rect 176658 237008 176714 237017
rect 176658 236943 176714 236952
rect 175924 235544 175976 235550
rect 175924 235486 175976 235492
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 175936 3534 175964 235486
rect 176672 11830 176700 236943
rect 176752 196648 176804 196654
rect 176752 196590 176804 196596
rect 176660 11824 176712 11830
rect 176660 11766 176712 11772
rect 176764 6914 176792 196590
rect 178052 16574 178080 239294
rect 179420 229832 179472 229838
rect 179420 229774 179472 229780
rect 179432 16574 179460 229774
rect 180800 220516 180852 220522
rect 180800 220458 180852 220464
rect 180812 16574 180840 220458
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 11824 177908 11830
rect 177856 11766 177908 11772
rect 176672 6886 176792 6914
rect 175924 3528 175976 3534
rect 175924 3470 175976 3476
rect 176672 480 176700 6886
rect 177868 480 177896 11766
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 239702
rect 184938 237280 184994 237289
rect 184938 237215 184994 237224
rect 183560 232824 183612 232830
rect 183560 232766 183612 232772
rect 183572 16574 183600 232766
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 480 184980 237215
rect 186320 227248 186372 227254
rect 186320 227190 186372 227196
rect 186332 16574 186360 227190
rect 186976 71738 187004 289167
rect 188342 237960 188398 237969
rect 188342 237895 188398 237904
rect 187700 217524 187752 217530
rect 187700 217466 187752 217472
rect 186964 71732 187016 71738
rect 186964 71674 187016 71680
rect 187712 16574 187740 217466
rect 188356 24138 188384 237895
rect 191840 236768 191892 236774
rect 191840 236710 191892 236716
rect 191104 232892 191156 232898
rect 191104 232834 191156 232840
rect 190460 207732 190512 207738
rect 190460 207674 190512 207680
rect 188344 24132 188396 24138
rect 188344 24074 188396 24080
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 186136 3528 186188 3534
rect 186136 3470 186188 3476
rect 186148 480 186176 3470
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189724 2984 189776 2990
rect 189724 2926 189776 2932
rect 189736 480 189764 2926
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 207674
rect 191116 2990 191144 232834
rect 191852 16574 191880 236710
rect 192496 85542 192524 289818
rect 193220 240848 193272 240854
rect 193220 240790 193272 240796
rect 192484 85536 192536 85542
rect 192484 85478 192536 85484
rect 191852 16546 192064 16574
rect 191104 2984 191156 2990
rect 191104 2926 191156 2932
rect 192036 480 192064 16546
rect 193232 3398 193260 240790
rect 194600 238128 194652 238134
rect 194600 238070 194652 238076
rect 194612 16574 194640 238070
rect 195256 59362 195284 291586
rect 197360 239828 197412 239834
rect 197360 239770 197412 239776
rect 195980 239216 196032 239222
rect 195980 239158 196032 239164
rect 195244 59356 195296 59362
rect 195244 59298 195296 59304
rect 195992 16574 196020 239158
rect 197372 16574 197400 239770
rect 198016 97986 198044 291654
rect 206282 291408 206338 291417
rect 206282 291343 206338 291352
rect 203524 289944 203576 289950
rect 203524 289886 203576 289892
rect 199384 289196 199436 289202
rect 199384 289138 199436 289144
rect 199396 164218 199424 289138
rect 202880 240916 202932 240922
rect 202880 240858 202932 240864
rect 200120 239284 200172 239290
rect 200120 239226 200172 239232
rect 199384 164212 199436 164218
rect 199384 164154 199436 164160
rect 198004 97980 198056 97986
rect 198004 97922 198056 97928
rect 200132 16574 200160 239226
rect 201498 237144 201554 237153
rect 201498 237079 201554 237088
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 200132 16546 200344 16574
rect 193312 4072 193364 4078
rect 193312 4014 193364 4020
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 193324 1442 193352 4014
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 193232 1414 193352 1442
rect 193232 480 193260 1414
rect 194428 480 194456 3334
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 199108 4140 199160 4146
rect 199108 4082 199160 4088
rect 199120 480 199148 4082
rect 200316 480 200344 16546
rect 201512 11830 201540 237079
rect 201592 206440 201644 206446
rect 201592 206382 201644 206388
rect 201500 11824 201552 11830
rect 201500 11766 201552 11772
rect 201604 6914 201632 206382
rect 202892 16574 202920 240858
rect 203536 137970 203564 289886
rect 204260 223100 204312 223106
rect 204260 223042 204312 223048
rect 203524 137964 203576 137970
rect 203524 137906 203576 137912
rect 204272 16574 204300 223042
rect 205640 213308 205692 213314
rect 205640 213250 205692 213256
rect 205652 16574 205680 213250
rect 206296 45558 206324 291343
rect 207020 239964 207072 239970
rect 207020 239906 207072 239912
rect 206376 238740 206428 238746
rect 206376 238682 206428 238688
rect 206388 160750 206416 238682
rect 206376 160744 206428 160750
rect 206376 160686 206428 160692
rect 206284 45552 206336 45558
rect 206284 45494 206336 45500
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202696 11824 202748 11830
rect 202696 11766 202748 11772
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11766
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 239906
rect 209700 238513 209728 318310
rect 210976 308440 211028 308446
rect 210976 308382 211028 308388
rect 210424 240100 210476 240106
rect 210424 240042 210476 240048
rect 209686 238504 209742 238513
rect 209686 238439 209742 238448
rect 209042 237824 209098 237833
rect 209042 237759 209098 237768
rect 208398 231296 208454 231305
rect 208398 231231 208454 231240
rect 208412 16574 208440 231231
rect 209056 90370 209084 237759
rect 209780 235680 209832 235686
rect 209780 235622 209832 235628
rect 209044 90364 209096 90370
rect 209044 90306 209096 90312
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 235622
rect 209870 224496 209926 224505
rect 209870 224431 209926 224440
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 224431
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210436 3602 210464 240042
rect 210988 236638 211016 308382
rect 210976 236632 211028 236638
rect 210976 236574 211028 236580
rect 210698 235920 210754 235929
rect 210698 235855 210754 235864
rect 210712 233889 210740 235855
rect 210698 233880 210754 233889
rect 210698 233815 210754 233824
rect 210988 232558 211016 236574
rect 211080 235929 211108 320554
rect 212170 318472 212226 318481
rect 212170 318407 212226 318416
rect 212078 318200 212134 318209
rect 212078 318135 212134 318144
rect 211986 307184 212042 307193
rect 211986 307119 212042 307128
rect 211804 289264 211856 289270
rect 211804 289206 211856 289212
rect 211066 235920 211122 235929
rect 211066 235855 211122 235864
rect 211160 235612 211212 235618
rect 211160 235554 211212 235560
rect 210976 232552 211028 232558
rect 210976 232494 211028 232500
rect 211172 16574 211200 235554
rect 211816 111790 211844 289206
rect 212000 236473 212028 307119
rect 212092 238746 212120 318135
rect 212080 238740 212132 238746
rect 212080 238682 212132 238688
rect 212184 237833 212212 318407
rect 212354 318336 212410 318345
rect 212264 318300 212316 318306
rect 212354 318271 212410 318280
rect 212264 318242 212316 318248
rect 212276 238542 212304 318242
rect 212264 238536 212316 238542
rect 212264 238478 212316 238484
rect 212170 237824 212226 237833
rect 212170 237759 212226 237768
rect 212368 237386 212396 318271
rect 212446 318064 212502 318073
rect 212446 317999 212502 318008
rect 212356 237380 212408 237386
rect 212356 237322 212408 237328
rect 211986 236464 212042 236473
rect 211986 236399 212042 236408
rect 212460 235958 212488 317999
rect 213368 316736 213420 316742
rect 213368 316678 213420 316684
rect 213276 309188 213328 309194
rect 213276 309130 213328 309136
rect 213288 241097 213316 309130
rect 213274 241088 213330 241097
rect 213274 241023 213330 241032
rect 213288 238754 213316 241023
rect 213380 239970 213408 316678
rect 213550 314392 213606 314401
rect 213550 314327 213606 314336
rect 213460 290012 213512 290018
rect 213460 289954 213512 289960
rect 213368 239964 213420 239970
rect 213368 239906 213420 239912
rect 213104 238726 213316 238754
rect 212448 235952 212500 235958
rect 212448 235894 212500 235900
rect 212460 235414 212488 235894
rect 212448 235408 212500 235414
rect 212448 235350 212500 235356
rect 213104 225593 213132 238726
rect 213368 238196 213420 238202
rect 213368 238138 213420 238144
rect 213184 237516 213236 237522
rect 213184 237458 213236 237464
rect 213090 225584 213146 225593
rect 213090 225519 213146 225528
rect 212538 221640 212594 221649
rect 212538 221575 212594 221584
rect 211804 111784 211856 111790
rect 211804 111726 211856 111732
rect 212552 16574 212580 221575
rect 211172 16546 211752 16574
rect 212552 16546 213132 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 210424 3596 210476 3602
rect 210424 3538 210476 3544
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213104 3482 213132 16546
rect 213196 3602 213224 237458
rect 213276 235408 213328 235414
rect 213276 235350 213328 235356
rect 213288 4078 213316 235350
rect 213380 21418 213408 238138
rect 213472 189038 213500 289954
rect 213564 236502 213592 314327
rect 213656 240553 213684 321535
rect 213642 240544 213698 240553
rect 213642 240479 213698 240488
rect 213552 236496 213604 236502
rect 213552 236438 213604 236444
rect 213564 232626 213592 236438
rect 213552 232620 213604 232626
rect 213552 232562 213604 232568
rect 213656 228313 213684 240479
rect 213748 235793 213776 321807
rect 215114 316704 215170 316713
rect 215114 316639 215170 316648
rect 215024 315308 215076 315314
rect 215024 315250 215076 315256
rect 213828 311976 213880 311982
rect 213828 311918 213880 311924
rect 213734 235784 213790 235793
rect 213734 235719 213790 235728
rect 213642 228304 213698 228313
rect 213642 228239 213698 228248
rect 213748 226953 213776 235719
rect 213734 226944 213790 226953
rect 213734 226879 213790 226888
rect 213840 223553 213868 311918
rect 214932 309936 214984 309942
rect 214932 309878 214984 309884
rect 214564 309800 214616 309806
rect 214564 309742 214616 309748
rect 214838 309768 214894 309777
rect 214470 307048 214526 307057
rect 214470 306983 214526 306992
rect 214380 240508 214432 240514
rect 214380 240450 214432 240456
rect 214392 239562 214420 240450
rect 214484 240446 214512 306983
rect 214472 240440 214524 240446
rect 214472 240382 214524 240388
rect 214380 239556 214432 239562
rect 214380 239498 214432 239504
rect 214484 236366 214512 240382
rect 214576 239494 214604 309742
rect 214838 309703 214894 309712
rect 214656 308508 214708 308514
rect 214656 308450 214708 308456
rect 214564 239488 214616 239494
rect 214564 239430 214616 239436
rect 214564 238264 214616 238270
rect 214564 238206 214616 238212
rect 213920 236360 213972 236366
rect 213920 236302 213972 236308
rect 214472 236360 214524 236366
rect 214472 236302 214524 236308
rect 213826 223544 213882 223553
rect 213826 223479 213882 223488
rect 213840 222873 213868 223479
rect 213826 222864 213882 222873
rect 213826 222799 213882 222808
rect 213460 189032 213512 189038
rect 213460 188974 213512 188980
rect 213368 21412 213420 21418
rect 213368 21354 213420 21360
rect 213932 16574 213960 236302
rect 214576 18630 214604 238206
rect 214668 238066 214696 308450
rect 214748 307216 214800 307222
rect 214748 307158 214800 307164
rect 214656 238060 214708 238066
rect 214656 238002 214708 238008
rect 214668 237930 214696 238002
rect 214656 237924 214708 237930
rect 214656 237866 214708 237872
rect 214760 236570 214788 307158
rect 214852 236609 214880 309703
rect 214944 237114 214972 309878
rect 214932 237108 214984 237114
rect 214932 237050 214984 237056
rect 215036 237046 215064 315250
rect 215128 237182 215156 316639
rect 217782 316568 217838 316577
rect 217782 316503 217838 316512
rect 217692 315376 217744 315382
rect 217598 315344 217654 315353
rect 217692 315318 217744 315324
rect 217598 315279 217654 315288
rect 216218 314256 216274 314265
rect 216218 314191 216274 314200
rect 216036 312724 216088 312730
rect 216036 312666 216088 312672
rect 215944 312588 215996 312594
rect 215944 312530 215996 312536
rect 215760 310004 215812 310010
rect 215760 309946 215812 309952
rect 215206 309904 215262 309913
rect 215206 309839 215262 309848
rect 215116 237176 215168 237182
rect 215116 237118 215168 237124
rect 215024 237040 215076 237046
rect 215024 236982 215076 236988
rect 214838 236600 214894 236609
rect 214748 236564 214800 236570
rect 214838 236535 214894 236544
rect 214748 236506 214800 236512
rect 214656 236020 214708 236026
rect 214656 235962 214708 235968
rect 214668 228478 214696 235962
rect 214852 229945 214880 236535
rect 215128 236026 215156 237118
rect 215116 236020 215168 236026
rect 215116 235962 215168 235968
rect 214838 229936 214894 229945
rect 214838 229871 214894 229880
rect 214656 228472 214708 228478
rect 214656 228414 214708 228420
rect 215220 224913 215248 309839
rect 215772 241534 215800 309946
rect 215852 307148 215904 307154
rect 215852 307090 215904 307096
rect 215760 241528 215812 241534
rect 215760 241470 215812 241476
rect 215576 240372 215628 240378
rect 215576 240314 215628 240320
rect 215588 239494 215616 240314
rect 215666 240272 215722 240281
rect 215666 240207 215722 240216
rect 215576 239488 215628 239494
rect 215576 239430 215628 239436
rect 215576 239080 215628 239086
rect 215576 239022 215628 239028
rect 215300 237380 215352 237386
rect 215300 237322 215352 237328
rect 214746 224904 214802 224913
rect 214746 224839 214802 224848
rect 215206 224904 215262 224913
rect 215206 224839 215262 224848
rect 214760 224233 214788 224839
rect 214746 224224 214802 224233
rect 214746 224159 214802 224168
rect 215312 164898 215340 237322
rect 215300 164892 215352 164898
rect 215300 164834 215352 164840
rect 214564 18624 214616 18630
rect 214564 18566 214616 18572
rect 213932 16546 214512 16574
rect 213276 4072 213328 4078
rect 213276 4014 213328 4020
rect 213184 3596 213236 3602
rect 213184 3538 213236 3544
rect 213104 3454 213408 3482
rect 213380 480 213408 3454
rect 214484 480 214512 16546
rect 215588 3942 215616 239022
rect 215680 231169 215708 240207
rect 215758 240000 215814 240009
rect 215758 239935 215814 239944
rect 215772 239057 215800 239935
rect 215758 239048 215814 239057
rect 215758 238983 215814 238992
rect 215864 236978 215892 307090
rect 215956 241097 215984 312530
rect 215942 241088 215998 241097
rect 215942 241023 215998 241032
rect 215956 240281 215984 241023
rect 215942 240272 215998 240281
rect 215942 240207 215998 240216
rect 215944 239556 215996 239562
rect 215944 239498 215996 239504
rect 215852 236972 215904 236978
rect 215852 236914 215904 236920
rect 215666 231160 215722 231169
rect 215666 231095 215722 231104
rect 215956 4010 215984 239498
rect 216048 239290 216076 312666
rect 216128 312656 216180 312662
rect 216128 312598 216180 312604
rect 216036 239284 216088 239290
rect 216036 239226 216088 239232
rect 216140 239154 216168 312598
rect 216232 240242 216260 314191
rect 216494 314120 216550 314129
rect 216494 314055 216550 314064
rect 216312 314016 216364 314022
rect 216312 313958 216364 313964
rect 216220 240236 216272 240242
rect 216220 240178 216272 240184
rect 216128 239148 216180 239154
rect 216128 239090 216180 239096
rect 216126 239048 216182 239057
rect 216126 238983 216182 238992
rect 216140 234614 216168 238983
rect 216232 237017 216260 240178
rect 216324 240009 216352 313958
rect 216404 313948 216456 313954
rect 216404 313890 216456 313896
rect 216310 240000 216366 240009
rect 216310 239935 216366 239944
rect 216312 239896 216364 239902
rect 216312 239838 216364 239844
rect 216218 237008 216274 237017
rect 216218 236943 216274 236952
rect 216324 236842 216352 239838
rect 216416 237998 216444 313890
rect 216404 237992 216456 237998
rect 216404 237934 216456 237940
rect 216508 237289 216536 314055
rect 216586 313984 216642 313993
rect 216586 313919 216642 313928
rect 216600 239902 216628 313919
rect 217508 311908 217560 311914
rect 217508 311850 217560 311856
rect 217416 309256 217468 309262
rect 217416 309198 217468 309204
rect 217324 307352 217376 307358
rect 217324 307294 217376 307300
rect 217232 291848 217284 291854
rect 217232 291790 217284 291796
rect 217138 240680 217194 240689
rect 217138 240615 217194 240624
rect 216588 239896 216640 239902
rect 216588 239838 216640 239844
rect 216588 239284 216640 239290
rect 216588 239226 216640 239232
rect 216600 239018 216628 239226
rect 216588 239012 216640 239018
rect 216588 238954 216640 238960
rect 216586 238096 216642 238105
rect 216586 238031 216642 238040
rect 216600 237386 216628 238031
rect 216588 237380 216640 237386
rect 216588 237322 216640 237328
rect 216494 237280 216550 237289
rect 216494 237215 216550 237224
rect 216312 236836 216364 236842
rect 216312 236778 216364 236784
rect 216140 234586 216352 234614
rect 216324 219434 216352 234586
rect 217152 232529 217180 240615
rect 217244 239426 217272 291790
rect 217232 239420 217284 239426
rect 217232 239362 217284 239368
rect 217336 238785 217364 307294
rect 217428 240281 217456 309198
rect 217520 240961 217548 311850
rect 217506 240952 217562 240961
rect 217506 240887 217562 240896
rect 217520 240689 217548 240887
rect 217506 240680 217562 240689
rect 217506 240615 217562 240624
rect 217612 240417 217640 315279
rect 217598 240408 217654 240417
rect 217598 240343 217654 240352
rect 217414 240272 217470 240281
rect 217414 240207 217470 240216
rect 217322 238776 217378 238785
rect 217322 238711 217378 238720
rect 217428 238626 217456 240207
rect 217244 238598 217456 238626
rect 217138 232520 217194 232529
rect 217138 232455 217194 232464
rect 217244 229809 217272 238598
rect 217416 238060 217468 238066
rect 217416 238002 217468 238008
rect 217322 235648 217378 235657
rect 217322 235583 217378 235592
rect 217230 229800 217286 229809
rect 217230 229735 217286 229744
rect 216678 226944 216734 226953
rect 216678 226879 216734 226888
rect 216140 219406 216352 219434
rect 216140 4146 216168 219406
rect 216692 16574 216720 226879
rect 216692 16546 216904 16574
rect 216128 4140 216180 4146
rect 216128 4082 216180 4088
rect 215944 4004 215996 4010
rect 215944 3946 215996 3952
rect 215576 3936 215628 3942
rect 215576 3878 215628 3884
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 215680 480 215708 3470
rect 216876 480 216904 16546
rect 217336 3466 217364 235583
rect 217428 17270 217456 238002
rect 217612 231441 217640 240343
rect 217704 240310 217732 315318
rect 217692 240304 217744 240310
rect 217692 240246 217744 240252
rect 217796 238882 217824 316503
rect 217874 314528 217930 314537
rect 217874 314463 217930 314472
rect 217784 238876 217836 238882
rect 217784 238818 217836 238824
rect 217888 236910 217916 314463
rect 217980 239630 218008 321943
rect 220634 321736 220690 321745
rect 220634 321671 220690 321680
rect 219164 320340 219216 320346
rect 219164 320282 219216 320288
rect 218980 318164 219032 318170
rect 218980 318106 219032 318112
rect 218796 316804 218848 316810
rect 218796 316746 218848 316752
rect 218612 309868 218664 309874
rect 218612 309810 218664 309816
rect 217968 239624 218020 239630
rect 217968 239566 218020 239572
rect 217876 236904 217928 236910
rect 217876 236846 217928 236852
rect 217598 231432 217654 231441
rect 217598 231367 217654 231376
rect 217888 228410 217916 236846
rect 218624 235754 218652 309810
rect 218704 304428 218756 304434
rect 218704 304370 218756 304376
rect 218716 240689 218744 304370
rect 218808 240990 218836 316746
rect 218888 314084 218940 314090
rect 218888 314026 218940 314032
rect 218796 240984 218848 240990
rect 218796 240926 218848 240932
rect 218808 240786 218836 240926
rect 218796 240780 218848 240786
rect 218796 240722 218848 240728
rect 218702 240680 218758 240689
rect 218702 240615 218758 240624
rect 218716 240514 218744 240615
rect 218704 240508 218756 240514
rect 218704 240450 218756 240456
rect 218704 239420 218756 239426
rect 218704 239362 218756 239368
rect 218612 235748 218664 235754
rect 218612 235690 218664 235696
rect 218060 234048 218112 234054
rect 218060 233990 218112 233996
rect 217876 228404 217928 228410
rect 217876 228346 217928 228352
rect 217416 17264 217468 17270
rect 217416 17206 217468 17212
rect 217324 3460 217376 3466
rect 217324 3402 217376 3408
rect 218072 480 218100 233990
rect 218152 230036 218204 230042
rect 218152 229978 218204 229984
rect 218164 16574 218192 229978
rect 218164 16546 218652 16574
rect 218624 3482 218652 16546
rect 218716 3806 218744 239362
rect 218900 237017 218928 314026
rect 218992 239698 219020 318106
rect 219072 318096 219124 318102
rect 219072 318038 219124 318044
rect 218980 239692 219032 239698
rect 218980 239634 219032 239640
rect 219084 239426 219112 318038
rect 219176 240514 219204 320282
rect 219348 320204 219400 320210
rect 219348 320146 219400 320152
rect 219254 316976 219310 316985
rect 219254 316911 219310 316920
rect 219268 240650 219296 316911
rect 219256 240644 219308 240650
rect 219256 240586 219308 240592
rect 219164 240508 219216 240514
rect 219164 240450 219216 240456
rect 219176 240134 219204 240450
rect 219360 240394 219388 320146
rect 220544 314152 220596 314158
rect 220544 314094 220596 314100
rect 220450 312488 220506 312497
rect 220450 312423 220506 312432
rect 220360 307080 220412 307086
rect 220360 307022 220412 307028
rect 220268 304360 220320 304366
rect 220268 304302 220320 304308
rect 220176 304292 220228 304298
rect 220176 304234 220228 304240
rect 220084 292596 220136 292602
rect 220084 292538 220136 292544
rect 219900 291372 219952 291378
rect 219900 291314 219952 291320
rect 219912 253230 219940 291314
rect 219992 290148 220044 290154
rect 219992 290090 220044 290096
rect 219900 253224 219952 253230
rect 219900 253166 219952 253172
rect 220004 241466 220032 290090
rect 219992 241460 220044 241466
rect 219992 241402 220044 241408
rect 220096 241346 220124 292538
rect 220004 241318 220124 241346
rect 219360 240366 219480 240394
rect 219176 240106 219388 240134
rect 219348 240100 219400 240106
rect 219348 240042 219400 240048
rect 219452 239986 219480 240366
rect 219360 239958 219480 239986
rect 219360 239902 219388 239958
rect 219164 239896 219216 239902
rect 219164 239838 219216 239844
rect 219348 239896 219400 239902
rect 219348 239838 219400 239844
rect 219176 239766 219204 239838
rect 219164 239760 219216 239766
rect 219164 239702 219216 239708
rect 219256 239760 219308 239766
rect 219256 239702 219308 239708
rect 219072 239420 219124 239426
rect 219072 239362 219124 239368
rect 219084 239222 219112 239362
rect 219072 239216 219124 239222
rect 219072 239158 219124 239164
rect 219176 239057 219204 239702
rect 219162 239048 219218 239057
rect 219162 238983 219218 238992
rect 219268 237833 219296 239702
rect 219348 239692 219400 239698
rect 219348 239634 219400 239640
rect 219360 239426 219388 239634
rect 219348 239420 219400 239426
rect 219348 239362 219400 239368
rect 219438 238232 219494 238241
rect 219438 238167 219494 238176
rect 219254 237824 219310 237833
rect 219254 237759 219310 237768
rect 218980 237652 219032 237658
rect 218980 237594 219032 237600
rect 218886 237008 218942 237017
rect 218886 236943 218942 236952
rect 218900 234614 218928 236943
rect 218808 234586 218928 234614
rect 218704 3800 218756 3806
rect 218704 3742 218756 3748
rect 218808 3738 218836 234586
rect 218992 169046 219020 237594
rect 218980 169040 219032 169046
rect 218980 168982 219032 168988
rect 219452 16574 219480 238167
rect 220004 237969 220032 241318
rect 220082 241224 220138 241233
rect 220082 241159 220138 241168
rect 220096 240553 220124 241159
rect 220188 240854 220216 304234
rect 220176 240848 220228 240854
rect 220176 240790 220228 240796
rect 220082 240544 220138 240553
rect 220082 240479 220138 240488
rect 220280 239834 220308 304302
rect 220372 241058 220400 307022
rect 220360 241052 220412 241058
rect 220360 240994 220412 241000
rect 220372 240922 220400 240994
rect 220360 240916 220412 240922
rect 220360 240858 220412 240864
rect 220358 240544 220414 240553
rect 220358 240479 220414 240488
rect 220372 240281 220400 240479
rect 220358 240272 220414 240281
rect 220358 240207 220414 240216
rect 220268 239828 220320 239834
rect 220268 239770 220320 239776
rect 220280 239290 220308 239770
rect 220268 239284 220320 239290
rect 220268 239226 220320 239232
rect 220360 238808 220412 238814
rect 220360 238750 220412 238756
rect 220268 238332 220320 238338
rect 220268 238274 220320 238280
rect 219990 237960 220046 237969
rect 219990 237895 220046 237904
rect 220004 234614 220032 237895
rect 220176 237720 220228 237726
rect 220176 237662 220228 237668
rect 220004 234586 220124 234614
rect 220096 232762 220124 234586
rect 220084 232756 220136 232762
rect 220084 232698 220136 232704
rect 220188 171834 220216 237662
rect 220280 175982 220308 238274
rect 220268 175976 220320 175982
rect 220268 175918 220320 175924
rect 220176 171828 220228 171834
rect 220176 171770 220228 171776
rect 219452 16546 220032 16574
rect 218796 3732 218848 3738
rect 218796 3674 218848 3680
rect 218624 3454 219296 3482
rect 219268 480 219296 3454
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220372 3874 220400 238750
rect 220464 238241 220492 312423
rect 220450 238232 220506 238241
rect 220450 238167 220506 238176
rect 220556 236706 220584 314094
rect 220648 239494 220676 321671
rect 220740 239601 220768 322079
rect 221922 318744 221978 318753
rect 221922 318679 221978 318688
rect 221740 317756 221792 317762
rect 221740 317698 221792 317704
rect 221648 311160 221700 311166
rect 221648 311102 221700 311108
rect 221556 301504 221608 301510
rect 221556 301446 221608 301452
rect 221464 298784 221516 298790
rect 221464 298726 221516 298732
rect 220912 291440 220964 291446
rect 220912 291382 220964 291388
rect 220924 286346 220952 291382
rect 220912 286340 220964 286346
rect 220912 286282 220964 286288
rect 221004 241528 221056 241534
rect 221004 241470 221056 241476
rect 220820 240644 220872 240650
rect 220820 240586 220872 240592
rect 220726 239592 220782 239601
rect 220726 239527 220782 239536
rect 220636 239488 220688 239494
rect 220636 239430 220688 239436
rect 220544 236700 220596 236706
rect 220544 236642 220596 236648
rect 220740 236298 220768 239527
rect 220832 237590 220860 240586
rect 220910 240272 220966 240281
rect 220910 240207 220966 240216
rect 220820 237584 220872 237590
rect 220820 237526 220872 237532
rect 220924 236570 220952 240207
rect 221016 239902 221044 241470
rect 221372 240780 221424 240786
rect 221372 240722 221424 240728
rect 221188 240508 221240 240514
rect 221188 240450 221240 240456
rect 221096 240304 221148 240310
rect 221096 240246 221148 240252
rect 221004 239896 221056 239902
rect 221004 239838 221056 239844
rect 221016 237318 221044 239838
rect 221108 237794 221136 240246
rect 221200 238649 221228 240450
rect 221280 239828 221332 239834
rect 221280 239770 221332 239776
rect 221186 238640 221242 238649
rect 221186 238575 221242 238584
rect 221188 238468 221240 238474
rect 221188 238410 221240 238416
rect 221200 238270 221228 238410
rect 221292 238270 221320 239770
rect 221384 238610 221412 240722
rect 221372 238604 221424 238610
rect 221372 238546 221424 238552
rect 221188 238264 221240 238270
rect 221188 238206 221240 238212
rect 221280 238264 221332 238270
rect 221280 238206 221332 238212
rect 221476 237862 221504 298726
rect 221568 238678 221596 301446
rect 221660 238950 221688 311102
rect 221752 240718 221780 317698
rect 221832 313880 221884 313886
rect 221832 313822 221884 313828
rect 221844 240786 221872 313822
rect 221832 240780 221884 240786
rect 221832 240722 221884 240728
rect 221740 240712 221792 240718
rect 221740 240654 221792 240660
rect 221740 240236 221792 240242
rect 221740 240178 221792 240184
rect 221648 238944 221700 238950
rect 221648 238886 221700 238892
rect 221556 238672 221608 238678
rect 221556 238614 221608 238620
rect 221752 238406 221780 240178
rect 221936 239970 221964 318679
rect 222200 307284 222252 307290
rect 222200 307226 222252 307232
rect 222016 291304 222068 291310
rect 222016 291246 222068 291252
rect 221924 239964 221976 239970
rect 221924 239906 221976 239912
rect 221740 238400 221792 238406
rect 221740 238342 221792 238348
rect 221648 238128 221700 238134
rect 221648 238070 221700 238076
rect 221464 237856 221516 237862
rect 221464 237798 221516 237804
rect 221096 237788 221148 237794
rect 221096 237730 221148 237736
rect 221004 237312 221056 237318
rect 221004 237254 221056 237260
rect 220912 236564 220964 236570
rect 220912 236506 220964 236512
rect 220728 236292 220780 236298
rect 220728 236234 220780 236240
rect 220820 235816 220872 235822
rect 220820 235758 220872 235764
rect 220832 16574 220860 235758
rect 221660 207670 221688 238070
rect 221936 229770 221964 239906
rect 221924 229764 221976 229770
rect 221924 229706 221976 229712
rect 221648 207664 221700 207670
rect 221648 207606 221700 207612
rect 222028 126274 222056 291246
rect 222108 291236 222160 291242
rect 222108 291178 222160 291184
rect 222016 126268 222068 126274
rect 222016 126210 222068 126216
rect 222120 87650 222148 291178
rect 222212 240106 222240 307226
rect 222292 295996 222344 296002
rect 222292 295938 222344 295944
rect 222304 241369 222332 295938
rect 223776 293078 223804 360198
rect 223948 293344 224000 293350
rect 223948 293286 224000 293292
rect 223764 293072 223816 293078
rect 223764 293014 223816 293020
rect 223960 292602 223988 293286
rect 223948 292596 224000 292602
rect 223948 292538 224000 292544
rect 223960 289884 223988 292538
rect 224236 291242 224264 363559
rect 225602 362264 225658 362273
rect 225602 362199 225658 362208
rect 225234 329080 225290 329089
rect 225234 329015 225290 329024
rect 225052 322244 225104 322250
rect 225052 322186 225104 322192
rect 224868 319728 224920 319734
rect 224868 319670 224920 319676
rect 224592 311500 224644 311506
rect 224592 311442 224644 311448
rect 224500 293072 224552 293078
rect 224500 293014 224552 293020
rect 224224 291236 224276 291242
rect 224224 291178 224276 291184
rect 224236 289898 224264 291178
rect 224512 289898 224540 293014
rect 224604 290057 224632 311442
rect 224590 290048 224646 290057
rect 224590 289983 224646 289992
rect 224236 289870 224342 289898
rect 224512 289870 224710 289898
rect 224880 289626 224908 319670
rect 225064 293078 225092 322186
rect 225248 306374 225276 329015
rect 225248 306346 225552 306374
rect 225052 293072 225104 293078
rect 225052 293014 225104 293020
rect 225052 291576 225104 291582
rect 225052 291518 225104 291524
rect 225064 289884 225092 291518
rect 225420 291236 225472 291242
rect 225420 291178 225472 291184
rect 225432 289884 225460 291178
rect 225524 290068 225552 306346
rect 225616 291242 225644 362199
rect 226340 358828 226392 358834
rect 226340 358770 226392 358776
rect 226352 293078 226380 358770
rect 226430 320784 226486 320793
rect 226430 320719 226486 320728
rect 225972 293072 226024 293078
rect 225972 293014 226024 293020
rect 226340 293072 226392 293078
rect 226340 293014 226392 293020
rect 225604 291236 225656 291242
rect 225604 291178 225656 291184
rect 225524 290040 225644 290068
rect 225616 289898 225644 290040
rect 225984 289898 226012 293014
rect 226444 291145 226472 320719
rect 226892 296744 226944 296750
rect 226892 296686 226944 296692
rect 226524 291508 226576 291514
rect 226524 291450 226576 291456
rect 226430 291136 226486 291145
rect 226430 291071 226486 291080
rect 225616 289870 225814 289898
rect 225984 289870 226182 289898
rect 226536 289884 226564 291450
rect 226904 289884 226932 296686
rect 226996 291582 227024 367503
rect 227732 306374 227760 367639
rect 227732 306346 227852 306374
rect 227076 293072 227128 293078
rect 227076 293014 227128 293020
rect 226984 291576 227036 291582
rect 226984 291518 227036 291524
rect 227088 289898 227116 293014
rect 227626 291136 227682 291145
rect 227626 291071 227682 291080
rect 227640 289921 227668 291071
rect 227626 289912 227682 289921
rect 227088 289870 227286 289898
rect 227824 289898 227852 306346
rect 228364 293480 228416 293486
rect 228364 293422 228416 293428
rect 227824 289870 228022 289898
rect 228376 289884 228404 293422
rect 228730 291544 228786 291553
rect 228730 291479 228786 291488
rect 228744 289884 228772 291479
rect 229112 289884 229140 372982
rect 229192 370660 229244 370666
rect 229192 370602 229244 370608
rect 229204 296714 229232 370602
rect 229284 369164 229336 369170
rect 229284 369106 229336 369112
rect 229296 306374 229324 369106
rect 229296 306346 230060 306374
rect 229468 298852 229520 298858
rect 229468 298794 229520 298800
rect 229204 296686 229324 296714
rect 229296 290086 229324 296686
rect 229284 290080 229336 290086
rect 229284 290022 229336 290028
rect 229480 289884 229508 298794
rect 229744 290080 229796 290086
rect 229744 290022 229796 290028
rect 229756 289898 229784 290022
rect 230032 289898 230060 306346
rect 230492 293078 230520 373322
rect 234632 373318 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299584 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700330 283880 703520
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 250444 514820 250496 514826
rect 250444 514762 250496 514768
rect 250456 406434 250484 514762
rect 250444 406428 250496 406434
rect 250444 406370 250496 406376
rect 255320 391264 255372 391270
rect 255320 391206 255372 391212
rect 255332 390590 255360 391206
rect 255320 390584 255372 390590
rect 255320 390526 255372 390532
rect 245660 383036 245712 383042
rect 245660 382978 245712 382984
rect 236644 375828 236696 375834
rect 236644 375770 236696 375776
rect 236000 375420 236052 375426
rect 236000 375362 236052 375368
rect 234712 374196 234764 374202
rect 234712 374138 234764 374144
rect 234620 373312 234672 373318
rect 234620 373254 234672 373260
rect 231122 371648 231178 371657
rect 231122 371583 231178 371592
rect 230572 327752 230624 327758
rect 230572 327694 230624 327700
rect 230480 293072 230532 293078
rect 230480 293014 230532 293020
rect 229756 289870 229862 289898
rect 230032 289870 230230 289898
rect 230584 289884 230612 327694
rect 231136 296750 231164 371583
rect 231952 370524 232004 370530
rect 231952 370466 232004 370472
rect 231860 370388 231912 370394
rect 231860 370330 231912 370336
rect 231124 296744 231176 296750
rect 231124 296686 231176 296692
rect 231676 293548 231728 293554
rect 231676 293490 231728 293496
rect 231124 293072 231176 293078
rect 231124 293014 231176 293020
rect 230940 291236 230992 291242
rect 230940 291178 230992 291184
rect 230952 289884 230980 291178
rect 231136 289898 231164 293014
rect 231136 289870 231334 289898
rect 231688 289884 231716 293490
rect 231872 292074 231900 370330
rect 231964 306374 231992 370466
rect 233240 368552 233292 368558
rect 233240 368494 233292 368500
rect 233056 315444 233108 315450
rect 233056 315386 233108 315392
rect 231964 306346 232636 306374
rect 231872 292046 232176 292074
rect 232044 291984 232096 291990
rect 232044 291926 232096 291932
rect 232056 289884 232084 291926
rect 232148 290170 232176 292046
rect 232228 291576 232280 291582
rect 232228 291518 232280 291524
rect 232240 290494 232268 291518
rect 232228 290488 232280 290494
rect 232228 290430 232280 290436
rect 232148 290142 232268 290170
rect 232240 289898 232268 290142
rect 232608 289898 232636 306346
rect 232964 297424 233016 297430
rect 232964 297366 233016 297372
rect 232240 289870 232438 289898
rect 232608 289870 232806 289898
rect 227626 289847 227682 289856
rect 224958 289640 225014 289649
rect 224880 289598 224958 289626
rect 232976 289626 233004 297366
rect 233068 289785 233096 315386
rect 233252 306374 233280 368494
rect 233252 306346 233372 306374
rect 233344 289898 233372 306346
rect 234724 296714 234752 374138
rect 235632 312860 235684 312866
rect 235632 312802 235684 312808
rect 234632 296686 234752 296714
rect 233884 293616 233936 293622
rect 233884 293558 233936 293564
rect 233344 289870 233542 289898
rect 233896 289884 233924 293558
rect 234252 292052 234304 292058
rect 234252 291994 234304 292000
rect 234264 289884 234292 291994
rect 234632 289884 234660 296686
rect 234988 292188 235040 292194
rect 234988 292130 235040 292136
rect 235000 289884 235028 292130
rect 235356 291916 235408 291922
rect 235356 291858 235408 291864
rect 235368 289884 235396 291858
rect 235644 289785 235672 312802
rect 235908 312792 235960 312798
rect 235908 312734 235960 312740
rect 235724 294636 235776 294642
rect 235724 294578 235776 294584
rect 235736 289884 235764 294578
rect 233054 289776 233110 289785
rect 233054 289711 233110 289720
rect 235630 289776 235686 289785
rect 235630 289711 235686 289720
rect 235920 289649 235948 312734
rect 236012 293078 236040 375362
rect 236092 370592 236144 370598
rect 236092 370534 236144 370540
rect 236104 306374 236132 370534
rect 236104 306346 236500 306374
rect 236092 293412 236144 293418
rect 236092 293354 236144 293360
rect 236000 293072 236052 293078
rect 236000 293014 236052 293020
rect 236104 289884 236132 293354
rect 236368 292120 236420 292126
rect 236368 292062 236420 292068
rect 236380 289898 236408 292062
rect 236472 290170 236500 306346
rect 236656 296714 236684 375770
rect 239404 375692 239456 375698
rect 239404 375634 239456 375640
rect 238760 375556 238812 375562
rect 238760 375498 238812 375504
rect 237378 370016 237434 370025
rect 237378 369951 237434 369960
rect 236564 296686 236684 296714
rect 236564 292194 236592 296686
rect 237012 293072 237064 293078
rect 237012 293014 237064 293020
rect 236552 292188 236604 292194
rect 236552 292130 236604 292136
rect 236472 290142 236684 290170
rect 236656 289898 236684 290142
rect 237024 289898 237052 293014
rect 237392 292074 237420 369951
rect 237472 319456 237524 319462
rect 237472 319398 237524 319404
rect 237484 306374 237512 319398
rect 237484 306346 238524 306374
rect 238300 292528 238352 292534
rect 238300 292470 238352 292476
rect 237392 292046 237788 292074
rect 237564 291984 237616 291990
rect 237564 291926 237616 291932
rect 236380 289870 236486 289898
rect 236656 289870 236854 289898
rect 237024 289870 237222 289898
rect 237576 289884 237604 291926
rect 237760 289898 237788 292046
rect 237760 289870 237958 289898
rect 238312 289884 238340 292470
rect 238496 289898 238524 306346
rect 238666 306368 238722 306377
rect 238772 306374 238800 375498
rect 238852 318436 238904 318442
rect 238852 318378 238904 318384
rect 238864 315489 238892 318378
rect 238850 315480 238906 315489
rect 238850 315415 238906 315424
rect 238772 306346 239260 306374
rect 238666 306303 238722 306312
rect 238680 296857 238708 306303
rect 238666 296848 238722 296857
rect 238666 296783 238722 296792
rect 238666 296712 238722 296721
rect 238666 296647 238722 296656
rect 238680 290329 238708 296647
rect 239034 293176 239090 293185
rect 239034 293111 239090 293120
rect 238666 290320 238722 290329
rect 238666 290255 238722 290264
rect 238496 289870 238694 289898
rect 239048 289884 239076 293111
rect 239232 289898 239260 306346
rect 239416 292534 239444 375634
rect 244280 375624 244332 375630
rect 244280 375566 244332 375572
rect 240140 375488 240192 375494
rect 240140 375430 240192 375436
rect 240152 301578 240180 375430
rect 243544 372088 243596 372094
rect 243544 372030 243596 372036
rect 242164 371272 242216 371278
rect 242164 371214 242216 371220
rect 241520 370796 241572 370802
rect 241520 370738 241572 370744
rect 240414 370424 240470 370433
rect 240414 370359 240470 370368
rect 240230 370152 240286 370161
rect 240230 370087 240286 370096
rect 240140 301572 240192 301578
rect 240140 301514 240192 301520
rect 240244 296714 240272 370087
rect 240428 306374 240456 370359
rect 240428 306346 241100 306374
rect 240324 301572 240376 301578
rect 240324 301514 240376 301520
rect 240152 296686 240272 296714
rect 239404 292528 239456 292534
rect 239404 292470 239456 292476
rect 239772 290692 239824 290698
rect 239772 290634 239824 290640
rect 239232 289870 239430 289898
rect 239784 289884 239812 290634
rect 240152 289884 240180 296686
rect 240336 289898 240364 301514
rect 240876 290624 240928 290630
rect 240876 290566 240928 290572
rect 240336 289870 240534 289898
rect 240888 289884 240916 290566
rect 241072 289898 241100 306346
rect 241532 293078 241560 370738
rect 241610 320648 241666 320657
rect 241610 320583 241666 320592
rect 241624 306374 241652 320583
rect 241624 306346 241836 306374
rect 241610 293312 241666 293321
rect 241610 293247 241666 293256
rect 241520 293072 241572 293078
rect 241520 293014 241572 293020
rect 241072 289870 241270 289898
rect 241624 289884 241652 293247
rect 241808 289898 241836 306346
rect 242176 298858 242204 371214
rect 242900 370320 242952 370326
rect 242900 370262 242952 370268
rect 242164 298852 242216 298858
rect 242164 298794 242216 298800
rect 242714 294808 242770 294817
rect 242714 294743 242770 294752
rect 242164 293072 242216 293078
rect 242164 293014 242216 293020
rect 242176 289898 242204 293014
rect 241808 289870 242006 289898
rect 242176 289870 242374 289898
rect 242728 289884 242756 294743
rect 242912 293078 242940 370262
rect 242990 321056 243046 321065
rect 242990 320991 243046 321000
rect 242900 293072 242952 293078
rect 242900 293014 242952 293020
rect 243004 293010 243032 320991
rect 243084 319320 243136 319326
rect 243084 319262 243136 319268
rect 242992 293004 243044 293010
rect 242992 292946 243044 292952
rect 243096 289884 243124 319262
rect 243556 293486 243584 372030
rect 244292 296154 244320 375566
rect 245016 372156 245068 372162
rect 245016 372098 245068 372104
rect 244924 370456 244976 370462
rect 244924 370398 244976 370404
rect 244370 319424 244426 319433
rect 244370 319359 244426 319368
rect 244384 306374 244412 319359
rect 244384 306346 244872 306374
rect 244292 296126 244780 296154
rect 244556 296064 244608 296070
rect 244556 296006 244608 296012
rect 243544 293480 243596 293486
rect 243544 293422 243596 293428
rect 243268 293072 243320 293078
rect 243268 293014 243320 293020
rect 243280 289898 243308 293014
rect 244004 293004 244056 293010
rect 244004 292946 244056 292952
rect 243820 290488 243872 290494
rect 243820 290430 243872 290436
rect 243280 289870 243478 289898
rect 243832 289884 243860 290430
rect 244016 289898 244044 292946
rect 244016 289870 244214 289898
rect 244568 289884 244596 296006
rect 244752 289898 244780 296126
rect 244844 290170 244872 306346
rect 244936 292194 244964 370398
rect 245028 293554 245056 372098
rect 245016 293548 245068 293554
rect 245016 293490 245068 293496
rect 244924 292188 244976 292194
rect 244924 292130 244976 292136
rect 244844 290142 245148 290170
rect 245120 289898 245148 290142
rect 244752 289870 244950 289898
rect 245120 289870 245318 289898
rect 245672 289884 245700 382978
rect 249800 375760 249852 375766
rect 249800 375702 249852 375708
rect 248420 373312 248472 373318
rect 248420 373254 248472 373260
rect 245752 372224 245804 372230
rect 245752 372166 245804 372172
rect 245764 301866 245792 372166
rect 247684 371544 247736 371550
rect 247684 371486 247736 371492
rect 245844 370252 245896 370258
rect 245844 370194 245896 370200
rect 245856 301986 245884 370194
rect 247040 370184 247092 370190
rect 247040 370126 247092 370132
rect 245936 369232 245988 369238
rect 245936 369174 245988 369180
rect 245948 306374 245976 369174
rect 245948 306346 246252 306374
rect 245844 301980 245896 301986
rect 245844 301922 245896 301928
rect 245764 301838 245976 301866
rect 245752 301776 245804 301782
rect 245752 301718 245804 301724
rect 245764 293078 245792 301718
rect 245948 296714 245976 301838
rect 245856 296686 245976 296714
rect 245752 293072 245804 293078
rect 245752 293014 245804 293020
rect 245856 289898 245884 296686
rect 246224 289898 246252 306346
rect 247052 293078 247080 370126
rect 247130 321328 247186 321337
rect 247130 321263 247186 321272
rect 247144 306374 247172 321263
rect 247224 318504 247276 318510
rect 247224 318446 247276 318452
rect 247236 314673 247264 318446
rect 247222 314664 247278 314673
rect 247222 314599 247278 314608
rect 247144 306346 247356 306374
rect 247132 304496 247184 304502
rect 247132 304438 247184 304444
rect 246580 293072 246632 293078
rect 246580 293014 246632 293020
rect 247040 293072 247092 293078
rect 247040 293014 247092 293020
rect 246592 289898 246620 293014
rect 245856 289870 246054 289898
rect 246224 289870 246422 289898
rect 246592 289870 246790 289898
rect 247144 289884 247172 304438
rect 247328 289898 247356 306346
rect 247696 296714 247724 371486
rect 248432 369238 248460 373254
rect 248420 369232 248472 369238
rect 248420 369174 248472 369180
rect 248418 321192 248474 321201
rect 248418 321127 248474 321136
rect 247604 296686 247724 296714
rect 247604 293622 247632 296686
rect 248236 293956 248288 293962
rect 248236 293898 248288 293904
rect 247592 293616 247644 293622
rect 247592 293558 247644 293564
rect 247684 293072 247736 293078
rect 247684 293014 247736 293020
rect 247696 289898 247724 293014
rect 247328 289870 247526 289898
rect 247696 289870 247894 289898
rect 248248 289884 248276 293898
rect 248432 289898 248460 321127
rect 248512 320476 248564 320482
rect 248512 320418 248564 320424
rect 248524 290170 248552 320418
rect 248696 319252 248748 319258
rect 248696 319194 248748 319200
rect 248604 319184 248656 319190
rect 248604 319126 248656 319132
rect 248616 292574 248644 319126
rect 248708 306374 248736 319194
rect 249616 311364 249668 311370
rect 249616 311306 249668 311312
rect 248708 306346 249564 306374
rect 248616 292546 249196 292574
rect 248524 290142 248828 290170
rect 248800 289898 248828 290142
rect 249168 289898 249196 292546
rect 249536 289898 249564 306346
rect 249628 290057 249656 311306
rect 249812 293078 249840 375702
rect 253204 374604 253256 374610
rect 253204 374546 253256 374552
rect 251178 374096 251234 374105
rect 251178 374031 251234 374040
rect 250444 371476 250496 371482
rect 250444 371418 250496 371424
rect 249890 368656 249946 368665
rect 249890 368591 249946 368600
rect 249800 293072 249852 293078
rect 249800 293014 249852 293020
rect 249614 290048 249670 290057
rect 249614 289983 249670 289992
rect 249904 289898 249932 368591
rect 249984 320408 250036 320414
rect 249984 320350 250036 320356
rect 249996 306374 250024 320350
rect 249996 306346 250392 306374
rect 250260 293072 250312 293078
rect 250260 293014 250312 293020
rect 250272 289898 250300 293014
rect 250364 292574 250392 306346
rect 250456 293962 250484 371418
rect 251088 311432 251140 311438
rect 251088 311374 251140 311380
rect 250996 311296 251048 311302
rect 250996 311238 251048 311244
rect 250720 311228 250772 311234
rect 250720 311170 250772 311176
rect 250444 293956 250496 293962
rect 250444 293898 250496 293904
rect 250364 292546 250668 292574
rect 250640 289898 250668 292546
rect 250732 290057 250760 311170
rect 250718 290048 250774 290057
rect 250718 289983 250774 289992
rect 248432 289870 248630 289898
rect 248800 289870 248998 289898
rect 249168 289870 249366 289898
rect 249536 289870 249734 289898
rect 249904 289870 250102 289898
rect 250272 289870 250470 289898
rect 250640 289870 250838 289898
rect 249248 289672 249300 289678
rect 235906 289640 235962 289649
rect 232976 289598 233174 289626
rect 224958 289575 225014 289584
rect 251008 289649 251036 311238
rect 251100 289785 251128 311374
rect 251192 289884 251220 374031
rect 251270 368928 251326 368937
rect 251270 368863 251326 368872
rect 251284 293078 251312 368863
rect 251362 367840 251418 367849
rect 251362 367775 251418 367784
rect 251272 293072 251324 293078
rect 251272 293014 251324 293020
rect 251376 289898 251404 367775
rect 252560 356720 252612 356726
rect 252560 356662 252612 356668
rect 251456 319388 251508 319394
rect 251456 319330 251508 319336
rect 251468 306374 251496 319330
rect 252468 312928 252520 312934
rect 252468 312870 252520 312876
rect 251468 306346 251772 306374
rect 251744 289898 251772 306346
rect 252100 293072 252152 293078
rect 252100 293014 252152 293020
rect 252112 289898 252140 293014
rect 251376 289870 251574 289898
rect 251744 289870 251942 289898
rect 252112 289870 252310 289898
rect 251086 289776 251142 289785
rect 251086 289711 251142 289720
rect 249248 289614 249300 289620
rect 250994 289640 251050 289649
rect 235906 289575 235962 289584
rect 249260 289542 249288 289614
rect 252480 289626 252508 312870
rect 252572 293010 252600 356662
rect 252650 320920 252706 320929
rect 252650 320855 252706 320864
rect 252664 293078 252692 320855
rect 252744 319524 252796 319530
rect 252744 319466 252796 319472
rect 252756 306374 252784 319466
rect 252756 306346 252876 306374
rect 252652 293072 252704 293078
rect 252652 293014 252704 293020
rect 252560 293004 252612 293010
rect 252560 292946 252612 292952
rect 252650 292088 252706 292097
rect 252650 292023 252706 292032
rect 252664 289884 252692 292023
rect 252848 289898 252876 306346
rect 253112 305040 253164 305046
rect 253112 304982 253164 304988
rect 253124 301782 253152 304982
rect 253112 301776 253164 301782
rect 253112 301718 253164 301724
rect 253216 296714 253244 374546
rect 253938 369064 253994 369073
rect 253938 368999 253994 369008
rect 253952 298926 253980 368999
rect 254122 368792 254178 368801
rect 254122 368727 254178 368736
rect 254030 320512 254086 320521
rect 254030 320447 254086 320456
rect 253940 298920 253992 298926
rect 253940 298862 253992 298868
rect 253124 296686 253244 296714
rect 253124 292126 253152 296686
rect 253204 293072 253256 293078
rect 253204 293014 253256 293020
rect 253112 292120 253164 292126
rect 253112 292062 253164 292068
rect 253216 289898 253244 293014
rect 253572 293004 253624 293010
rect 253572 292946 253624 292952
rect 253584 289898 253612 292946
rect 254044 289898 254072 320447
rect 254136 290306 254164 368727
rect 254214 319560 254270 319569
rect 254214 319495 254270 319504
rect 254228 306374 254256 319495
rect 254228 306346 255084 306374
rect 254676 298920 254728 298926
rect 254676 298862 254728 298868
rect 254136 290278 254348 290306
rect 254320 289898 254348 290278
rect 254688 289898 254716 298862
rect 255056 289898 255084 306346
rect 255332 292574 255360 390526
rect 266372 383042 266400 697546
rect 289084 632120 289136 632126
rect 289084 632062 289136 632068
rect 266360 383036 266412 383042
rect 266360 382978 266412 382984
rect 262128 376780 262180 376786
rect 262128 376722 262180 376728
rect 255964 374468 256016 374474
rect 255964 374410 256016 374416
rect 255412 369300 255464 369306
rect 255412 369242 255464 369248
rect 255424 297362 255452 369242
rect 255504 323604 255556 323610
rect 255504 323546 255556 323552
rect 255516 306374 255544 323546
rect 255516 306346 255820 306374
rect 255412 297356 255464 297362
rect 255412 297298 255464 297304
rect 255332 292546 255452 292574
rect 255424 289898 255452 292546
rect 255792 289898 255820 306346
rect 255976 290698 256004 374410
rect 257344 374400 257396 374406
rect 257344 374342 257396 374348
rect 256700 372632 256752 372638
rect 256700 372574 256752 372580
rect 256516 310208 256568 310214
rect 256516 310150 256568 310156
rect 256240 310072 256292 310078
rect 256240 310014 256292 310020
rect 256148 291508 256200 291514
rect 256148 291450 256200 291456
rect 255964 290692 256016 290698
rect 255964 290634 256016 290640
rect 252848 289870 253046 289898
rect 253216 289870 253414 289898
rect 253584 289870 253782 289898
rect 254044 289870 254150 289898
rect 254320 289870 254518 289898
rect 254688 289870 254886 289898
rect 255056 289870 255254 289898
rect 255424 289870 255622 289898
rect 255792 289870 255990 289898
rect 256160 289814 256188 291450
rect 256148 289808 256200 289814
rect 256252 289785 256280 310014
rect 256332 297356 256384 297362
rect 256332 297298 256384 297304
rect 256344 289884 256372 297298
rect 256528 290057 256556 310150
rect 256608 310140 256660 310146
rect 256608 310082 256660 310088
rect 256514 290048 256570 290057
rect 256514 289983 256570 289992
rect 256516 289808 256568 289814
rect 256148 289750 256200 289756
rect 256238 289776 256294 289785
rect 256238 289711 256294 289720
rect 256514 289776 256516 289785
rect 256568 289776 256570 289785
rect 256514 289711 256570 289720
rect 256620 289649 256648 310082
rect 256712 297498 256740 372574
rect 256790 345672 256846 345681
rect 256790 345607 256846 345616
rect 256804 345098 256832 345607
rect 256792 345092 256844 345098
rect 256792 345034 256844 345040
rect 256804 299538 256832 345034
rect 256884 324964 256936 324970
rect 256884 324906 256936 324912
rect 256792 299532 256844 299538
rect 256792 299474 256844 299480
rect 256700 297492 256752 297498
rect 256700 297434 256752 297440
rect 256896 297362 256924 324906
rect 256974 319696 257030 319705
rect 256974 319631 257030 319640
rect 256884 297356 256936 297362
rect 256884 297298 256936 297304
rect 256988 289762 257016 319631
rect 257252 297492 257304 297498
rect 257252 297434 257304 297440
rect 257068 297356 257120 297362
rect 257068 297298 257120 297304
rect 257080 289884 257108 297298
rect 257264 289898 257292 297434
rect 257356 290630 257384 374342
rect 259644 374332 259696 374338
rect 259644 374274 259696 374280
rect 258816 373176 258868 373182
rect 258816 373118 258868 373124
rect 257436 373108 257488 373114
rect 257436 373050 257488 373056
rect 257448 372638 257476 373050
rect 258724 372972 258776 372978
rect 258724 372914 258776 372920
rect 257436 372632 257488 372638
rect 257436 372574 257488 372580
rect 258356 364404 258408 364410
rect 258356 364346 258408 364352
rect 258368 358086 258396 364346
rect 258356 358080 258408 358086
rect 258356 358022 258408 358028
rect 258172 318776 258224 318782
rect 258172 318718 258224 318724
rect 257620 299532 257672 299538
rect 257620 299474 257672 299480
rect 257344 290624 257396 290630
rect 257344 290566 257396 290572
rect 257632 289898 257660 299474
rect 258184 294710 258212 318718
rect 258368 299474 258396 358022
rect 258276 299446 258396 299474
rect 258172 294704 258224 294710
rect 258172 294646 258224 294652
rect 258276 294522 258304 299446
rect 258540 294704 258592 294710
rect 258540 294646 258592 294652
rect 258184 294494 258304 294522
rect 257264 289870 257462 289898
rect 257632 289870 257830 289898
rect 258184 289884 258212 294494
rect 258552 289884 258580 294646
rect 258736 293282 258764 372914
rect 258828 318782 258856 373118
rect 259552 372836 259604 372842
rect 259552 372778 259604 372784
rect 258816 318776 258868 318782
rect 258816 318718 258868 318724
rect 258816 301776 258868 301782
rect 258816 301718 258868 301724
rect 258828 300830 258856 301718
rect 258816 300824 258868 300830
rect 258816 300766 258868 300772
rect 259092 300824 259144 300830
rect 259092 300766 259144 300772
rect 258724 293276 258776 293282
rect 258724 293218 258776 293224
rect 258736 292574 258764 293218
rect 258736 292546 258948 292574
rect 258920 289884 258948 292546
rect 259104 289898 259132 300766
rect 259104 289870 259302 289898
rect 259564 289814 259592 372778
rect 259656 306374 259684 374274
rect 260104 374128 260156 374134
rect 260104 374070 260156 374076
rect 259656 306346 259868 306374
rect 259644 292528 259696 292534
rect 259644 292470 259696 292476
rect 259656 291582 259684 292470
rect 259644 291576 259696 291582
rect 259644 291518 259696 291524
rect 259656 289884 259684 291518
rect 259840 290154 259868 306346
rect 260116 291446 260144 374070
rect 261024 372768 261076 372774
rect 261024 372710 261076 372716
rect 260196 370728 260248 370734
rect 260196 370670 260248 370676
rect 260208 292534 260236 370670
rect 260930 319832 260986 319841
rect 260930 319767 260986 319776
rect 260288 305720 260340 305726
rect 260288 305662 260340 305668
rect 260196 292528 260248 292534
rect 260196 292470 260248 292476
rect 260300 292058 260328 305662
rect 260288 292052 260340 292058
rect 260288 291994 260340 292000
rect 260104 291440 260156 291446
rect 260104 291382 260156 291388
rect 260116 290170 260144 291382
rect 259828 290148 259880 290154
rect 260116 290142 260236 290170
rect 259828 290090 259880 290096
rect 259840 289898 259868 290090
rect 260208 289898 260236 290142
rect 260944 290018 260972 319767
rect 261036 306374 261064 372710
rect 261484 326392 261536 326398
rect 261484 326334 261536 326340
rect 261036 306346 261340 306374
rect 260932 290012 260984 290018
rect 260932 289954 260984 289960
rect 260944 289898 260972 289954
rect 259840 289870 260038 289898
rect 260208 289870 260406 289898
rect 260944 289870 261142 289898
rect 261312 289814 261340 306346
rect 261496 291378 261524 326334
rect 262140 292534 262168 376722
rect 275100 375896 275152 375902
rect 275100 375838 275152 375844
rect 262496 374944 262548 374950
rect 262496 374886 262548 374892
rect 262404 373244 262456 373250
rect 262404 373186 262456 373192
rect 262312 372904 262364 372910
rect 262312 372846 262364 372852
rect 262128 292528 262180 292534
rect 262128 292470 262180 292476
rect 262324 291786 262352 372846
rect 262312 291780 262364 291786
rect 262312 291722 262364 291728
rect 261484 291372 261536 291378
rect 261484 291314 261536 291320
rect 261496 289884 261524 291314
rect 262128 289944 262180 289950
rect 262416 289898 262444 373186
rect 262508 290154 262536 374886
rect 264888 374264 264940 374270
rect 264888 374206 264940 374212
rect 263598 372872 263654 372881
rect 263598 372807 263654 372816
rect 263612 306374 263640 372807
rect 264244 366376 264296 366382
rect 264244 366318 264296 366324
rect 263612 306346 263916 306374
rect 262588 292528 262640 292534
rect 262588 292470 262640 292476
rect 262600 291854 262628 292470
rect 263692 292052 263744 292058
rect 263692 291994 263744 292000
rect 262588 291848 262640 291854
rect 262588 291790 262640 291796
rect 262496 290148 262548 290154
rect 262496 290090 262548 290096
rect 262180 289892 262444 289898
rect 262128 289886 262444 289892
rect 262140 289870 262444 289886
rect 262508 289882 262536 290090
rect 262600 289884 262628 291790
rect 262772 291780 262824 291786
rect 262772 291722 262824 291728
rect 262784 289898 262812 291722
rect 263704 291718 263732 291994
rect 263692 291712 263744 291718
rect 263692 291654 263744 291660
rect 263324 290148 263376 290154
rect 263324 290090 263376 290096
rect 262496 289876 262548 289882
rect 262496 289818 262548 289824
rect 262784 289870 262982 289898
rect 263336 289884 263364 290090
rect 263704 289884 263732 291654
rect 263888 289898 263916 306346
rect 264256 292534 264284 366318
rect 264336 319592 264388 319598
rect 264336 319534 264388 319540
rect 264244 292528 264296 292534
rect 264244 292470 264296 292476
rect 264348 291417 264376 319534
rect 264796 292528 264848 292534
rect 264796 292470 264848 292476
rect 264808 291650 264836 292470
rect 264796 291644 264848 291650
rect 264796 291586 264848 291592
rect 264334 291408 264390 291417
rect 264334 291343 264390 291352
rect 264348 289898 264376 291343
rect 263888 289870 264086 289898
rect 264348 289870 264454 289898
rect 264808 289884 264836 291586
rect 264900 290902 264928 374206
rect 264978 372736 265034 372745
rect 264978 372671 265034 372680
rect 264888 290896 264940 290902
rect 264888 290838 264940 290844
rect 264900 290562 264928 290838
rect 264888 290556 264940 290562
rect 264888 290498 264940 290504
rect 256726 289734 257016 289762
rect 259552 289808 259604 289814
rect 259552 289750 259604 289756
rect 260564 289808 260616 289814
rect 261300 289808 261352 289814
rect 260616 289756 260774 289762
rect 260564 289750 260774 289756
rect 261300 289750 261352 289756
rect 261668 289808 261720 289814
rect 261720 289756 261878 289762
rect 261668 289750 261878 289756
rect 252558 289640 252614 289649
rect 252480 289598 252558 289626
rect 250994 289575 251050 289584
rect 252558 289575 252614 289584
rect 256606 289640 256662 289649
rect 256606 289575 256662 289584
rect 259564 289542 259592 289750
rect 260576 289734 260774 289750
rect 261312 289542 261340 289750
rect 261680 289734 261878 289750
rect 262784 289610 262812 289870
rect 263888 289649 263916 289870
rect 264992 289649 265020 372671
rect 272616 320544 272668 320550
rect 272616 320486 272668 320492
rect 269764 319660 269816 319666
rect 269764 319602 269816 319608
rect 268384 315580 268436 315586
rect 268384 315522 268436 315528
rect 265900 291848 265952 291854
rect 265900 291790 265952 291796
rect 265912 291281 265940 291790
rect 265898 291272 265954 291281
rect 265898 291207 265954 291216
rect 265532 290896 265584 290902
rect 265532 290838 265584 290844
rect 265544 289884 265572 290838
rect 265912 289884 265940 291207
rect 263874 289640 263930 289649
rect 262772 289604 262824 289610
rect 263874 289575 263930 289584
rect 264978 289640 265034 289649
rect 264978 289575 265034 289584
rect 262772 289546 262824 289552
rect 249248 289536 249300 289542
rect 249248 289478 249300 289484
rect 259552 289536 259604 289542
rect 259552 289478 259604 289484
rect 261300 289536 261352 289542
rect 261300 289478 261352 289484
rect 265162 289368 265218 289377
rect 265162 289303 265218 289312
rect 222476 289196 222528 289202
rect 222476 289138 222528 289144
rect 222488 288862 222516 289138
rect 222476 288856 222528 288862
rect 222476 288798 222528 288804
rect 267554 272504 267610 272513
rect 267554 272439 267610 272448
rect 267568 244225 267596 272439
rect 267646 250472 267702 250481
rect 267646 250407 267702 250416
rect 267554 244216 267610 244225
rect 267554 244151 267610 244160
rect 267554 244080 267610 244089
rect 267554 244015 267610 244024
rect 267568 241641 267596 244015
rect 267554 241632 267610 241641
rect 267554 241567 267610 241576
rect 222290 241360 222346 241369
rect 222290 241295 222346 241304
rect 267464 241324 267516 241330
rect 267464 241266 267516 241272
rect 267476 241233 267504 241266
rect 267660 241262 267688 250407
rect 267922 246256 267978 246265
rect 267922 246191 267978 246200
rect 267830 243536 267886 243545
rect 267830 243471 267886 243480
rect 267648 241256 267700 241262
rect 267462 241224 267518 241233
rect 267648 241198 267700 241204
rect 267462 241159 267518 241168
rect 267740 241188 267792 241194
rect 267740 241130 267792 241136
rect 267556 241120 267608 241126
rect 267648 241120 267700 241126
rect 267556 241062 267608 241068
rect 267646 241088 267648 241097
rect 267700 241088 267702 241097
rect 222292 240916 222344 240922
rect 222292 240858 222344 240864
rect 222304 240650 222332 240858
rect 267568 240718 267596 241062
rect 267646 241023 267702 241032
rect 267752 240990 267780 241130
rect 267740 240984 267792 240990
rect 267740 240926 267792 240932
rect 267740 240848 267792 240854
rect 267740 240790 267792 240796
rect 267556 240712 267608 240718
rect 267556 240654 267608 240660
rect 267752 240650 267780 240790
rect 222292 240644 222344 240650
rect 222292 240586 222344 240592
rect 267740 240644 267792 240650
rect 267740 240586 267792 240592
rect 267740 240372 267792 240378
rect 267740 240314 267792 240320
rect 222292 240304 222344 240310
rect 222290 240272 222292 240281
rect 222344 240272 222346 240281
rect 222290 240207 222346 240216
rect 222290 240136 222346 240145
rect 222200 240100 222252 240106
rect 267752 240122 267780 240314
rect 222290 240071 222346 240080
rect 222200 240042 222252 240048
rect 222212 239850 222240 240042
rect 222304 240038 222332 240071
rect 222292 240032 222344 240038
rect 222292 239974 222344 239980
rect 222384 239964 222436 239970
rect 222534 239952 222562 240108
rect 222436 239924 222562 239952
rect 222384 239906 222436 239912
rect 222212 239822 222516 239850
rect 222200 239760 222252 239766
rect 222200 239702 222252 239708
rect 222212 239193 222240 239702
rect 222292 239624 222344 239630
rect 222292 239566 222344 239572
rect 222198 239184 222254 239193
rect 222198 239119 222254 239128
rect 222304 229094 222332 239566
rect 222382 236328 222438 236337
rect 222382 236263 222438 236272
rect 222212 229066 222332 229094
rect 222212 215966 222240 229066
rect 222396 220794 222424 236263
rect 222384 220788 222436 220794
rect 222384 220730 222436 220736
rect 222200 215960 222252 215966
rect 222200 215902 222252 215908
rect 222200 181552 222252 181558
rect 222200 181494 222252 181500
rect 222108 87644 222160 87650
rect 222108 87586 222160 87592
rect 222212 16574 222240 181494
rect 222488 174554 222516 239822
rect 222626 239465 222654 240108
rect 222718 239902 222746 240108
rect 222810 239902 222838 240108
rect 222902 239970 222930 240108
rect 222890 239964 222942 239970
rect 222890 239906 222942 239912
rect 222706 239896 222758 239902
rect 222706 239838 222758 239844
rect 222798 239896 222850 239902
rect 222798 239838 222850 239844
rect 222752 239760 222804 239766
rect 222750 239728 222752 239737
rect 222804 239728 222806 239737
rect 222750 239663 222806 239672
rect 222994 239544 223022 240108
rect 223086 239907 223114 240108
rect 223072 239898 223128 239907
rect 223178 239902 223206 240108
rect 223072 239833 223128 239842
rect 223166 239896 223218 239902
rect 223166 239838 223218 239844
rect 223270 239748 223298 240108
rect 223362 239970 223390 240108
rect 223454 239970 223482 240108
rect 223350 239964 223402 239970
rect 223350 239906 223402 239912
rect 223442 239964 223494 239970
rect 223442 239906 223494 239912
rect 223546 239834 223574 240108
rect 223638 239850 223666 240108
rect 223730 239970 223758 240108
rect 223718 239964 223770 239970
rect 223718 239906 223770 239912
rect 223534 239828 223586 239834
rect 223638 239822 223712 239850
rect 223534 239770 223586 239776
rect 223118 239728 223174 239737
rect 223118 239663 223120 239672
rect 223172 239663 223174 239672
rect 223224 239720 223298 239748
rect 223394 239728 223450 239737
rect 223120 239634 223172 239640
rect 222764 239516 223022 239544
rect 222612 239456 222668 239465
rect 222612 239391 222668 239400
rect 222764 237794 222792 239516
rect 222934 239456 222990 239465
rect 222934 239391 222990 239400
rect 222842 239320 222898 239329
rect 222842 239255 222898 239264
rect 222856 238921 222884 239255
rect 222842 238912 222898 238921
rect 222842 238847 222898 238856
rect 222842 237824 222898 237833
rect 222752 237788 222804 237794
rect 222842 237759 222898 237768
rect 222752 237730 222804 237736
rect 222568 237380 222620 237386
rect 222568 237322 222620 237328
rect 222580 181490 222608 237322
rect 222660 237244 222712 237250
rect 222660 237186 222712 237192
rect 222672 189786 222700 237186
rect 222764 202162 222792 237730
rect 222752 202156 222804 202162
rect 222752 202098 222804 202104
rect 222660 189780 222712 189786
rect 222660 189722 222712 189728
rect 222568 181484 222620 181490
rect 222568 181426 222620 181432
rect 222476 174548 222528 174554
rect 222476 174490 222528 174496
rect 222856 22778 222884 237759
rect 222948 227050 222976 239391
rect 223132 237386 223160 239634
rect 223224 239193 223252 239720
rect 223394 239663 223396 239672
rect 223448 239663 223450 239672
rect 223580 239692 223632 239698
rect 223396 239634 223448 239640
rect 223580 239634 223632 239640
rect 223302 239456 223358 239465
rect 223302 239391 223358 239400
rect 223210 239184 223266 239193
rect 223210 239119 223266 239128
rect 223316 237658 223344 239391
rect 223304 237652 223356 237658
rect 223304 237594 223356 237600
rect 223120 237380 223172 237386
rect 223120 237322 223172 237328
rect 223028 237312 223080 237318
rect 223028 237254 223080 237260
rect 222936 227044 222988 227050
rect 222936 226986 222988 226992
rect 222936 220788 222988 220794
rect 222936 220730 222988 220736
rect 222948 220250 222976 220730
rect 222936 220244 222988 220250
rect 222936 220186 222988 220192
rect 222948 203590 222976 220186
rect 223040 210458 223068 237254
rect 223408 237250 223436 239634
rect 223488 239624 223540 239630
rect 223592 239601 223620 239634
rect 223488 239566 223540 239572
rect 223578 239592 223634 239601
rect 223500 238513 223528 239566
rect 223578 239527 223634 239536
rect 223486 238504 223542 238513
rect 223486 238439 223542 238448
rect 223684 237833 223712 239822
rect 223822 239816 223850 240108
rect 223914 239902 223942 240108
rect 224006 239902 224034 240108
rect 223902 239896 223954 239902
rect 223902 239838 223954 239844
rect 223994 239896 224046 239902
rect 223994 239838 224046 239844
rect 223776 239788 223850 239816
rect 223670 237824 223726 237833
rect 223670 237759 223726 237768
rect 223396 237244 223448 237250
rect 223396 237186 223448 237192
rect 223672 236564 223724 236570
rect 223776 236552 223804 239788
rect 223854 239728 223910 239737
rect 224098 239680 224126 240108
rect 224190 239907 224218 240108
rect 224176 239898 224232 239907
rect 224282 239902 224310 240108
rect 224374 239902 224402 240108
rect 224176 239833 224232 239842
rect 224270 239896 224322 239902
rect 224270 239838 224322 239844
rect 224362 239896 224414 239902
rect 224362 239838 224414 239844
rect 224316 239760 224368 239766
rect 223854 239663 223856 239672
rect 223908 239663 223910 239672
rect 223856 239634 223908 239640
rect 224052 239652 224126 239680
rect 224314 239728 224316 239737
rect 224466 239748 224494 240108
rect 224558 239970 224586 240108
rect 224650 239970 224678 240108
rect 224742 239970 224770 240108
rect 224834 239970 224862 240108
rect 224546 239964 224598 239970
rect 224546 239906 224598 239912
rect 224638 239964 224690 239970
rect 224638 239906 224690 239912
rect 224730 239964 224782 239970
rect 224730 239906 224782 239912
rect 224822 239964 224874 239970
rect 224822 239906 224874 239912
rect 224592 239828 224644 239834
rect 224592 239770 224644 239776
rect 224730 239828 224782 239834
rect 224926 239816 224954 240108
rect 225018 239970 225046 240108
rect 225006 239964 225058 239970
rect 225006 239906 225058 239912
rect 225110 239850 225138 240108
rect 225202 239873 225230 240108
rect 225294 239970 225322 240108
rect 225386 239970 225414 240108
rect 225282 239964 225334 239970
rect 225282 239906 225334 239912
rect 225374 239964 225426 239970
rect 225374 239906 225426 239912
rect 225064 239822 225138 239850
rect 225188 239864 225244 239873
rect 224926 239788 225000 239816
rect 224730 239770 224782 239776
rect 224368 239728 224370 239737
rect 224314 239663 224370 239672
rect 224420 239720 224494 239748
rect 223946 239592 224002 239601
rect 223946 239527 224002 239536
rect 223960 238202 223988 239527
rect 223948 238196 224000 238202
rect 223948 238138 224000 238144
rect 223776 236524 223896 236552
rect 223672 236506 223724 236512
rect 223580 236292 223632 236298
rect 223580 236234 223632 236240
rect 223592 224262 223620 236234
rect 223580 224256 223632 224262
rect 223580 224198 223632 224204
rect 223028 210452 223080 210458
rect 223028 210394 223080 210400
rect 222936 203584 222988 203590
rect 222936 203526 222988 203532
rect 223684 184210 223712 236506
rect 223762 236328 223818 236337
rect 223762 236263 223818 236272
rect 223776 220833 223804 236263
rect 223868 221814 223896 236524
rect 224052 235793 224080 239652
rect 224224 239624 224276 239630
rect 224144 239584 224224 239612
rect 224144 237590 224172 239584
rect 224224 239566 224276 239572
rect 224328 238474 224356 239663
rect 224316 238468 224368 238474
rect 224316 238410 224368 238416
rect 224420 237912 224448 239720
rect 224500 239624 224552 239630
rect 224604 239601 224632 239770
rect 224742 239714 224770 239770
rect 224972 239748 225000 239788
rect 224696 239686 224770 239714
rect 224880 239720 225000 239748
rect 224500 239566 224552 239572
rect 224590 239592 224646 239601
rect 224512 238377 224540 239566
rect 224590 239527 224646 239536
rect 224590 238640 224646 238649
rect 224590 238575 224646 238584
rect 224604 238474 224632 238575
rect 224592 238468 224644 238474
rect 224592 238410 224644 238416
rect 224498 238368 224554 238377
rect 224498 238303 224554 238312
rect 224328 237884 224448 237912
rect 224132 237584 224184 237590
rect 224132 237526 224184 237532
rect 224038 235784 224094 235793
rect 224038 235719 224094 235728
rect 224144 235634 224172 237526
rect 224224 236360 224276 236366
rect 224224 236302 224276 236308
rect 223960 235606 224172 235634
rect 223856 221808 223908 221814
rect 223856 221750 223908 221756
rect 223762 220824 223818 220833
rect 223762 220759 223818 220768
rect 223960 199442 223988 235606
rect 224040 235204 224092 235210
rect 224040 235146 224092 235152
rect 224052 219337 224080 235146
rect 224132 221808 224184 221814
rect 224132 221750 224184 221756
rect 224144 221474 224172 221750
rect 224132 221468 224184 221474
rect 224132 221410 224184 221416
rect 224236 219434 224264 236302
rect 224144 219406 224264 219434
rect 224038 219328 224094 219337
rect 224038 219263 224094 219272
rect 224052 213246 224080 219263
rect 224040 213240 224092 213246
rect 224040 213182 224092 213188
rect 223948 199436 224000 199442
rect 223948 199378 224000 199384
rect 223672 184204 223724 184210
rect 223672 184146 223724 184152
rect 222844 22772 222896 22778
rect 222844 22714 222896 22720
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 220360 3868 220412 3874
rect 220360 3810 220412 3816
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 224144 13122 224172 219406
rect 224328 219298 224356 237884
rect 224408 237788 224460 237794
rect 224408 237730 224460 237736
rect 224316 219292 224368 219298
rect 224316 219234 224368 219240
rect 224328 217326 224356 219234
rect 224316 217320 224368 217326
rect 224316 217262 224368 217268
rect 224316 215348 224368 215354
rect 224316 215290 224368 215296
rect 224132 13116 224184 13122
rect 224132 13058 224184 13064
rect 224328 11762 224356 215290
rect 224420 167686 224448 237730
rect 224512 236366 224540 238303
rect 224592 236972 224644 236978
rect 224592 236914 224644 236920
rect 224500 236360 224552 236366
rect 224500 236302 224552 236308
rect 224604 236201 224632 236914
rect 224590 236192 224646 236201
rect 224590 236127 224646 236136
rect 224696 235210 224724 239686
rect 224776 239624 224828 239630
rect 224776 239566 224828 239572
rect 224788 237318 224816 239566
rect 224880 237794 224908 239720
rect 224868 237788 224920 237794
rect 224868 237730 224920 237736
rect 224880 237697 224908 237730
rect 224866 237688 224922 237697
rect 224866 237623 224922 237632
rect 224960 237652 225012 237658
rect 224960 237594 225012 237600
rect 224868 237584 224920 237590
rect 224868 237526 224920 237532
rect 224776 237312 224828 237318
rect 224776 237254 224828 237260
rect 224684 235204 224736 235210
rect 224684 235146 224736 235152
rect 224498 220824 224554 220833
rect 224498 220759 224554 220768
rect 224512 220561 224540 220759
rect 224498 220552 224554 220561
rect 224498 220487 224554 220496
rect 224512 209098 224540 220487
rect 224880 216510 224908 237526
rect 224972 237046 225000 237594
rect 224960 237040 225012 237046
rect 224960 236982 225012 236988
rect 224972 236348 225000 236982
rect 225064 236473 225092 239822
rect 225478 239816 225506 240108
rect 225570 239970 225598 240108
rect 225662 239970 225690 240108
rect 225558 239964 225610 239970
rect 225558 239906 225610 239912
rect 225650 239964 225702 239970
rect 225650 239906 225702 239912
rect 225188 239799 225244 239808
rect 225432 239788 225506 239816
rect 225604 239828 225656 239834
rect 225144 239760 225196 239766
rect 225144 239702 225196 239708
rect 225156 237658 225184 239702
rect 225236 239692 225288 239698
rect 225236 239634 225288 239640
rect 225248 239306 225276 239634
rect 225328 239624 225380 239630
rect 225326 239592 225328 239601
rect 225380 239592 225382 239601
rect 225326 239527 225382 239536
rect 225248 239278 225368 239306
rect 225236 238536 225288 238542
rect 225236 238478 225288 238484
rect 225144 237652 225196 237658
rect 225144 237594 225196 237600
rect 225248 237368 225276 238478
rect 225340 237436 225368 239278
rect 225432 237590 225460 239788
rect 225754 239816 225782 240108
rect 225604 239770 225656 239776
rect 225708 239788 225782 239816
rect 225512 239624 225564 239630
rect 225512 239566 225564 239572
rect 225524 239057 225552 239566
rect 225510 239048 225566 239057
rect 225510 238983 225566 238992
rect 225420 237584 225472 237590
rect 225420 237526 225472 237532
rect 225340 237408 225460 237436
rect 225248 237340 225368 237368
rect 225144 237312 225196 237318
rect 225144 237254 225196 237260
rect 225050 236464 225106 236473
rect 225050 236399 225106 236408
rect 224972 236320 225092 236348
rect 224958 236192 225014 236201
rect 224958 236127 225014 236136
rect 224868 216504 224920 216510
rect 224868 216446 224920 216452
rect 224880 215354 224908 216446
rect 224972 216034 225000 236127
rect 225064 222902 225092 236320
rect 225052 222896 225104 222902
rect 225052 222838 225104 222844
rect 225052 216164 225104 216170
rect 225052 216106 225104 216112
rect 224960 216028 225012 216034
rect 224960 215970 225012 215976
rect 224868 215348 224920 215354
rect 224868 215290 224920 215296
rect 224500 209092 224552 209098
rect 224500 209034 224552 209040
rect 224408 167680 224460 167686
rect 224408 167622 224460 167628
rect 225064 16574 225092 216106
rect 225156 193866 225184 237254
rect 225236 231532 225288 231538
rect 225236 231474 225288 231480
rect 225248 220697 225276 231474
rect 225234 220688 225290 220697
rect 225234 220623 225290 220632
rect 225248 214606 225276 220623
rect 225236 214600 225288 214606
rect 225236 214542 225288 214548
rect 225144 193860 225196 193866
rect 225144 193802 225196 193808
rect 225340 180130 225368 237340
rect 225432 237114 225460 237408
rect 225420 237108 225472 237114
rect 225420 237050 225472 237056
rect 225432 218754 225460 237050
rect 225420 218748 225472 218754
rect 225420 218690 225472 218696
rect 225524 211818 225552 238983
rect 225616 238950 225644 239770
rect 225604 238944 225656 238950
rect 225604 238886 225656 238892
rect 225616 229094 225644 238886
rect 225708 238746 225736 239788
rect 225846 239680 225874 240108
rect 225938 239748 225966 240108
rect 226030 239873 226058 240108
rect 226122 239902 226150 240108
rect 226214 239970 226242 240108
rect 226202 239964 226254 239970
rect 226202 239906 226254 239912
rect 226110 239896 226162 239902
rect 226016 239864 226072 239873
rect 226110 239838 226162 239844
rect 226016 239799 226072 239808
rect 225938 239737 226104 239748
rect 225938 239728 226118 239737
rect 225938 239720 226062 239728
rect 225846 239652 225966 239680
rect 226306 239680 226334 240108
rect 226398 239873 226426 240108
rect 226384 239864 226440 239873
rect 226384 239799 226440 239808
rect 226490 239748 226518 240108
rect 226582 239902 226610 240108
rect 226674 239902 226702 240108
rect 226766 239902 226794 240108
rect 226570 239896 226622 239902
rect 226570 239838 226622 239844
rect 226662 239896 226714 239902
rect 226662 239838 226714 239844
rect 226754 239896 226806 239902
rect 226754 239838 226806 239844
rect 226858 239850 226886 240108
rect 226950 239970 226978 240108
rect 227042 239970 227070 240108
rect 226938 239964 226990 239970
rect 226938 239906 226990 239912
rect 227030 239964 227082 239970
rect 227030 239906 227082 239912
rect 227134 239873 227162 240108
rect 227226 239902 227254 240108
rect 227318 239907 227346 240108
rect 227410 239970 227438 240108
rect 227398 239964 227450 239970
rect 227214 239896 227266 239902
rect 226982 239864 227038 239873
rect 226858 239822 226982 239850
rect 226982 239799 227038 239808
rect 227120 239864 227176 239873
rect 227214 239838 227266 239844
rect 227304 239898 227360 239907
rect 227398 239906 227450 239912
rect 227502 239902 227530 240108
rect 227594 239902 227622 240108
rect 227686 239907 227714 240108
rect 227778 239970 227806 240108
rect 227766 239964 227818 239970
rect 227304 239833 227360 239842
rect 227490 239896 227542 239902
rect 227490 239838 227542 239844
rect 227582 239896 227634 239902
rect 227582 239838 227634 239844
rect 227672 239898 227728 239907
rect 227766 239906 227818 239912
rect 227672 239833 227728 239842
rect 227120 239799 227176 239808
rect 226062 239663 226118 239672
rect 225938 239578 225966 239652
rect 226260 239652 226334 239680
rect 226444 239720 226518 239748
rect 226892 239760 226944 239766
rect 226706 239728 226762 239737
rect 225892 239550 225966 239578
rect 226064 239624 226116 239630
rect 226064 239566 226116 239572
rect 225696 238740 225748 238746
rect 225696 238682 225748 238688
rect 225892 235929 225920 239550
rect 225972 238740 226024 238746
rect 225972 238682 226024 238688
rect 225984 238270 226012 238682
rect 225972 238264 226024 238270
rect 225972 238206 226024 238212
rect 226076 237946 226104 239566
rect 226260 238542 226288 239652
rect 226340 238876 226392 238882
rect 226340 238818 226392 238824
rect 226248 238536 226300 238542
rect 226154 238504 226210 238513
rect 226248 238478 226300 238484
rect 226154 238439 226210 238448
rect 225984 237918 226104 237946
rect 225984 236910 226012 237918
rect 226064 237788 226116 237794
rect 226064 237730 226116 237736
rect 225972 236904 226024 236910
rect 225972 236846 226024 236852
rect 225878 235920 225934 235929
rect 225878 235855 225934 235864
rect 226076 231538 226104 237730
rect 226168 237658 226196 238439
rect 226156 237652 226208 237658
rect 226156 237594 226208 237600
rect 226168 235550 226196 237594
rect 226248 237312 226300 237318
rect 226248 237254 226300 237260
rect 226260 236706 226288 237254
rect 226248 236700 226300 236706
rect 226248 236642 226300 236648
rect 226156 235544 226208 235550
rect 226156 235486 226208 235492
rect 226064 231532 226116 231538
rect 226064 231474 226116 231480
rect 225616 229066 225828 229094
rect 225512 211812 225564 211818
rect 225512 211754 225564 211760
rect 225800 192506 225828 229066
rect 226352 224330 226380 238818
rect 226444 230654 226472 239720
rect 226616 239692 226668 239698
rect 226890 239728 226892 239737
rect 227122 239760 227174 239766
rect 226944 239728 226946 239737
rect 226706 239663 226762 239672
rect 226800 239692 226852 239698
rect 226616 239634 226668 239640
rect 226628 238610 226656 239634
rect 226720 239630 226748 239663
rect 226890 239663 226946 239672
rect 226996 239720 227122 239748
rect 226800 239634 226852 239640
rect 226708 239624 226760 239630
rect 226708 239566 226760 239572
rect 226812 238785 226840 239634
rect 226892 239624 226944 239630
rect 226892 239566 226944 239572
rect 226798 238776 226854 238785
rect 226720 238734 226798 238762
rect 226616 238604 226668 238610
rect 226616 238546 226668 238552
rect 226522 238504 226578 238513
rect 226522 238439 226578 238448
rect 226432 230648 226484 230654
rect 226432 230590 226484 230596
rect 226536 227186 226564 238439
rect 226628 238270 226656 238546
rect 226616 238264 226668 238270
rect 226616 238206 226668 238212
rect 226614 238096 226670 238105
rect 226614 238031 226670 238040
rect 226628 233730 226656 238031
rect 226720 233866 226748 238734
rect 226798 238711 226854 238720
rect 226798 238232 226854 238241
rect 226798 238167 226854 238176
rect 226812 235278 226840 238167
rect 226904 236638 226932 239566
rect 226996 237794 227024 239720
rect 227122 239702 227174 239708
rect 227536 239760 227588 239766
rect 227870 239748 227898 240108
rect 227962 239873 227990 240108
rect 228054 239902 228082 240108
rect 228146 239970 228174 240108
rect 228134 239964 228186 239970
rect 228134 239906 228186 239912
rect 228238 239902 228266 240108
rect 228042 239896 228094 239902
rect 227948 239864 228004 239873
rect 228042 239838 228094 239844
rect 228226 239896 228278 239902
rect 228226 239838 228278 239844
rect 227948 239799 228004 239808
rect 228330 239748 228358 240108
rect 227536 239702 227588 239708
rect 227626 239728 227682 239737
rect 227352 239692 227404 239698
rect 227352 239634 227404 239640
rect 227258 239592 227314 239601
rect 227076 239556 227128 239562
rect 227076 239498 227128 239504
rect 227168 239556 227220 239562
rect 227258 239527 227260 239536
rect 227168 239498 227220 239504
rect 227312 239527 227314 239536
rect 227260 239498 227312 239504
rect 227088 238542 227116 239498
rect 227180 238882 227208 239498
rect 227168 238876 227220 238882
rect 227168 238818 227220 238824
rect 227076 238536 227128 238542
rect 227076 238478 227128 238484
rect 227260 238196 227312 238202
rect 227260 238138 227312 238144
rect 227272 237969 227300 238138
rect 227258 237960 227314 237969
rect 227258 237895 227314 237904
rect 226984 237788 227036 237794
rect 226984 237730 227036 237736
rect 226892 236632 226944 236638
rect 226892 236574 226944 236580
rect 226800 235272 226852 235278
rect 226800 235214 226852 235220
rect 226720 233838 226932 233866
rect 226628 233702 226748 233730
rect 226616 233640 226668 233646
rect 226616 233582 226668 233588
rect 226524 227180 226576 227186
rect 226524 227122 226576 227128
rect 226340 224324 226392 224330
rect 226340 224266 226392 224272
rect 226628 222902 226656 233582
rect 226720 229094 226748 233702
rect 226720 229066 226840 229094
rect 226616 222896 226668 222902
rect 226616 222838 226668 222844
rect 226340 220448 226392 220454
rect 226340 220390 226392 220396
rect 226352 220114 226380 220390
rect 226340 220108 226392 220114
rect 226340 220050 226392 220056
rect 225788 192500 225840 192506
rect 225788 192442 225840 192448
rect 225328 180124 225380 180130
rect 225328 180066 225380 180072
rect 226812 177342 226840 229066
rect 226904 206310 226932 233838
rect 227364 233646 227392 239634
rect 227548 239578 227576 239702
rect 227870 239720 227944 239748
rect 227626 239663 227682 239672
rect 227456 239550 227576 239578
rect 227352 233640 227404 233646
rect 227352 233582 227404 233588
rect 227456 230738 227484 239550
rect 227536 238264 227588 238270
rect 227536 238206 227588 238212
rect 227180 230710 227484 230738
rect 227076 222896 227128 222902
rect 227076 222838 227128 222844
rect 226984 220788 227036 220794
rect 226984 220730 227036 220736
rect 226996 220386 227024 220730
rect 226984 220380 227036 220386
rect 226984 220322 227036 220328
rect 226996 211886 227024 220322
rect 226984 211880 227036 211886
rect 226984 211822 227036 211828
rect 226892 206304 226944 206310
rect 226892 206246 226944 206252
rect 226982 199472 227038 199481
rect 226982 199407 227038 199416
rect 226800 177336 226852 177342
rect 226800 177278 226852 177284
rect 226338 156632 226394 156641
rect 226338 156567 226394 156576
rect 225064 16546 225184 16574
rect 224316 11756 224368 11762
rect 224316 11698 224368 11704
rect 223948 3120 224000 3126
rect 223948 3062 224000 3068
rect 223960 480 223988 3062
rect 225156 480 225184 16546
rect 226352 3466 226380 156567
rect 226432 3596 226484 3602
rect 226432 3538 226484 3544
rect 226340 3460 226392 3466
rect 226340 3402 226392 3408
rect 226444 1850 226472 3538
rect 226996 3126 227024 199407
rect 227088 198014 227116 222838
rect 227180 220454 227208 230710
rect 227260 230648 227312 230654
rect 227260 230590 227312 230596
rect 227272 220794 227300 230590
rect 227548 229094 227576 238206
rect 227640 238134 227668 239663
rect 227720 239624 227772 239630
rect 227718 239592 227720 239601
rect 227772 239592 227774 239601
rect 227718 239527 227774 239536
rect 227916 239034 227944 239720
rect 228284 239720 228358 239748
rect 228422 239748 228450 240108
rect 228514 239873 228542 240108
rect 228606 239902 228634 240108
rect 228698 239970 228726 240108
rect 228686 239964 228738 239970
rect 228686 239906 228738 239912
rect 228594 239896 228646 239902
rect 228500 239864 228556 239873
rect 228790 239873 228818 240108
rect 228882 239970 228910 240108
rect 228974 239970 229002 240108
rect 228870 239964 228922 239970
rect 228870 239906 228922 239912
rect 228962 239964 229014 239970
rect 228962 239906 229014 239912
rect 229066 239902 229094 240108
rect 229054 239896 229106 239902
rect 228594 239838 228646 239844
rect 228776 239864 228832 239873
rect 228500 239799 228556 239808
rect 228776 239799 228832 239808
rect 229052 239864 229054 239873
rect 229106 239864 229108 239873
rect 229052 239799 229108 239808
rect 228548 239760 228600 239766
rect 228422 239720 228496 239748
rect 228180 239692 228232 239698
rect 228100 239652 228180 239680
rect 227916 239006 228036 239034
rect 227902 238912 227958 238921
rect 227902 238847 227958 238856
rect 227718 238776 227774 238785
rect 227718 238711 227774 238720
rect 227628 238128 227680 238134
rect 227628 238070 227680 238076
rect 227732 233322 227760 238711
rect 227916 235994 227944 238847
rect 228008 238105 228036 239006
rect 227994 238096 228050 238105
rect 227994 238031 228050 238040
rect 227824 235966 227944 235994
rect 227994 236056 228050 236065
rect 227994 235991 228050 236000
rect 227824 233442 227852 235966
rect 227904 233844 227956 233850
rect 227904 233786 227956 233792
rect 227916 233458 227944 233786
rect 228008 233646 228036 235991
rect 227996 233640 228048 233646
rect 227996 233582 228048 233588
rect 227812 233436 227864 233442
rect 227916 233430 228036 233458
rect 227812 233378 227864 233384
rect 227732 233294 227944 233322
rect 227812 233096 227864 233102
rect 227812 233038 227864 233044
rect 227720 232212 227772 232218
rect 227720 232154 227772 232160
rect 227364 229066 227576 229094
rect 227260 220788 227312 220794
rect 227260 220730 227312 220736
rect 227168 220448 227220 220454
rect 227168 220390 227220 220396
rect 227076 198008 227128 198014
rect 227076 197950 227128 197956
rect 227364 155242 227392 229066
rect 227352 155236 227404 155242
rect 227352 155178 227404 155184
rect 227732 6914 227760 232154
rect 227824 8974 227852 233038
rect 227812 8968 227864 8974
rect 227812 8910 227864 8916
rect 227732 6886 227852 6914
rect 227536 3460 227588 3466
rect 227536 3402 227588 3408
rect 226984 3120 227036 3126
rect 226984 3062 227036 3068
rect 226352 1822 226472 1850
rect 226352 480 226380 1822
rect 227548 480 227576 3402
rect 227824 490 227852 6886
rect 227916 4826 227944 233294
rect 228008 219201 228036 233430
rect 228100 220794 228128 239652
rect 228180 239634 228232 239640
rect 228180 239556 228232 239562
rect 228180 239498 228232 239504
rect 228192 239465 228220 239498
rect 228178 239456 228234 239465
rect 228178 239391 228234 239400
rect 228284 233986 228312 239720
rect 228364 239556 228416 239562
rect 228364 239498 228416 239504
rect 228376 239465 228404 239498
rect 228362 239456 228418 239465
rect 228362 239391 228418 239400
rect 228364 239080 228416 239086
rect 228364 239022 228416 239028
rect 228376 236298 228404 239022
rect 228364 236292 228416 236298
rect 228364 236234 228416 236240
rect 228468 235994 228496 239720
rect 228548 239702 228600 239708
rect 228824 239760 228876 239766
rect 229008 239760 229060 239766
rect 228824 239702 228876 239708
rect 228914 239728 228970 239737
rect 228376 235966 228496 235994
rect 228272 233980 228324 233986
rect 228272 233922 228324 233928
rect 228376 233866 228404 235966
rect 228192 233838 228404 233866
rect 228560 233850 228588 239702
rect 228640 239624 228692 239630
rect 228640 239566 228692 239572
rect 228732 239624 228784 239630
rect 228732 239566 228784 239572
rect 228548 233844 228600 233850
rect 228088 220788 228140 220794
rect 228088 220730 228140 220736
rect 228192 220590 228220 233838
rect 228548 233786 228600 233792
rect 228652 233730 228680 239566
rect 228744 237726 228772 239566
rect 228836 237969 228864 239702
rect 229158 239748 229186 240108
rect 229008 239702 229060 239708
rect 229112 239720 229186 239748
rect 229250 239748 229278 240108
rect 229342 239873 229370 240108
rect 229328 239864 229384 239873
rect 229328 239799 229384 239808
rect 229434 239748 229462 240108
rect 229250 239720 229324 239748
rect 228914 239663 228970 239672
rect 228928 238338 228956 239663
rect 229020 238921 229048 239702
rect 229006 238912 229062 238921
rect 229006 238847 229062 238856
rect 229006 238640 229062 238649
rect 229006 238575 229008 238584
rect 229060 238575 229062 238584
rect 229008 238546 229060 238552
rect 228916 238332 228968 238338
rect 228916 238274 228968 238280
rect 228914 238232 228970 238241
rect 228914 238167 228970 238176
rect 228822 237960 228878 237969
rect 228822 237895 228878 237904
rect 228732 237720 228784 237726
rect 228732 237662 228784 237668
rect 228732 236904 228784 236910
rect 228732 236846 228784 236852
rect 228744 236609 228772 236846
rect 228730 236600 228786 236609
rect 228730 236535 228786 236544
rect 228732 235272 228784 235278
rect 228732 235214 228784 235220
rect 228284 233702 228680 233730
rect 228284 220833 228312 233702
rect 228456 233640 228508 233646
rect 228456 233582 228508 233588
rect 228364 223236 228416 223242
rect 228364 223178 228416 223184
rect 228376 222970 228404 223178
rect 228364 222964 228416 222970
rect 228364 222906 228416 222912
rect 228270 220824 228326 220833
rect 228270 220759 228326 220768
rect 228180 220584 228232 220590
rect 228180 220526 228232 220532
rect 227994 219192 228050 219201
rect 227994 219127 228050 219136
rect 228008 217394 228036 219127
rect 227996 217388 228048 217394
rect 227996 217330 228048 217336
rect 228192 209774 228220 220526
rect 228192 209746 228404 209774
rect 228376 159390 228404 209746
rect 228468 178702 228496 233582
rect 228744 232218 228772 235214
rect 228824 233980 228876 233986
rect 228824 233922 228876 233928
rect 228732 232212 228784 232218
rect 228732 232154 228784 232160
rect 228836 223242 228864 233922
rect 228928 231130 228956 238167
rect 229112 237930 229140 239720
rect 229192 239624 229244 239630
rect 229192 239566 229244 239572
rect 229100 237924 229152 237930
rect 229100 237866 229152 237872
rect 229204 235958 229232 239566
rect 229192 235952 229244 235958
rect 229192 235894 229244 235900
rect 228916 231124 228968 231130
rect 228916 231066 228968 231072
rect 228824 223236 228876 223242
rect 228824 223178 228876 223184
rect 229296 222154 229324 239720
rect 229388 239720 229462 239748
rect 229526 239748 229554 240108
rect 229618 239902 229646 240108
rect 229606 239896 229658 239902
rect 229606 239838 229658 239844
rect 229710 239748 229738 240108
rect 229526 239720 229600 239748
rect 229388 236502 229416 239720
rect 229466 239456 229522 239465
rect 229466 239391 229522 239400
rect 229480 239193 229508 239391
rect 229466 239184 229522 239193
rect 229466 239119 229522 239128
rect 229466 238640 229522 238649
rect 229466 238575 229522 238584
rect 229480 238474 229508 238575
rect 229468 238468 229520 238474
rect 229468 238410 229520 238416
rect 229376 236496 229428 236502
rect 229376 236438 229428 236444
rect 229572 234122 229600 239720
rect 229664 239720 229738 239748
rect 229664 237425 229692 239720
rect 229802 239578 229830 240108
rect 229894 239850 229922 240108
rect 229986 239970 230014 240108
rect 229974 239964 230026 239970
rect 229974 239906 230026 239912
rect 230078 239902 230106 240108
rect 230066 239896 230118 239902
rect 229894 239822 229968 239850
rect 230066 239838 230118 239844
rect 230170 239850 230198 240108
rect 230262 239970 230290 240108
rect 230250 239964 230302 239970
rect 230250 239906 230302 239912
rect 230354 239902 230382 240108
rect 230342 239896 230394 239902
rect 230170 239822 230244 239850
rect 230342 239838 230394 239844
rect 230446 239850 230474 240108
rect 230538 239970 230566 240108
rect 230526 239964 230578 239970
rect 230526 239906 230578 239912
rect 230446 239822 230520 239850
rect 229802 239550 229876 239578
rect 229742 239184 229798 239193
rect 229742 239119 229744 239128
rect 229796 239119 229798 239128
rect 229744 239090 229796 239096
rect 229650 237416 229706 237425
rect 229650 237351 229706 237360
rect 229560 234116 229612 234122
rect 229560 234058 229612 234064
rect 229848 234002 229876 239550
rect 229940 238474 229968 239822
rect 230020 239760 230072 239766
rect 230020 239702 230072 239708
rect 230112 239760 230164 239766
rect 230216 239737 230244 239822
rect 230296 239760 230348 239766
rect 230112 239702 230164 239708
rect 230202 239728 230258 239737
rect 229928 238468 229980 238474
rect 229928 238410 229980 238416
rect 229388 233974 229876 234002
rect 229388 225758 229416 233974
rect 229940 233866 229968 238410
rect 230032 237182 230060 239702
rect 230124 238785 230152 239702
rect 230388 239760 230440 239766
rect 230296 239702 230348 239708
rect 230386 239728 230388 239737
rect 230440 239728 230442 239737
rect 230202 239663 230258 239672
rect 230110 238776 230166 238785
rect 230110 238711 230166 238720
rect 230110 238232 230166 238241
rect 230110 238167 230166 238176
rect 230020 237176 230072 237182
rect 230020 237118 230072 237124
rect 229744 233844 229796 233850
rect 229744 233786 229796 233792
rect 229848 233838 229968 233866
rect 229376 225752 229428 225758
rect 229376 225694 229428 225700
rect 229284 222148 229336 222154
rect 229284 222090 229336 222096
rect 228730 220824 228786 220833
rect 228548 220788 228600 220794
rect 228730 220759 228786 220768
rect 228548 220730 228600 220736
rect 228560 220318 228588 220730
rect 228548 220312 228600 220318
rect 228548 220254 228600 220260
rect 228560 195294 228588 220254
rect 228744 219881 228772 220759
rect 228730 219872 228786 219881
rect 228730 219807 228786 219816
rect 228744 204950 228772 219807
rect 228732 204944 228784 204950
rect 228732 204886 228784 204892
rect 228548 195288 228600 195294
rect 228548 195230 228600 195236
rect 228456 178696 228508 178702
rect 228456 178638 228508 178644
rect 228364 159384 228416 159390
rect 228364 159326 228416 159332
rect 229756 7614 229784 233786
rect 229848 170406 229876 233838
rect 230124 229094 230152 238167
rect 230216 238066 230244 239663
rect 230204 238060 230256 238066
rect 230204 238002 230256 238008
rect 230204 234116 230256 234122
rect 230204 234058 230256 234064
rect 229940 229066 230152 229094
rect 229940 173194 229968 229066
rect 230020 225752 230072 225758
rect 230020 225694 230072 225700
rect 230032 225418 230060 225694
rect 230020 225412 230072 225418
rect 230020 225354 230072 225360
rect 230032 191146 230060 225354
rect 230112 222148 230164 222154
rect 230112 222090 230164 222096
rect 230124 221678 230152 222090
rect 230112 221672 230164 221678
rect 230112 221614 230164 221620
rect 230124 210526 230152 221614
rect 230216 219026 230244 234058
rect 230308 219230 230336 239702
rect 230386 239663 230442 239672
rect 230388 239624 230440 239630
rect 230386 239592 230388 239601
rect 230440 239592 230442 239601
rect 230386 239527 230442 239536
rect 230386 239184 230442 239193
rect 230386 239119 230442 239128
rect 230400 238406 230428 239119
rect 230492 238406 230520 239822
rect 230630 239748 230658 240108
rect 230722 239850 230750 240108
rect 230814 239970 230842 240108
rect 230802 239964 230854 239970
rect 230802 239906 230854 239912
rect 230906 239902 230934 240108
rect 230894 239896 230946 239902
rect 230722 239822 230796 239850
rect 230894 239838 230946 239844
rect 230630 239720 230704 239748
rect 230768 239737 230796 239822
rect 230998 239748 231026 240108
rect 230572 239556 230624 239562
rect 230572 239498 230624 239504
rect 230388 238400 230440 238406
rect 230388 238342 230440 238348
rect 230480 238400 230532 238406
rect 230480 238342 230532 238348
rect 230492 238184 230520 238342
rect 230400 238156 230520 238184
rect 230400 233850 230428 238156
rect 230480 238060 230532 238066
rect 230480 238002 230532 238008
rect 230492 235754 230520 238002
rect 230480 235748 230532 235754
rect 230480 235690 230532 235696
rect 230388 233844 230440 233850
rect 230388 233786 230440 233792
rect 230492 221542 230520 235690
rect 230584 235482 230612 239498
rect 230676 237561 230704 239720
rect 230754 239728 230810 239737
rect 230952 239720 231026 239748
rect 231090 239748 231118 240108
rect 231182 239873 231210 240108
rect 231274 239970 231302 240108
rect 231366 239970 231394 240108
rect 231458 239970 231486 240108
rect 231262 239964 231314 239970
rect 231262 239906 231314 239912
rect 231354 239964 231406 239970
rect 231354 239906 231406 239912
rect 231446 239964 231498 239970
rect 231446 239906 231498 239912
rect 231168 239864 231224 239873
rect 231550 239850 231578 240108
rect 231642 239970 231670 240108
rect 231630 239964 231682 239970
rect 231630 239906 231682 239912
rect 231734 239850 231762 240108
rect 231826 239902 231854 240108
rect 231918 239902 231946 240108
rect 231168 239799 231224 239808
rect 231412 239822 231578 239850
rect 231688 239822 231762 239850
rect 231814 239896 231866 239902
rect 231814 239838 231866 239844
rect 231906 239896 231958 239902
rect 232010 239873 232038 240108
rect 232102 239902 232130 240108
rect 232090 239896 232142 239902
rect 231906 239838 231958 239844
rect 231996 239864 232052 239873
rect 231090 239720 231164 239748
rect 230810 239686 230888 239714
rect 230754 239663 230810 239672
rect 230756 239624 230808 239630
rect 230756 239566 230808 239572
rect 230662 237552 230718 237561
rect 230662 237487 230718 237496
rect 230572 235476 230624 235482
rect 230572 235418 230624 235424
rect 230768 228138 230796 239566
rect 230860 235346 230888 239686
rect 230952 238270 230980 239720
rect 231032 239624 231084 239630
rect 231032 239566 231084 239572
rect 230940 238264 230992 238270
rect 230940 238206 230992 238212
rect 230848 235340 230900 235346
rect 230848 235282 230900 235288
rect 230848 229152 230900 229158
rect 230848 229094 230900 229100
rect 230756 228132 230808 228138
rect 230756 228074 230808 228080
rect 230480 221536 230532 221542
rect 230480 221478 230532 221484
rect 230296 219224 230348 219230
rect 230296 219166 230348 219172
rect 230204 219020 230256 219026
rect 230204 218962 230256 218968
rect 230216 214674 230244 218962
rect 230308 218822 230336 219166
rect 230296 218816 230348 218822
rect 230296 218758 230348 218764
rect 230204 214668 230256 214674
rect 230204 214610 230256 214616
rect 230112 210520 230164 210526
rect 230112 210462 230164 210468
rect 230020 191140 230072 191146
rect 230020 191082 230072 191088
rect 229928 173188 229980 173194
rect 229928 173130 229980 173136
rect 229836 170400 229888 170406
rect 229836 170342 229888 170348
rect 229744 7608 229796 7614
rect 229744 7550 229796 7556
rect 230860 6914 230888 229094
rect 230952 10334 230980 238206
rect 231044 238066 231072 239566
rect 231032 238060 231084 238066
rect 231032 238002 231084 238008
rect 231032 237924 231084 237930
rect 231032 237866 231084 237872
rect 231044 227118 231072 237866
rect 231136 236910 231164 239720
rect 231214 239728 231270 239737
rect 231214 239663 231270 239672
rect 231124 236904 231176 236910
rect 231124 236846 231176 236852
rect 231124 236768 231176 236774
rect 231124 236710 231176 236716
rect 231032 227112 231084 227118
rect 231032 227054 231084 227060
rect 230940 10328 230992 10334
rect 230940 10270 230992 10276
rect 230860 6886 231072 6914
rect 227904 4820 227956 4826
rect 227904 4762 227956 4768
rect 229836 3460 229888 3466
rect 229836 3402 229888 3408
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 227824 462 228312 490
rect 229848 480 229876 3402
rect 231044 480 231072 6886
rect 231136 6186 231164 236710
rect 231228 234614 231256 239663
rect 231308 239624 231360 239630
rect 231306 239592 231308 239601
rect 231360 239592 231362 239601
rect 231306 239527 231362 239536
rect 231412 237590 231440 239822
rect 231492 239760 231544 239766
rect 231492 239702 231544 239708
rect 231584 239760 231636 239766
rect 231584 239702 231636 239708
rect 231504 238785 231532 239702
rect 231490 238776 231546 238785
rect 231490 238711 231546 238720
rect 231400 237584 231452 237590
rect 231400 237526 231452 237532
rect 231412 236774 231440 237526
rect 231400 236768 231452 236774
rect 231400 236710 231452 236716
rect 231228 234586 231348 234614
rect 231320 232694 231348 234586
rect 231308 232688 231360 232694
rect 231308 232630 231360 232636
rect 231308 228132 231360 228138
rect 231308 228074 231360 228080
rect 231320 186998 231348 228074
rect 231308 186992 231360 186998
rect 231308 186934 231360 186940
rect 231504 185638 231532 238711
rect 231596 219094 231624 239702
rect 231688 238105 231716 239822
rect 232090 239838 232142 239844
rect 231996 239799 232052 239808
rect 231768 239760 231820 239766
rect 232194 239748 232222 240108
rect 231768 239702 231820 239708
rect 231872 239720 232222 239748
rect 232286 239748 232314 240108
rect 232378 239816 232406 240108
rect 232470 239970 232498 240108
rect 232458 239964 232510 239970
rect 232458 239906 232510 239912
rect 232562 239816 232590 240108
rect 232654 239907 232682 240108
rect 232746 239970 232774 240108
rect 232838 239970 232866 240108
rect 232734 239964 232786 239970
rect 232640 239898 232696 239907
rect 232734 239906 232786 239912
rect 232826 239964 232878 239970
rect 232826 239906 232878 239912
rect 232930 239907 232958 240108
rect 233022 239970 233050 240108
rect 233010 239964 233062 239970
rect 232640 239833 232696 239842
rect 232916 239898 232972 239907
rect 233010 239906 233062 239912
rect 232378 239788 232452 239816
rect 232286 239720 232360 239748
rect 231780 238338 231808 239702
rect 231872 239154 231900 239720
rect 231952 239624 232004 239630
rect 231952 239566 232004 239572
rect 232136 239624 232188 239630
rect 232136 239566 232188 239572
rect 231860 239148 231912 239154
rect 231860 239090 231912 239096
rect 231860 238536 231912 238542
rect 231860 238478 231912 238484
rect 231768 238332 231820 238338
rect 231768 238274 231820 238280
rect 231674 238096 231730 238105
rect 231674 238031 231730 238040
rect 231780 237930 231808 238274
rect 231872 238134 231900 238478
rect 231860 238128 231912 238134
rect 231860 238070 231912 238076
rect 231964 237969 231992 239566
rect 232148 239290 232176 239566
rect 232228 239556 232280 239562
rect 232228 239498 232280 239504
rect 232044 239284 232096 239290
rect 232044 239226 232096 239232
rect 232136 239284 232188 239290
rect 232136 239226 232188 239232
rect 232056 239154 232084 239226
rect 232240 239170 232268 239498
rect 232044 239148 232096 239154
rect 232044 239090 232096 239096
rect 232148 239142 232268 239170
rect 232148 238950 232176 239142
rect 232136 238944 232188 238950
rect 232136 238886 232188 238892
rect 232044 238536 232096 238542
rect 232044 238478 232096 238484
rect 231950 237960 232006 237969
rect 231768 237924 231820 237930
rect 231950 237895 232006 237904
rect 231768 237866 231820 237872
rect 231860 236700 231912 236706
rect 231860 236642 231912 236648
rect 231768 234252 231820 234258
rect 231768 234194 231820 234200
rect 231780 229094 231808 234194
rect 231872 233866 231900 236642
rect 231872 233838 231992 233866
rect 231780 229066 231900 229094
rect 231584 219088 231636 219094
rect 231584 219030 231636 219036
rect 231596 216102 231624 219030
rect 231584 216096 231636 216102
rect 231584 216038 231636 216044
rect 231492 185632 231544 185638
rect 231492 185574 231544 185580
rect 231124 6180 231176 6186
rect 231124 6122 231176 6128
rect 228284 354 228312 462
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 231872 354 231900 229066
rect 231964 205018 231992 233838
rect 232056 222193 232084 238478
rect 232148 236706 232176 238886
rect 232332 236978 232360 239720
rect 232424 237318 232452 239788
rect 232516 239788 232590 239816
rect 232780 239828 232832 239834
rect 232916 239833 232972 239842
rect 232412 237312 232464 237318
rect 232412 237254 232464 237260
rect 232320 236972 232372 236978
rect 232320 236914 232372 236920
rect 232136 236700 232188 236706
rect 232136 236642 232188 236648
rect 232332 229094 232360 236914
rect 232516 235346 232544 239788
rect 233114 239816 233142 240108
rect 233206 239970 233234 240108
rect 233298 239970 233326 240108
rect 233194 239964 233246 239970
rect 233194 239906 233246 239912
rect 233286 239964 233338 239970
rect 233286 239906 233338 239912
rect 232780 239770 232832 239776
rect 233068 239788 233142 239816
rect 232596 239692 232648 239698
rect 232596 239634 232648 239640
rect 232608 239601 232636 239634
rect 232688 239624 232740 239630
rect 232594 239592 232650 239601
rect 232688 239566 232740 239572
rect 232594 239527 232650 239536
rect 232700 239476 232728 239566
rect 232608 239448 232728 239476
rect 232608 238202 232636 239448
rect 232792 239408 232820 239770
rect 232964 239760 233016 239766
rect 232964 239702 233016 239708
rect 232870 239592 232926 239601
rect 232870 239527 232926 239536
rect 232700 239380 232820 239408
rect 232596 238196 232648 238202
rect 232596 238138 232648 238144
rect 232504 235340 232556 235346
rect 232504 235282 232556 235288
rect 232700 230382 232728 239380
rect 232780 239284 232832 239290
rect 232780 239226 232832 239232
rect 232792 238202 232820 239226
rect 232884 238542 232912 239527
rect 232872 238536 232924 238542
rect 232872 238478 232924 238484
rect 232780 238196 232832 238202
rect 232780 238138 232832 238144
rect 232688 230376 232740 230382
rect 232688 230318 232740 230324
rect 232596 229764 232648 229770
rect 232596 229706 232648 229712
rect 232332 229066 232544 229094
rect 232042 222184 232098 222193
rect 232042 222119 232098 222128
rect 231952 205012 232004 205018
rect 231952 204954 232004 204960
rect 232516 158030 232544 229066
rect 232608 166326 232636 229706
rect 232700 192574 232728 230318
rect 232792 200802 232820 238138
rect 232872 235340 232924 235346
rect 232872 235282 232924 235288
rect 232884 230246 232912 235282
rect 232976 233986 233004 239702
rect 232964 233980 233016 233986
rect 232964 233922 233016 233928
rect 232872 230240 232924 230246
rect 232872 230182 232924 230188
rect 232884 229094 232912 230182
rect 232976 229770 233004 233922
rect 232964 229764 233016 229770
rect 232964 229706 233016 229712
rect 232884 229066 233004 229094
rect 232870 222184 232926 222193
rect 232870 222119 232926 222128
rect 232884 209166 232912 222119
rect 232976 220182 233004 229066
rect 233068 227458 233096 239788
rect 233390 239748 233418 240108
rect 233482 239970 233510 240108
rect 233470 239964 233522 239970
rect 233470 239906 233522 239912
rect 233574 239748 233602 240108
rect 233666 239873 233694 240108
rect 233758 239902 233786 240108
rect 233850 239970 233878 240108
rect 233838 239964 233890 239970
rect 233838 239906 233890 239912
rect 233942 239907 233970 240108
rect 234034 239970 234062 240108
rect 234022 239964 234074 239970
rect 233746 239896 233798 239902
rect 233652 239864 233708 239873
rect 233746 239838 233798 239844
rect 233928 239898 233984 239907
rect 234022 239906 234074 239912
rect 233928 239833 233984 239842
rect 234126 239816 234154 240108
rect 233652 239799 233708 239808
rect 234080 239788 234154 239816
rect 233700 239760 233752 239766
rect 233146 239728 233202 239737
rect 233390 239720 233464 239748
rect 233574 239720 233648 239748
rect 233146 239663 233148 239672
rect 233200 239663 233202 239672
rect 233148 239634 233200 239640
rect 233436 239290 233464 239720
rect 233516 239624 233568 239630
rect 233516 239566 233568 239572
rect 233424 239284 233476 239290
rect 233424 239226 233476 239232
rect 233148 238740 233200 238746
rect 233148 238682 233200 238688
rect 233160 238542 233188 238682
rect 233330 238640 233386 238649
rect 233330 238575 233386 238584
rect 233148 238536 233200 238542
rect 233148 238478 233200 238484
rect 233240 231328 233292 231334
rect 233240 231270 233292 231276
rect 233056 227452 233108 227458
rect 233056 227394 233108 227400
rect 233068 225622 233096 227394
rect 233056 225616 233108 225622
rect 233056 225558 233108 225564
rect 232964 220176 233016 220182
rect 232964 220118 233016 220124
rect 232872 209160 232924 209166
rect 232872 209102 232924 209108
rect 232780 200796 232832 200802
rect 232780 200738 232832 200744
rect 232688 192568 232740 192574
rect 232688 192510 232740 192516
rect 232596 166320 232648 166326
rect 232596 166262 232648 166268
rect 232504 158024 232556 158030
rect 232504 157966 232556 157972
rect 233252 16574 233280 231270
rect 233344 218890 233372 238575
rect 233436 223038 233464 239226
rect 233528 235385 233556 239566
rect 233514 235376 233570 235385
rect 233514 235311 233570 235320
rect 233620 233918 233648 239720
rect 233700 239702 233752 239708
rect 233712 239601 233740 239702
rect 233792 239624 233844 239630
rect 233698 239592 233754 239601
rect 233792 239566 233844 239572
rect 233698 239527 233754 239536
rect 233700 238876 233752 238882
rect 233700 238818 233752 238824
rect 233712 237454 233740 238818
rect 233700 237448 233752 237454
rect 233700 237390 233752 237396
rect 233608 233912 233660 233918
rect 233608 233854 233660 233860
rect 233804 233594 233832 239566
rect 233976 239556 234028 239562
rect 233976 239498 234028 239504
rect 233988 234326 234016 239498
rect 233976 234320 234028 234326
rect 233976 234262 234028 234268
rect 233528 233566 233832 233594
rect 233528 224330 233556 233566
rect 233608 233504 233660 233510
rect 233608 233446 233660 233452
rect 233620 224913 233648 233446
rect 233884 230988 233936 230994
rect 233884 230930 233936 230936
rect 233700 230784 233752 230790
rect 233700 230726 233752 230732
rect 233712 226710 233740 230726
rect 233896 228546 233924 230930
rect 233884 228540 233936 228546
rect 233884 228482 233936 228488
rect 233700 226704 233752 226710
rect 233700 226646 233752 226652
rect 233988 225690 234016 234262
rect 234080 233238 234108 239788
rect 234218 239748 234246 240108
rect 234310 239873 234338 240108
rect 234402 239970 234430 240108
rect 234390 239964 234442 239970
rect 234390 239906 234442 239912
rect 234296 239864 234352 239873
rect 234494 239850 234522 240108
rect 234296 239799 234352 239808
rect 234448 239822 234522 239850
rect 234172 239720 234246 239748
rect 234172 233510 234200 239720
rect 234344 239692 234396 239698
rect 234344 239634 234396 239640
rect 234252 238740 234304 238746
rect 234252 238682 234304 238688
rect 234264 238649 234292 238682
rect 234250 238640 234306 238649
rect 234250 238575 234306 238584
rect 234356 234614 234384 239634
rect 234448 237017 234476 239822
rect 234586 239748 234614 240108
rect 234678 239873 234706 240108
rect 234664 239864 234720 239873
rect 234664 239799 234720 239808
rect 234770 239816 234798 240108
rect 234862 239970 234890 240108
rect 234850 239964 234902 239970
rect 234850 239906 234902 239912
rect 234954 239850 234982 240108
rect 235046 239970 235074 240108
rect 235034 239964 235086 239970
rect 235034 239906 235086 239912
rect 235138 239850 235166 240108
rect 235230 239902 235258 240108
rect 235322 239970 235350 240108
rect 235310 239964 235362 239970
rect 235310 239906 235362 239912
rect 234954 239822 235028 239850
rect 234770 239788 234844 239816
rect 234586 239720 234752 239748
rect 234620 239624 234672 239630
rect 234618 239592 234620 239601
rect 234672 239592 234674 239601
rect 234618 239527 234674 239536
rect 234724 239034 234752 239720
rect 234540 239006 234752 239034
rect 234434 237008 234490 237017
rect 234434 236943 234490 236952
rect 234264 234598 234384 234614
rect 234252 234592 234384 234598
rect 234304 234586 234384 234592
rect 234252 234534 234304 234540
rect 234160 233504 234212 233510
rect 234160 233446 234212 233452
rect 234068 233232 234120 233238
rect 234068 233174 234120 233180
rect 234080 230994 234108 233174
rect 234068 230988 234120 230994
rect 234068 230930 234120 230936
rect 234264 229094 234292 234534
rect 234344 234524 234396 234530
rect 234344 234466 234396 234472
rect 234356 233918 234384 234466
rect 234344 233912 234396 233918
rect 234344 233854 234396 233860
rect 234540 230790 234568 239006
rect 234620 238876 234672 238882
rect 234620 238818 234672 238824
rect 234632 238649 234660 238818
rect 234618 238640 234674 238649
rect 234618 238575 234674 238584
rect 234712 237924 234764 237930
rect 234712 237866 234764 237872
rect 234620 237380 234672 237386
rect 234620 237322 234672 237328
rect 234528 230784 234580 230790
rect 234528 230726 234580 230732
rect 234080 229066 234292 229094
rect 233976 225684 234028 225690
rect 233976 225626 234028 225632
rect 233606 224904 233662 224913
rect 233606 224839 233662 224848
rect 233620 224482 233648 224839
rect 233620 224454 234016 224482
rect 233516 224324 233568 224330
rect 233516 224266 233568 224272
rect 233424 223032 233476 223038
rect 233424 222974 233476 222980
rect 233528 219434 233556 224266
rect 233528 219406 233924 219434
rect 233332 218884 233384 218890
rect 233332 218826 233384 218832
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 233896 14482 233924 219406
rect 233988 217462 234016 224454
rect 233976 217456 234028 217462
rect 233976 217398 234028 217404
rect 233976 207596 234028 207602
rect 233976 207538 234028 207544
rect 233884 14476 233936 14482
rect 233884 14418 233936 14424
rect 233988 3602 234016 207538
rect 234080 162178 234108 229066
rect 234160 227044 234212 227050
rect 234160 226986 234212 226992
rect 234172 226710 234200 226986
rect 234160 226704 234212 226710
rect 234160 226646 234212 226652
rect 234172 206378 234200 226646
rect 234160 206372 234212 206378
rect 234160 206314 234212 206320
rect 234068 162172 234120 162178
rect 234068 162114 234120 162120
rect 233976 3596 234028 3602
rect 233976 3538 234028 3544
rect 234632 480 234660 237322
rect 234724 16574 234752 237866
rect 234816 234569 234844 239788
rect 234896 239760 234948 239766
rect 234896 239702 234948 239708
rect 234908 234841 234936 239702
rect 235000 239222 235028 239822
rect 235092 239822 235166 239850
rect 235218 239896 235270 239902
rect 235218 239838 235270 239844
rect 234988 239216 235040 239222
rect 234988 239158 235040 239164
rect 234894 234832 234950 234841
rect 234894 234767 234950 234776
rect 235092 234614 235120 239822
rect 235414 239816 235442 240108
rect 235506 239970 235534 240108
rect 235494 239964 235546 239970
rect 235494 239906 235546 239912
rect 235598 239816 235626 240108
rect 235368 239788 235442 239816
rect 235552 239788 235626 239816
rect 235172 239760 235224 239766
rect 235172 239702 235224 239708
rect 235184 238814 235212 239702
rect 235264 239692 235316 239698
rect 235264 239634 235316 239640
rect 235172 238808 235224 238814
rect 235172 238750 235224 238756
rect 235184 236366 235212 238750
rect 235172 236360 235224 236366
rect 235172 236302 235224 236308
rect 234908 234586 235120 234614
rect 234802 234560 234858 234569
rect 234802 234495 234858 234504
rect 234804 234456 234856 234462
rect 234804 234398 234856 234404
rect 234816 224398 234844 234398
rect 234908 224534 234936 234586
rect 235276 233050 235304 239634
rect 235368 234462 235396 239788
rect 235448 239556 235500 239562
rect 235448 239498 235500 239504
rect 235460 236298 235488 239498
rect 235448 236292 235500 236298
rect 235448 236234 235500 236240
rect 235356 234456 235408 234462
rect 235356 234398 235408 234404
rect 235000 233022 235304 233050
rect 235000 229906 235028 233022
rect 235552 229974 235580 239788
rect 235690 239748 235718 240108
rect 235782 239902 235810 240108
rect 235874 239970 235902 240108
rect 235862 239964 235914 239970
rect 235862 239906 235914 239912
rect 235770 239896 235822 239902
rect 235966 239873 235994 240108
rect 236058 239970 236086 240108
rect 236046 239964 236098 239970
rect 236046 239906 236098 239912
rect 235770 239838 235822 239844
rect 235952 239864 236008 239873
rect 235952 239799 236008 239808
rect 235908 239760 235960 239766
rect 235690 239737 235764 239748
rect 235690 239728 235778 239737
rect 235690 239720 235722 239728
rect 235644 239672 235722 239680
rect 235908 239702 235960 239708
rect 235998 239728 236054 239737
rect 235644 239663 235778 239672
rect 235816 239692 235868 239698
rect 235644 239652 235764 239663
rect 235644 236745 235672 239652
rect 235736 239603 235764 239652
rect 235816 239634 235868 239640
rect 235828 238134 235856 239634
rect 235816 238128 235868 238134
rect 235816 238070 235868 238076
rect 235724 237516 235776 237522
rect 235724 237458 235776 237464
rect 235630 236736 235686 236745
rect 235630 236671 235686 236680
rect 235736 235482 235764 237458
rect 235724 235476 235776 235482
rect 235724 235418 235776 235424
rect 235828 235006 235856 238070
rect 235816 235000 235868 235006
rect 235816 234942 235868 234948
rect 235724 234116 235776 234122
rect 235724 234058 235776 234064
rect 235736 232830 235764 234058
rect 235724 232824 235776 232830
rect 235724 232766 235776 232772
rect 235540 229968 235592 229974
rect 235540 229910 235592 229916
rect 234988 229900 235040 229906
rect 234988 229842 235040 229848
rect 234896 224528 234948 224534
rect 234896 224470 234948 224476
rect 234804 224392 234856 224398
rect 234804 224334 234856 224340
rect 235000 219434 235028 229842
rect 235080 229220 235132 229226
rect 235080 229162 235132 229168
rect 235092 228614 235120 229162
rect 235552 229094 235580 229910
rect 235920 229634 235948 239702
rect 236150 239680 236178 240108
rect 236242 239970 236270 240108
rect 236334 239970 236362 240108
rect 236230 239964 236282 239970
rect 236230 239906 236282 239912
rect 236322 239964 236374 239970
rect 236322 239906 236374 239912
rect 236426 239714 236454 240108
rect 236518 239902 236546 240108
rect 236506 239896 236558 239902
rect 236610 239873 236638 240108
rect 236702 239970 236730 240108
rect 236794 239970 236822 240108
rect 236690 239964 236742 239970
rect 236690 239906 236742 239912
rect 236782 239964 236834 239970
rect 236782 239906 236834 239912
rect 236506 239838 236558 239844
rect 236596 239864 236652 239873
rect 236596 239799 236652 239808
rect 235998 239663 236054 239672
rect 236012 236842 236040 239663
rect 236104 239652 236178 239680
rect 236380 239686 236454 239714
rect 236552 239760 236604 239766
rect 236886 239748 236914 240108
rect 236978 239907 237006 240108
rect 236964 239898 237020 239907
rect 237070 239902 237098 240108
rect 236964 239833 237020 239842
rect 237058 239896 237110 239902
rect 237058 239838 237110 239844
rect 237162 239816 237190 240108
rect 237254 239970 237282 240108
rect 237242 239964 237294 239970
rect 237242 239906 237294 239912
rect 237346 239850 237374 240108
rect 237300 239822 237374 239850
rect 237438 239850 237466 240108
rect 237530 239970 237558 240108
rect 237518 239964 237570 239970
rect 237518 239906 237570 239912
rect 237438 239822 237512 239850
rect 237162 239788 237236 239816
rect 236604 239720 236684 239748
rect 236552 239702 236604 239708
rect 236104 238218 236132 239652
rect 236184 239556 236236 239562
rect 236184 239498 236236 239504
rect 236196 239193 236224 239498
rect 236182 239184 236238 239193
rect 236182 239119 236238 239128
rect 236104 238190 236316 238218
rect 236184 238060 236236 238066
rect 236184 238002 236236 238008
rect 236000 236836 236052 236842
rect 236000 236778 236052 236784
rect 236196 235550 236224 238002
rect 236000 235544 236052 235550
rect 236000 235486 236052 235492
rect 236184 235544 236236 235550
rect 236184 235486 236236 235492
rect 236012 232898 236040 235486
rect 236092 234660 236144 234666
rect 236092 234602 236144 234608
rect 236000 232892 236052 232898
rect 236000 232834 236052 232840
rect 236000 231192 236052 231198
rect 236000 231134 236052 231140
rect 235908 229628 235960 229634
rect 235908 229570 235960 229576
rect 235920 229226 235948 229570
rect 235908 229220 235960 229226
rect 235908 229162 235960 229168
rect 235460 229066 235580 229094
rect 235080 228608 235132 228614
rect 235080 228550 235132 228556
rect 235000 219406 235396 219434
rect 235262 218104 235318 218113
rect 235262 218039 235318 218048
rect 234724 16546 235212 16574
rect 235184 3482 235212 16546
rect 235276 3670 235304 218039
rect 235368 198082 235396 219406
rect 235460 214742 235488 229066
rect 235632 224528 235684 224534
rect 235632 224470 235684 224476
rect 235540 224392 235592 224398
rect 235540 224334 235592 224340
rect 235448 214736 235500 214742
rect 235448 214678 235500 214684
rect 235552 210594 235580 224334
rect 235644 211954 235672 224470
rect 235632 211948 235684 211954
rect 235632 211890 235684 211896
rect 235540 210588 235592 210594
rect 235540 210530 235592 210536
rect 235356 198076 235408 198082
rect 235356 198018 235408 198024
rect 236012 16574 236040 231134
rect 236104 222018 236132 234602
rect 236288 229498 236316 238190
rect 236380 229838 236408 239686
rect 236552 239624 236604 239630
rect 236458 239592 236514 239601
rect 236552 239566 236604 239572
rect 236458 239527 236514 239536
rect 236472 239494 236500 239527
rect 236460 239488 236512 239494
rect 236460 239430 236512 239436
rect 236460 238808 236512 238814
rect 236460 238750 236512 238756
rect 236472 234666 236500 238750
rect 236564 237289 236592 239566
rect 236656 238814 236684 239720
rect 236840 239720 236914 239748
rect 237012 239760 237064 239766
rect 236736 239556 236788 239562
rect 236736 239498 236788 239504
rect 236644 238808 236696 238814
rect 236644 238750 236696 238756
rect 236642 238096 236698 238105
rect 236642 238031 236698 238040
rect 236550 237280 236606 237289
rect 236550 237215 236606 237224
rect 236460 234660 236512 234666
rect 236460 234602 236512 234608
rect 236552 234456 236604 234462
rect 236552 234398 236604 234404
rect 236564 234054 236592 234398
rect 236552 234048 236604 234054
rect 236552 233990 236604 233996
rect 236552 231532 236604 231538
rect 236552 231474 236604 231480
rect 236564 230042 236592 231474
rect 236552 230036 236604 230042
rect 236552 229978 236604 229984
rect 236368 229832 236420 229838
rect 236368 229774 236420 229780
rect 236656 229770 236684 238031
rect 236748 234122 236776 239498
rect 236840 237522 236868 239720
rect 237064 239708 237144 239714
rect 237012 239702 237144 239708
rect 237024 239686 237144 239702
rect 236828 237516 236880 237522
rect 236828 237458 236880 237464
rect 237116 234614 237144 239686
rect 237208 238066 237236 239788
rect 237300 239737 237328 239822
rect 237286 239728 237342 239737
rect 237286 239663 237342 239672
rect 237288 239624 237340 239630
rect 237288 239566 237340 239572
rect 237196 238060 237248 238066
rect 237196 238002 237248 238008
rect 237116 234586 237236 234614
rect 236736 234116 236788 234122
rect 236736 234058 236788 234064
rect 236736 230444 236788 230450
rect 236736 230386 236788 230392
rect 236644 229764 236696 229770
rect 236644 229706 236696 229712
rect 236276 229492 236328 229498
rect 236276 229434 236328 229440
rect 236092 222012 236144 222018
rect 236092 221954 236144 221960
rect 236104 220522 236132 221954
rect 236092 220516 236144 220522
rect 236092 220458 236144 220464
rect 236288 219434 236316 229434
rect 236656 227254 236684 229706
rect 236644 227248 236696 227254
rect 236644 227190 236696 227196
rect 236288 219406 236684 219434
rect 236656 196654 236684 219406
rect 236748 207738 236776 230386
rect 237208 221746 237236 234586
rect 237300 230450 237328 239566
rect 237484 236994 237512 239822
rect 237622 239816 237650 240108
rect 237714 239850 237742 240108
rect 237806 239970 237834 240108
rect 237794 239964 237846 239970
rect 237794 239906 237846 239912
rect 237714 239834 237788 239850
rect 237714 239828 237800 239834
rect 237714 239822 237748 239828
rect 237576 239788 237650 239816
rect 237576 237998 237604 239788
rect 237898 239816 237926 240108
rect 237990 239970 238018 240108
rect 238082 239970 238110 240108
rect 237978 239964 238030 239970
rect 237978 239906 238030 239912
rect 238070 239964 238122 239970
rect 238070 239906 238122 239912
rect 238174 239873 238202 240108
rect 238266 239970 238294 240108
rect 238254 239964 238306 239970
rect 238254 239906 238306 239912
rect 237748 239770 237800 239776
rect 237852 239788 237926 239816
rect 238160 239864 238216 239873
rect 238358 239816 238386 240108
rect 238216 239808 238248 239816
rect 238160 239799 238248 239808
rect 238174 239788 238248 239799
rect 237656 239692 237708 239698
rect 237656 239634 237708 239640
rect 237748 239692 237800 239698
rect 237748 239634 237800 239640
rect 237668 239086 237696 239634
rect 237760 239154 237788 239634
rect 237852 239578 237880 239788
rect 238024 239624 238076 239630
rect 237852 239550 237972 239578
rect 238024 239566 238076 239572
rect 237944 239329 237972 239550
rect 237930 239320 237986 239329
rect 237930 239255 237986 239264
rect 237748 239148 237800 239154
rect 237748 239090 237800 239096
rect 237932 239148 237984 239154
rect 237932 239090 237984 239096
rect 237656 239080 237708 239086
rect 237656 239022 237708 239028
rect 237944 238898 237972 239090
rect 238036 239018 238064 239566
rect 238116 239352 238168 239358
rect 238116 239294 238168 239300
rect 238024 239012 238076 239018
rect 238024 238954 238076 238960
rect 237944 238870 238064 238898
rect 237932 238808 237984 238814
rect 237932 238750 237984 238756
rect 237564 237992 237616 237998
rect 237564 237934 237616 237940
rect 237564 237176 237616 237182
rect 237564 237118 237616 237124
rect 237392 236966 237512 236994
rect 237392 235414 237420 236966
rect 237472 236700 237524 236706
rect 237472 236642 237524 236648
rect 237380 235408 237432 235414
rect 237380 235350 237432 235356
rect 237288 230444 237340 230450
rect 237288 230386 237340 230392
rect 237300 230110 237328 230386
rect 237288 230104 237340 230110
rect 237288 230046 237340 230052
rect 237378 222184 237434 222193
rect 237378 222119 237434 222128
rect 237196 221740 237248 221746
rect 237196 221682 237248 221688
rect 237208 217530 237236 221682
rect 237196 217524 237248 217530
rect 237196 217466 237248 217472
rect 236736 207732 236788 207738
rect 236736 207674 236788 207680
rect 236644 196648 236696 196654
rect 236644 196590 236696 196596
rect 237392 16574 237420 222119
rect 237484 206446 237512 236642
rect 237576 235278 237604 237118
rect 237656 235816 237708 235822
rect 237656 235758 237708 235764
rect 237564 235272 237616 235278
rect 237564 235214 237616 235220
rect 237668 235074 237696 235758
rect 237656 235068 237708 235074
rect 237656 235010 237708 235016
rect 237564 233912 237616 233918
rect 237564 233854 237616 233860
rect 237576 221882 237604 233854
rect 237944 231305 237972 238750
rect 238036 237374 238064 238870
rect 238128 238134 238156 239294
rect 238116 238128 238168 238134
rect 238116 238070 238168 238076
rect 238036 237346 238156 237374
rect 238128 236706 238156 237346
rect 238220 237153 238248 239788
rect 238312 239788 238386 239816
rect 238206 237144 238262 237153
rect 238206 237079 238262 237088
rect 238116 236700 238168 236706
rect 238116 236642 238168 236648
rect 237930 231296 237986 231305
rect 237930 231231 237986 231240
rect 238312 230994 238340 239788
rect 238450 239748 238478 240108
rect 238542 239834 238570 240108
rect 238530 239828 238582 239834
rect 238530 239770 238582 239776
rect 238404 239737 238478 239748
rect 238390 239728 238478 239737
rect 238446 239720 238478 239728
rect 238634 239714 238662 240108
rect 238726 239873 238754 240108
rect 238818 239902 238846 240108
rect 238910 239902 238938 240108
rect 238806 239896 238858 239902
rect 238712 239864 238768 239873
rect 238806 239838 238858 239844
rect 238898 239896 238950 239902
rect 238898 239838 238950 239844
rect 238712 239799 238768 239808
rect 239002 239816 239030 240108
rect 239094 239970 239122 240108
rect 239082 239964 239134 239970
rect 239082 239906 239134 239912
rect 239186 239902 239214 240108
rect 239174 239896 239226 239902
rect 239278 239873 239306 240108
rect 239370 239902 239398 240108
rect 239462 239970 239490 240108
rect 239554 239970 239582 240108
rect 239450 239964 239502 239970
rect 239450 239906 239502 239912
rect 239542 239964 239594 239970
rect 239542 239906 239594 239912
rect 239358 239896 239410 239902
rect 239174 239838 239226 239844
rect 239264 239864 239320 239873
rect 239002 239788 239076 239816
rect 239358 239838 239410 239844
rect 239264 239799 239320 239808
rect 239496 239828 239548 239834
rect 238634 239686 238708 239714
rect 238390 239663 238446 239672
rect 238392 239556 238444 239562
rect 238392 239498 238444 239504
rect 238484 239556 238536 239562
rect 238484 239498 238536 239504
rect 238404 239154 238432 239498
rect 238392 239148 238444 239154
rect 238392 239090 238444 239096
rect 238496 238542 238524 239498
rect 238574 239456 238630 239465
rect 238574 239391 238630 239400
rect 238484 238536 238536 238542
rect 238484 238478 238536 238484
rect 238588 237374 238616 239391
rect 238680 238814 238708 239686
rect 238944 239692 238996 239698
rect 238944 239634 238996 239640
rect 238760 239624 238812 239630
rect 238760 239566 238812 239572
rect 238668 238808 238720 238814
rect 238668 238750 238720 238756
rect 238404 237346 238616 237374
rect 238404 233918 238432 237346
rect 238772 235686 238800 239566
rect 238852 239556 238904 239562
rect 238852 239498 238904 239504
rect 238864 239329 238892 239498
rect 238850 239320 238906 239329
rect 238850 239255 238906 239264
rect 238760 235680 238812 235686
rect 238760 235622 238812 235628
rect 238956 235618 238984 239634
rect 238944 235612 238996 235618
rect 238944 235554 238996 235560
rect 238392 233912 238444 233918
rect 238392 233854 238444 233860
rect 238760 232824 238812 232830
rect 238760 232766 238812 232772
rect 238484 232756 238536 232762
rect 238484 232698 238536 232704
rect 237656 230988 237708 230994
rect 237656 230930 237708 230936
rect 238300 230988 238352 230994
rect 238300 230930 238352 230936
rect 237668 223106 237696 230930
rect 238024 229356 238076 229362
rect 238024 229298 238076 229304
rect 237656 223100 237708 223106
rect 237656 223042 237708 223048
rect 237564 221876 237616 221882
rect 237564 221818 237616 221824
rect 237576 213314 237604 221818
rect 237564 213308 237616 213314
rect 237564 213250 237616 213256
rect 237472 206440 237524 206446
rect 237472 206382 237524 206388
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 235264 3664 235316 3670
rect 235264 3606 235316 3612
rect 235184 3454 235856 3482
rect 235828 480 235856 3454
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 238036 3534 238064 229298
rect 238496 222193 238524 232698
rect 238482 222184 238538 222193
rect 238482 222119 238538 222128
rect 238772 16574 238800 232766
rect 239048 229094 239076 239788
rect 239496 239770 239548 239776
rect 239128 239760 239180 239766
rect 239220 239760 239272 239766
rect 239128 239702 239180 239708
rect 239218 239728 239220 239737
rect 239272 239728 239274 239737
rect 239508 239714 239536 239770
rect 239646 239748 239674 240108
rect 239738 239970 239766 240108
rect 239830 239970 239858 240108
rect 239726 239964 239778 239970
rect 239726 239906 239778 239912
rect 239818 239964 239870 239970
rect 239818 239906 239870 239912
rect 239922 239850 239950 240108
rect 240014 239970 240042 240108
rect 240002 239964 240054 239970
rect 240002 239906 240054 239912
rect 240106 239902 240134 240108
rect 240198 239970 240226 240108
rect 240186 239964 240238 239970
rect 240186 239906 240238 239912
rect 240290 239902 240318 240108
rect 239772 239828 239824 239834
rect 239772 239770 239824 239776
rect 239876 239822 239950 239850
rect 240094 239896 240146 239902
rect 240094 239838 240146 239844
rect 240278 239896 240330 239902
rect 240278 239838 240330 239844
rect 239646 239720 239720 239748
rect 239140 229566 239168 239702
rect 239218 239663 239274 239672
rect 239324 239686 239536 239714
rect 239218 239320 239274 239329
rect 239218 239255 239274 239264
rect 239232 238746 239260 239255
rect 239220 238740 239272 238746
rect 239220 238682 239272 238688
rect 239220 238128 239272 238134
rect 239220 238070 239272 238076
rect 239232 236910 239260 238070
rect 239220 236904 239272 236910
rect 239220 236846 239272 236852
rect 239324 231538 239352 239686
rect 239496 239624 239548 239630
rect 239496 239566 239548 239572
rect 239404 239556 239456 239562
rect 239404 239498 239456 239504
rect 239416 234462 239444 239498
rect 239508 238610 239536 239566
rect 239588 238944 239640 238950
rect 239588 238886 239640 238892
rect 239600 238814 239628 238886
rect 239588 238808 239640 238814
rect 239588 238750 239640 238756
rect 239496 238604 239548 238610
rect 239496 238546 239548 238552
rect 239494 237960 239550 237969
rect 239494 237895 239550 237904
rect 239508 237386 239536 237895
rect 239496 237380 239548 237386
rect 239496 237322 239548 237328
rect 239692 235074 239720 239720
rect 239680 235068 239732 235074
rect 239680 235010 239732 235016
rect 239404 234456 239456 234462
rect 239404 234398 239456 234404
rect 239784 233866 239812 239770
rect 239416 233838 239812 233866
rect 239312 231532 239364 231538
rect 239312 231474 239364 231480
rect 239416 230926 239444 233838
rect 239876 232966 239904 239822
rect 239956 239760 240008 239766
rect 239956 239702 240008 239708
rect 240140 239760 240192 239766
rect 240382 239748 240410 240108
rect 240140 239702 240192 239708
rect 240336 239720 240410 239748
rect 239588 232960 239640 232966
rect 239588 232902 239640 232908
rect 239864 232960 239916 232966
rect 239864 232902 239916 232908
rect 239404 230920 239456 230926
rect 239404 230862 239456 230868
rect 239128 229560 239180 229566
rect 239128 229502 239180 229508
rect 239140 229362 239168 229502
rect 239128 229356 239180 229362
rect 239128 229298 239180 229304
rect 238864 229066 239076 229094
rect 238864 221785 238892 229066
rect 238850 221776 238906 221785
rect 238850 221711 238906 221720
rect 239416 181558 239444 230862
rect 239496 230512 239548 230518
rect 239496 230454 239548 230460
rect 239508 207602 239536 230454
rect 239600 216170 239628 232902
rect 239968 230994 239996 239702
rect 240048 239692 240100 239698
rect 240048 239634 240100 239640
rect 240060 239601 240088 239634
rect 240046 239592 240102 239601
rect 240046 239527 240102 239536
rect 240152 237182 240180 239702
rect 240232 239692 240284 239698
rect 240232 239634 240284 239640
rect 240244 238066 240272 239634
rect 240232 238060 240284 238066
rect 240232 238002 240284 238008
rect 240140 237176 240192 237182
rect 240140 237118 240192 237124
rect 240336 235994 240364 239720
rect 240474 239680 240502 240108
rect 240566 239748 240594 240108
rect 240658 239907 240686 240108
rect 240750 239970 240778 240108
rect 240738 239964 240790 239970
rect 240644 239898 240700 239907
rect 240738 239906 240790 239912
rect 240644 239833 240700 239842
rect 240842 239816 240870 240108
rect 240934 239970 240962 240108
rect 240922 239964 240974 239970
rect 240922 239906 240974 239912
rect 241026 239816 241054 240108
rect 240796 239788 240870 239816
rect 240980 239788 241054 239816
rect 240692 239760 240744 239766
rect 240566 239720 240640 239748
rect 240474 239652 240548 239680
rect 240416 238060 240468 238066
rect 240416 238002 240468 238008
rect 240244 235966 240364 235994
rect 239956 230988 240008 230994
rect 239956 230930 240008 230936
rect 239968 230518 239996 230930
rect 239956 230512 240008 230518
rect 239956 230454 240008 230460
rect 240048 229152 240100 229158
rect 240048 229094 240100 229100
rect 240244 229094 240272 235966
rect 240324 231940 240376 231946
rect 240324 231882 240376 231888
rect 240060 229066 240272 229094
rect 240060 225758 240088 229066
rect 240336 227254 240364 231882
rect 240428 231470 240456 238002
rect 240520 234258 240548 239652
rect 240508 234252 240560 234258
rect 240508 234194 240560 234200
rect 240416 231464 240468 231470
rect 240416 231406 240468 231412
rect 240612 231334 240640 239720
rect 240692 239702 240744 239708
rect 240704 232762 240732 239702
rect 240692 232756 240744 232762
rect 240692 232698 240744 232704
rect 240796 231554 240824 239788
rect 240876 238740 240928 238746
rect 240876 238682 240928 238688
rect 240888 231946 240916 238682
rect 240980 232830 241008 239788
rect 241118 239748 241146 240108
rect 241210 239970 241238 240108
rect 241198 239964 241250 239970
rect 241198 239906 241250 239912
rect 241302 239902 241330 240108
rect 241290 239896 241342 239902
rect 241290 239838 241342 239844
rect 241072 239720 241146 239748
rect 241244 239760 241296 239766
rect 240968 232824 241020 232830
rect 240968 232766 241020 232772
rect 240876 231940 240928 231946
rect 240876 231882 240928 231888
rect 240796 231526 240916 231554
rect 240784 231464 240836 231470
rect 240784 231406 240836 231412
rect 240600 231328 240652 231334
rect 240600 231270 240652 231276
rect 240324 227248 240376 227254
rect 240324 227190 240376 227196
rect 240140 226364 240192 226370
rect 240140 226306 240192 226312
rect 240048 225752 240100 225758
rect 240048 225694 240100 225700
rect 239588 216164 239640 216170
rect 239588 216106 239640 216112
rect 239496 207596 239548 207602
rect 239496 207538 239548 207544
rect 239404 181552 239456 181558
rect 239404 181494 239456 181500
rect 238772 16546 239352 16574
rect 238024 3528 238076 3534
rect 238024 3470 238076 3476
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 226306
rect 240796 3466 240824 231406
rect 240888 231198 240916 231526
rect 240876 231192 240928 231198
rect 240876 231134 240928 231140
rect 241072 226914 241100 239720
rect 241394 239748 241422 240108
rect 241486 239970 241514 240108
rect 241474 239964 241526 239970
rect 241474 239906 241526 239912
rect 241578 239748 241606 240108
rect 241394 239720 241468 239748
rect 241244 239702 241296 239708
rect 241152 239624 241204 239630
rect 241152 239566 241204 239572
rect 241060 226908 241112 226914
rect 241060 226850 241112 226856
rect 241072 226370 241100 226850
rect 241060 226364 241112 226370
rect 241060 226306 241112 226312
rect 241164 222154 241192 239566
rect 241256 232762 241284 239702
rect 241334 239592 241390 239601
rect 241334 239527 241336 239536
rect 241388 239527 241390 239536
rect 241336 239498 241388 239504
rect 241348 236706 241376 239498
rect 241440 238746 241468 239720
rect 241532 239720 241606 239748
rect 241428 238740 241480 238746
rect 241428 238682 241480 238688
rect 241532 238542 241560 239720
rect 241670 239680 241698 240108
rect 241762 239873 241790 240108
rect 241854 239902 241882 240108
rect 241946 239970 241974 240108
rect 242038 239970 242066 240108
rect 241934 239964 241986 239970
rect 241934 239906 241986 239912
rect 242026 239964 242078 239970
rect 242026 239906 242078 239912
rect 241842 239896 241894 239902
rect 241748 239864 241804 239873
rect 241842 239838 241894 239844
rect 242038 239816 242066 239906
rect 241748 239799 241804 239808
rect 241762 239748 241790 239799
rect 241992 239788 242066 239816
rect 241762 239720 241836 239748
rect 241670 239652 241744 239680
rect 241612 239556 241664 239562
rect 241612 239498 241664 239504
rect 241520 238536 241572 238542
rect 241520 238478 241572 238484
rect 241336 236700 241388 236706
rect 241336 236642 241388 236648
rect 241624 235994 241652 239498
rect 241532 235966 241652 235994
rect 241532 234054 241560 235966
rect 241610 235920 241666 235929
rect 241610 235855 241666 235864
rect 241520 234048 241572 234054
rect 241520 233990 241572 233996
rect 241520 233912 241572 233918
rect 241520 233854 241572 233860
rect 241244 232756 241296 232762
rect 241244 232698 241296 232704
rect 241428 232756 241480 232762
rect 241428 232698 241480 232704
rect 241336 227520 241388 227526
rect 241336 227462 241388 227468
rect 241348 227254 241376 227462
rect 241336 227248 241388 227254
rect 241336 227190 241388 227196
rect 241152 222148 241204 222154
rect 241152 222090 241204 222096
rect 241348 3534 241376 227190
rect 241336 3528 241388 3534
rect 241336 3470 241388 3476
rect 241440 3466 241468 232698
rect 241532 224262 241560 233854
rect 241520 224256 241572 224262
rect 241520 224198 241572 224204
rect 241520 222148 241572 222154
rect 241520 222090 241572 222096
rect 241532 221542 241560 222090
rect 241520 221536 241572 221542
rect 241520 221478 241572 221484
rect 241532 16574 241560 221478
rect 241624 162178 241652 235855
rect 241716 226846 241744 239652
rect 241808 231810 241836 239720
rect 241888 239692 241940 239698
rect 241888 239634 241940 239640
rect 241900 233918 241928 239634
rect 241992 239193 242020 239788
rect 242130 239748 242158 240108
rect 242222 239816 242250 240108
rect 242314 239970 242342 240108
rect 242406 239970 242434 240108
rect 242302 239964 242354 239970
rect 242302 239906 242354 239912
rect 242394 239964 242446 239970
rect 242394 239906 242446 239912
rect 242498 239873 242526 240108
rect 242590 239970 242618 240108
rect 242578 239964 242630 239970
rect 242578 239906 242630 239912
rect 242346 239864 242402 239873
rect 242222 239788 242296 239816
rect 242346 239799 242402 239808
rect 242484 239864 242540 239873
rect 242682 239816 242710 240108
rect 242774 239873 242802 240108
rect 242484 239799 242540 239808
rect 242084 239720 242158 239748
rect 241978 239184 242034 239193
rect 241978 239119 242034 239128
rect 241980 238740 242032 238746
rect 241980 238682 242032 238688
rect 241888 233912 241940 233918
rect 241888 233854 241940 233860
rect 241992 233170 242020 238682
rect 242084 235994 242112 239720
rect 242164 239624 242216 239630
rect 242164 239566 242216 239572
rect 242176 237930 242204 239566
rect 242268 238746 242296 239788
rect 242256 238740 242308 238746
rect 242256 238682 242308 238688
rect 242164 237924 242216 237930
rect 242164 237866 242216 237872
rect 242360 236745 242388 239799
rect 242636 239788 242710 239816
rect 242760 239864 242816 239873
rect 242760 239799 242816 239808
rect 242440 239760 242492 239766
rect 242440 239702 242492 239708
rect 242530 239728 242586 239737
rect 242452 238649 242480 239702
rect 242530 239663 242532 239672
rect 242584 239663 242586 239672
rect 242532 239634 242584 239640
rect 242544 239494 242572 239634
rect 242532 239488 242584 239494
rect 242532 239430 242584 239436
rect 242438 238640 242494 238649
rect 242438 238575 242494 238584
rect 242346 236736 242402 236745
rect 242346 236671 242402 236680
rect 242084 235966 242204 235994
rect 241980 233164 242032 233170
rect 241980 233106 242032 233112
rect 242176 233034 242204 235966
rect 242636 234614 242664 239788
rect 242866 239714 242894 240108
rect 242958 239902 242986 240108
rect 242946 239896 242998 239902
rect 243050 239873 243078 240108
rect 242946 239838 242998 239844
rect 243036 239864 243092 239873
rect 243036 239799 243092 239808
rect 242992 239760 243044 239766
rect 242866 239686 242940 239714
rect 243142 239748 243170 240108
rect 243234 239902 243262 240108
rect 243222 239896 243274 239902
rect 243222 239838 243274 239844
rect 243326 239850 243354 240108
rect 243418 239970 243446 240108
rect 243510 239970 243538 240108
rect 243406 239964 243458 239970
rect 243406 239906 243458 239912
rect 243498 239964 243550 239970
rect 243498 239906 243550 239912
rect 243326 239822 243400 239850
rect 243142 239720 243216 239748
rect 242992 239702 243044 239708
rect 242808 239624 242860 239630
rect 242912 239601 242940 239686
rect 242808 239566 242860 239572
rect 242898 239592 242954 239601
rect 242716 239488 242768 239494
rect 242716 239430 242768 239436
rect 242544 234586 242664 234614
rect 242728 234614 242756 239430
rect 242820 238066 242848 239566
rect 243004 239578 243032 239702
rect 243188 239601 243216 239720
rect 243372 239714 243400 239822
rect 243452 239828 243504 239834
rect 243602 239816 243630 240108
rect 243452 239770 243504 239776
rect 243556 239788 243630 239816
rect 243280 239686 243400 239714
rect 243174 239592 243230 239601
rect 243004 239550 243124 239578
rect 242898 239527 242954 239536
rect 242992 239488 243044 239494
rect 242992 239430 243044 239436
rect 243004 238678 243032 239430
rect 242992 238672 243044 238678
rect 242992 238614 243044 238620
rect 242808 238060 242860 238066
rect 242808 238002 242860 238008
rect 242820 237862 242848 238002
rect 242808 237856 242860 237862
rect 242808 237798 242860 237804
rect 242728 234586 242848 234614
rect 242256 234048 242308 234054
rect 242256 233990 242308 233996
rect 242164 233028 242216 233034
rect 242164 232970 242216 232976
rect 242268 232354 242296 233990
rect 242544 232558 242572 234586
rect 242716 233164 242768 233170
rect 242716 233106 242768 233112
rect 242532 232552 242584 232558
rect 242532 232494 242584 232500
rect 242728 232422 242756 233106
rect 242716 232416 242768 232422
rect 242716 232358 242768 232364
rect 242256 232348 242308 232354
rect 242256 232290 242308 232296
rect 241796 231804 241848 231810
rect 241796 231746 241848 231752
rect 241704 226840 241756 226846
rect 241704 226782 241756 226788
rect 242728 214606 242756 232358
rect 242716 214600 242768 214606
rect 242716 214542 242768 214548
rect 241612 162172 241664 162178
rect 241612 162114 241664 162120
rect 242820 33794 242848 234586
rect 243004 229094 243032 238614
rect 243096 237658 243124 239550
rect 243174 239527 243230 239536
rect 243084 237652 243136 237658
rect 243084 237594 243136 237600
rect 243084 236836 243136 236842
rect 243084 236778 243136 236784
rect 243096 229702 243124 236778
rect 243188 234054 243216 239527
rect 243280 235346 243308 239686
rect 243360 239624 243412 239630
rect 243360 239566 243412 239572
rect 243372 239465 243400 239566
rect 243358 239456 243414 239465
rect 243358 239391 243414 239400
rect 243464 236774 243492 239770
rect 243452 236768 243504 236774
rect 243452 236710 243504 236716
rect 243268 235340 243320 235346
rect 243268 235282 243320 235288
rect 243176 234048 243228 234054
rect 243176 233990 243228 233996
rect 243556 233714 243584 239788
rect 243694 239748 243722 240108
rect 243648 239720 243722 239748
rect 243786 239748 243814 240108
rect 243878 239816 243906 240108
rect 243970 239970 243998 240108
rect 243958 239964 244010 239970
rect 243958 239906 244010 239912
rect 244062 239816 244090 240108
rect 244154 239902 244182 240108
rect 244142 239896 244194 239902
rect 244142 239838 244194 239844
rect 243878 239788 243952 239816
rect 243786 239720 243860 239748
rect 243544 233708 243596 233714
rect 243544 233650 243596 233656
rect 243648 231962 243676 239720
rect 243832 238134 243860 239720
rect 243820 238128 243872 238134
rect 243820 238070 243872 238076
rect 243924 232626 243952 239788
rect 244016 239788 244090 239816
rect 244246 239816 244274 240108
rect 244338 239970 244366 240108
rect 244326 239964 244378 239970
rect 244326 239906 244378 239912
rect 244430 239850 244458 240108
rect 244522 239970 244550 240108
rect 244614 239970 244642 240108
rect 244510 239964 244562 239970
rect 244510 239906 244562 239912
rect 244602 239964 244654 239970
rect 244602 239906 244654 239912
rect 244706 239902 244734 240108
rect 244694 239896 244746 239902
rect 244430 239822 244504 239850
rect 244694 239838 244746 239844
rect 244246 239788 244320 239816
rect 244016 235278 244044 239788
rect 244096 239692 244148 239698
rect 244096 239634 244148 239640
rect 244188 239692 244240 239698
rect 244188 239634 244240 239640
rect 244004 235272 244056 235278
rect 244004 235214 244056 235220
rect 243912 232620 243964 232626
rect 243912 232562 243964 232568
rect 243556 231934 243676 231962
rect 243084 229696 243136 229702
rect 243084 229638 243136 229644
rect 242912 229066 243032 229094
rect 242808 33788 242860 33794
rect 242808 33730 242860 33736
rect 242912 16574 242940 229066
rect 243556 225486 243584 231934
rect 243636 231804 243688 231810
rect 243636 231746 243688 231752
rect 243544 225480 243596 225486
rect 243544 225422 243596 225428
rect 241532 16546 241744 16574
rect 242912 16546 243032 16574
rect 240784 3460 240836 3466
rect 240784 3402 240836 3408
rect 241428 3460 241480 3466
rect 241428 3402 241480 3408
rect 241716 480 241744 16546
rect 243004 3602 243032 16546
rect 242992 3596 243044 3602
rect 242992 3538 243044 3544
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 243648 3262 243676 231746
rect 244108 223038 244136 239634
rect 244200 236842 244228 239634
rect 244292 238649 244320 239788
rect 244372 239760 244424 239766
rect 244372 239702 244424 239708
rect 244278 238640 244334 238649
rect 244278 238575 244334 238584
rect 244188 236836 244240 236842
rect 244188 236778 244240 236784
rect 244280 236700 244332 236706
rect 244280 236642 244332 236648
rect 244188 234048 244240 234054
rect 244188 233990 244240 233996
rect 244096 223032 244148 223038
rect 244096 222974 244148 222980
rect 244200 215966 244228 233990
rect 244188 215960 244240 215966
rect 244188 215902 244240 215908
rect 244292 16574 244320 236642
rect 244384 235414 244412 239702
rect 244372 235408 244424 235414
rect 244372 235350 244424 235356
rect 244476 230738 244504 239822
rect 244798 239748 244826 240108
rect 244890 239902 244918 240108
rect 244878 239896 244930 239902
rect 244878 239838 244930 239844
rect 244982 239850 245010 240108
rect 245074 239970 245102 240108
rect 245062 239964 245114 239970
rect 245062 239906 245114 239912
rect 244982 239822 245056 239850
rect 244924 239760 244976 239766
rect 244798 239720 244872 239748
rect 244740 239624 244792 239630
rect 244740 239566 244792 239572
rect 244648 239420 244700 239426
rect 244648 239362 244700 239368
rect 244556 238740 244608 238746
rect 244556 238682 244608 238688
rect 244568 231010 244596 238682
rect 244660 237374 244688 239362
rect 244752 238746 244780 239566
rect 244740 238740 244792 238746
rect 244740 238682 244792 238688
rect 244844 238649 244872 239720
rect 244924 239702 244976 239708
rect 244830 238640 244886 238649
rect 244830 238575 244886 238584
rect 244832 238128 244884 238134
rect 244832 238070 244884 238076
rect 244660 237346 244780 237374
rect 244752 235994 244780 237346
rect 244844 236230 244872 238070
rect 244936 236842 244964 239702
rect 245028 238746 245056 239822
rect 245166 239816 245194 240108
rect 245120 239788 245194 239816
rect 245258 239816 245286 240108
rect 245350 239970 245378 240108
rect 245442 239970 245470 240108
rect 245534 239970 245562 240108
rect 245338 239964 245390 239970
rect 245338 239906 245390 239912
rect 245430 239964 245482 239970
rect 245430 239906 245482 239912
rect 245522 239964 245574 239970
rect 245522 239906 245574 239912
rect 245384 239828 245436 239834
rect 245258 239788 245332 239816
rect 245016 238740 245068 238746
rect 245016 238682 245068 238688
rect 244924 236836 244976 236842
rect 244924 236778 244976 236784
rect 244832 236224 244884 236230
rect 244832 236166 244884 236172
rect 244752 235966 244872 235994
rect 244844 231266 244872 235966
rect 245120 233850 245148 239788
rect 245198 239728 245254 239737
rect 245198 239663 245200 239672
rect 245252 239663 245254 239672
rect 245200 239634 245252 239640
rect 245198 239592 245254 239601
rect 245198 239527 245200 239536
rect 245252 239527 245254 239536
rect 245200 239498 245252 239504
rect 245200 238740 245252 238746
rect 245200 238682 245252 238688
rect 245108 233844 245160 233850
rect 245108 233786 245160 233792
rect 244832 231260 244884 231266
rect 244832 231202 244884 231208
rect 244568 230982 244780 231010
rect 244476 230710 244596 230738
rect 244464 230036 244516 230042
rect 244464 229978 244516 229984
rect 244372 229424 244424 229430
rect 244372 229366 244424 229372
rect 244384 209166 244412 229366
rect 244476 218890 244504 229978
rect 244568 227050 244596 230710
rect 244556 227044 244608 227050
rect 244556 226986 244608 226992
rect 244752 224954 244780 230982
rect 245212 230042 245240 238682
rect 245200 230036 245252 230042
rect 245200 229978 245252 229984
rect 245304 229430 245332 239788
rect 245626 239816 245654 240108
rect 245718 239970 245746 240108
rect 245706 239964 245758 239970
rect 245706 239906 245758 239912
rect 245810 239850 245838 240108
rect 245384 239770 245436 239776
rect 245488 239788 245654 239816
rect 245764 239822 245838 239850
rect 245396 233918 245424 239770
rect 245488 238649 245516 239788
rect 245568 239692 245620 239698
rect 245568 239634 245620 239640
rect 245660 239692 245712 239698
rect 245660 239634 245712 239640
rect 245474 238640 245530 238649
rect 245474 238575 245530 238584
rect 245580 237930 245608 239634
rect 245568 237924 245620 237930
rect 245568 237866 245620 237872
rect 245384 233912 245436 233918
rect 245384 233854 245436 233860
rect 245672 232898 245700 239634
rect 245764 238610 245792 239822
rect 245902 239748 245930 240108
rect 245994 239902 246022 240108
rect 245982 239896 246034 239902
rect 245982 239838 246034 239844
rect 246086 239816 246114 240108
rect 246178 239970 246206 240108
rect 246270 239970 246298 240108
rect 246362 239970 246390 240108
rect 246166 239964 246218 239970
rect 246166 239906 246218 239912
rect 246258 239964 246310 239970
rect 246258 239906 246310 239912
rect 246350 239964 246402 239970
rect 246350 239906 246402 239912
rect 246210 239864 246266 239873
rect 246086 239788 246160 239816
rect 246210 239799 246212 239808
rect 245856 239720 245930 239748
rect 245752 238604 245804 238610
rect 245752 238546 245804 238552
rect 245752 238128 245804 238134
rect 245752 238070 245804 238076
rect 245660 232892 245712 232898
rect 245660 232834 245712 232840
rect 245660 231872 245712 231878
rect 245660 231814 245712 231820
rect 245292 229424 245344 229430
rect 245292 229366 245344 229372
rect 244568 224926 244780 224954
rect 244568 220182 244596 224926
rect 245566 223136 245622 223145
rect 245566 223071 245622 223080
rect 244922 220824 244978 220833
rect 244922 220759 244978 220768
rect 244556 220176 244608 220182
rect 244556 220118 244608 220124
rect 244464 218884 244516 218890
rect 244464 218826 244516 218832
rect 244372 209160 244424 209166
rect 244372 209102 244424 209108
rect 244292 16546 244872 16574
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 244844 3482 244872 16546
rect 244936 4010 244964 220759
rect 244924 4004 244976 4010
rect 244924 3946 244976 3952
rect 243636 3256 243688 3262
rect 243636 3198 243688 3204
rect 244108 480 244136 3470
rect 244844 3454 245240 3482
rect 245580 3466 245608 223071
rect 245672 16574 245700 231814
rect 245764 208350 245792 238070
rect 245856 217870 245884 239720
rect 246028 239692 246080 239698
rect 246028 239634 246080 239640
rect 246040 239601 246068 239634
rect 246026 239592 246082 239601
rect 246026 239527 246082 239536
rect 245936 239488 245988 239494
rect 245936 239430 245988 239436
rect 245948 236706 245976 239430
rect 246028 238740 246080 238746
rect 246028 238682 246080 238688
rect 245936 236700 245988 236706
rect 245936 236642 245988 236648
rect 246040 228750 246068 238682
rect 246132 237794 246160 239788
rect 246264 239799 246266 239808
rect 246212 239770 246264 239776
rect 246454 239714 246482 240108
rect 246546 239970 246574 240108
rect 246534 239964 246586 239970
rect 246534 239906 246586 239912
rect 246638 239748 246666 240108
rect 246730 239850 246758 240108
rect 246822 239970 246850 240108
rect 246914 239970 246942 240108
rect 246810 239964 246862 239970
rect 246810 239906 246862 239912
rect 246902 239964 246954 239970
rect 246902 239906 246954 239912
rect 246730 239822 246804 239850
rect 246408 239686 246482 239714
rect 246592 239720 246666 239748
rect 246776 239737 246804 239822
rect 247006 239816 247034 240108
rect 246960 239788 247034 239816
rect 247098 239816 247126 240108
rect 247190 239970 247218 240108
rect 247178 239964 247230 239970
rect 247178 239906 247230 239912
rect 247282 239816 247310 240108
rect 247374 239970 247402 240108
rect 247362 239964 247414 239970
rect 247362 239906 247414 239912
rect 247466 239850 247494 240108
rect 247558 239970 247586 240108
rect 247546 239964 247598 239970
rect 247546 239906 247598 239912
rect 247098 239788 247172 239816
rect 246762 239728 246818 239737
rect 246212 239624 246264 239630
rect 246212 239566 246264 239572
rect 246120 237788 246172 237794
rect 246120 237730 246172 237736
rect 246224 235994 246252 239566
rect 246408 238626 246436 239686
rect 246488 239624 246540 239630
rect 246488 239566 246540 239572
rect 246500 238746 246528 239566
rect 246592 238746 246620 239720
rect 246762 239663 246818 239672
rect 246672 239624 246724 239630
rect 246672 239566 246724 239572
rect 246488 238740 246540 238746
rect 246488 238682 246540 238688
rect 246580 238740 246632 238746
rect 246580 238682 246632 238688
rect 246316 238598 246436 238626
rect 246316 238134 246344 238598
rect 246396 238536 246448 238542
rect 246396 238478 246448 238484
rect 246304 238128 246356 238134
rect 246304 238070 246356 238076
rect 246132 235966 246252 235994
rect 246132 230042 246160 235966
rect 246408 232694 246436 238478
rect 246684 235994 246712 239566
rect 246856 239556 246908 239562
rect 246856 239498 246908 239504
rect 246764 238740 246816 238746
rect 246764 238682 246816 238688
rect 246776 236570 246804 238682
rect 246764 236564 246816 236570
rect 246764 236506 246816 236512
rect 246592 235966 246712 235994
rect 246592 235686 246620 235966
rect 246580 235680 246632 235686
rect 246580 235622 246632 235628
rect 246762 234560 246818 234569
rect 246762 234495 246818 234504
rect 246396 232688 246448 232694
rect 246396 232630 246448 232636
rect 246408 231878 246436 232630
rect 246396 231872 246448 231878
rect 246396 231814 246448 231820
rect 246120 230036 246172 230042
rect 246120 229978 246172 229984
rect 246028 228744 246080 228750
rect 246028 228686 246080 228692
rect 246776 227254 246804 234495
rect 246868 228818 246896 239498
rect 246960 238649 246988 239788
rect 247040 239692 247092 239698
rect 247040 239634 247092 239640
rect 246946 238640 247002 238649
rect 246946 238575 247002 238584
rect 246948 238060 247000 238066
rect 246948 238002 247000 238008
rect 246960 237318 246988 238002
rect 246948 237312 247000 237318
rect 246948 237254 247000 237260
rect 246948 236768 247000 236774
rect 246948 236710 247000 236716
rect 246856 228812 246908 228818
rect 246856 228754 246908 228760
rect 246764 227248 246816 227254
rect 246764 227190 246816 227196
rect 246776 224954 246804 227190
rect 246776 224926 246896 224954
rect 245844 217864 245896 217870
rect 245844 217806 245896 217812
rect 245752 208344 245804 208350
rect 245752 208286 245804 208292
rect 245672 16546 245976 16574
rect 245212 480 245240 3454
rect 245568 3460 245620 3466
rect 245568 3402 245620 3408
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 246868 3670 246896 224926
rect 246856 3664 246908 3670
rect 246856 3606 246908 3612
rect 246960 3602 246988 236710
rect 247052 228886 247080 239634
rect 247144 234054 247172 239788
rect 247236 239788 247310 239816
rect 247420 239822 247494 239850
rect 247132 234048 247184 234054
rect 247132 233990 247184 233996
rect 247040 228880 247092 228886
rect 247040 228822 247092 228828
rect 247040 226840 247092 226846
rect 247040 226782 247092 226788
rect 247052 16574 247080 226782
rect 247236 224954 247264 239788
rect 247420 239714 247448 239822
rect 247650 239816 247678 240108
rect 247604 239788 247678 239816
rect 247420 239686 247540 239714
rect 247408 239624 247460 239630
rect 247408 239566 247460 239572
rect 247316 239284 247368 239290
rect 247316 239226 247368 239232
rect 247328 227186 247356 239226
rect 247420 238882 247448 239566
rect 247408 238876 247460 238882
rect 247408 238818 247460 238824
rect 247408 238740 247460 238746
rect 247408 238682 247460 238688
rect 247420 233102 247448 238682
rect 247512 234394 247540 239686
rect 247604 238746 247632 239788
rect 247742 239612 247770 240108
rect 247834 239873 247862 240108
rect 247820 239864 247876 239873
rect 247926 239850 247954 240108
rect 248018 239970 248046 240108
rect 248110 239970 248138 240108
rect 248006 239964 248058 239970
rect 248006 239906 248058 239912
rect 248098 239964 248150 239970
rect 248098 239906 248150 239912
rect 247926 239822 248092 239850
rect 247820 239799 247876 239808
rect 247868 239760 247920 239766
rect 247866 239728 247868 239737
rect 247960 239760 248012 239766
rect 247920 239728 247922 239737
rect 248064 239737 248092 239822
rect 247960 239702 248012 239708
rect 248050 239728 248106 239737
rect 247866 239663 247922 239672
rect 247696 239584 247770 239612
rect 247592 238740 247644 238746
rect 247592 238682 247644 238688
rect 247500 234388 247552 234394
rect 247500 234330 247552 234336
rect 247408 233096 247460 233102
rect 247408 233038 247460 233044
rect 247696 228954 247724 239584
rect 247880 239170 247908 239663
rect 247972 239358 248000 239702
rect 248202 239714 248230 240108
rect 248050 239663 248106 239672
rect 248156 239686 248230 239714
rect 248052 239624 248104 239630
rect 248052 239566 248104 239572
rect 248064 239465 248092 239566
rect 248050 239456 248106 239465
rect 248050 239391 248106 239400
rect 247960 239352 248012 239358
rect 247960 239294 248012 239300
rect 248156 239290 248184 239686
rect 248294 239612 248322 240108
rect 248386 239850 248414 240108
rect 248478 239970 248506 240108
rect 248466 239964 248518 239970
rect 248466 239906 248518 239912
rect 248570 239850 248598 240108
rect 248662 239970 248690 240108
rect 248650 239964 248702 239970
rect 248650 239906 248702 239912
rect 248386 239822 248460 239850
rect 248248 239584 248322 239612
rect 248248 239290 248276 239584
rect 248328 239488 248380 239494
rect 248328 239430 248380 239436
rect 248144 239284 248196 239290
rect 248144 239226 248196 239232
rect 248236 239284 248288 239290
rect 248236 239226 248288 239232
rect 247880 239142 248276 239170
rect 248052 238876 248104 238882
rect 248052 238818 248104 238824
rect 248064 231606 248092 238818
rect 248052 231600 248104 231606
rect 248052 231542 248104 231548
rect 247684 228948 247736 228954
rect 247684 228890 247736 228896
rect 247316 227180 247368 227186
rect 247316 227122 247368 227128
rect 247236 224926 248184 224954
rect 248156 211070 248184 224926
rect 248248 217326 248276 239142
rect 248340 235994 248368 239430
rect 248432 238649 248460 239822
rect 248524 239822 248598 239850
rect 248418 238640 248474 238649
rect 248418 238575 248474 238584
rect 248524 238542 248552 239822
rect 248754 239816 248782 240108
rect 248708 239788 248782 239816
rect 248604 239760 248656 239766
rect 248604 239702 248656 239708
rect 248616 238649 248644 239702
rect 248602 238640 248658 238649
rect 248602 238575 248658 238584
rect 248512 238536 248564 238542
rect 248512 238478 248564 238484
rect 248708 235994 248736 239788
rect 248846 239748 248874 240108
rect 248938 239970 248966 240108
rect 249030 239970 249058 240108
rect 248926 239964 248978 239970
rect 248926 239906 248978 239912
rect 249018 239964 249070 239970
rect 249018 239906 249070 239912
rect 248972 239828 249024 239834
rect 249122 239816 249150 240108
rect 249214 239850 249242 240108
rect 249306 239970 249334 240108
rect 249398 239970 249426 240108
rect 249294 239964 249346 239970
rect 249294 239906 249346 239912
rect 249386 239964 249438 239970
rect 249386 239906 249438 239912
rect 249490 239850 249518 240108
rect 249214 239822 249288 239850
rect 248972 239770 249024 239776
rect 249076 239788 249150 239816
rect 248340 235966 248460 235994
rect 248328 232348 248380 232354
rect 248328 232290 248380 232296
rect 248236 217320 248288 217326
rect 248236 217262 248288 217268
rect 248144 211064 248196 211070
rect 248144 211006 248196 211012
rect 247052 16546 247632 16574
rect 246948 3596 247000 3602
rect 246948 3538 247000 3544
rect 247604 480 247632 16546
rect 248340 4146 248368 232290
rect 248432 230178 248460 235966
rect 248616 235966 248736 235994
rect 248800 239720 248874 239748
rect 248800 235994 248828 239720
rect 248880 239624 248932 239630
rect 248878 239592 248880 239601
rect 248932 239592 248934 239601
rect 248878 239527 248934 239536
rect 248880 239488 248932 239494
rect 248880 239430 248932 239436
rect 248892 239086 248920 239430
rect 248880 239080 248932 239086
rect 248880 239022 248932 239028
rect 248800 235966 248920 235994
rect 248420 230172 248472 230178
rect 248420 230114 248472 230120
rect 248616 225894 248644 235966
rect 248892 231742 248920 235966
rect 248880 231736 248932 231742
rect 248880 231678 248932 231684
rect 248604 225888 248656 225894
rect 248604 225830 248656 225836
rect 248984 224954 249012 239770
rect 249076 239494 249104 239788
rect 249260 239737 249288 239822
rect 249352 239822 249518 239850
rect 249246 239728 249302 239737
rect 249246 239663 249302 239672
rect 249248 239556 249300 239562
rect 249248 239498 249300 239504
rect 249064 239488 249116 239494
rect 249064 239430 249116 239436
rect 249156 239352 249208 239358
rect 249156 239294 249208 239300
rect 249064 238604 249116 238610
rect 249064 238546 249116 238552
rect 249076 237522 249104 238546
rect 249064 237516 249116 237522
rect 249064 237458 249116 237464
rect 249168 228614 249196 239294
rect 249260 229022 249288 239498
rect 249352 239465 249380 239822
rect 249582 239748 249610 240108
rect 249674 239902 249702 240108
rect 249662 239896 249714 239902
rect 249766 239873 249794 240108
rect 249662 239838 249714 239844
rect 249752 239864 249808 239873
rect 249752 239799 249808 239808
rect 249858 239748 249886 240108
rect 249444 239720 249610 239748
rect 249720 239720 249886 239748
rect 249950 239748 249978 240108
rect 250042 239816 250070 240108
rect 250134 239970 250162 240108
rect 250122 239964 250174 239970
rect 250122 239906 250174 239912
rect 250042 239788 250116 239816
rect 249950 239720 250024 239748
rect 249338 239456 249394 239465
rect 249338 239391 249394 239400
rect 249340 239284 249392 239290
rect 249340 239226 249392 239232
rect 249352 237114 249380 239226
rect 249340 237108 249392 237114
rect 249340 237050 249392 237056
rect 249444 234614 249472 239720
rect 249522 239592 249578 239601
rect 249522 239527 249578 239536
rect 249352 234586 249472 234614
rect 249248 229016 249300 229022
rect 249248 228958 249300 228964
rect 249156 228608 249208 228614
rect 249156 228550 249208 228556
rect 248524 224926 249012 224954
rect 248524 223514 248552 224926
rect 248512 223508 248564 223514
rect 248512 223450 248564 223456
rect 249352 216646 249380 234586
rect 249536 224954 249564 239527
rect 249616 239420 249668 239426
rect 249616 239362 249668 239368
rect 249628 238610 249656 239362
rect 249616 238604 249668 238610
rect 249616 238546 249668 238552
rect 249720 238066 249748 239720
rect 249800 239624 249852 239630
rect 249800 239566 249852 239572
rect 249708 238060 249760 238066
rect 249708 238002 249760 238008
rect 249708 237652 249760 237658
rect 249708 237594 249760 237600
rect 249614 236192 249670 236201
rect 249614 236127 249670 236136
rect 249444 224926 249564 224954
rect 249340 216640 249392 216646
rect 249340 216582 249392 216588
rect 249444 196654 249472 224926
rect 249524 224256 249576 224262
rect 249524 224198 249576 224204
rect 249432 196648 249484 196654
rect 249432 196590 249484 196596
rect 248328 4140 248380 4146
rect 248328 4082 248380 4088
rect 249536 3398 249564 224198
rect 249628 7614 249656 236127
rect 249720 233442 249748 237594
rect 249708 233436 249760 233442
rect 249708 233378 249760 233384
rect 249616 7608 249668 7614
rect 249616 7550 249668 7556
rect 249720 3806 249748 233378
rect 249812 233170 249840 239566
rect 249996 237912 250024 239720
rect 250088 239465 250116 239788
rect 250226 239748 250254 240108
rect 250318 239970 250346 240108
rect 250410 239970 250438 240108
rect 250306 239964 250358 239970
rect 250306 239906 250358 239912
rect 250398 239964 250450 239970
rect 250398 239906 250450 239912
rect 250502 239748 250530 240108
rect 250594 239970 250622 240108
rect 250686 239970 250714 240108
rect 250582 239964 250634 239970
rect 250582 239906 250634 239912
rect 250674 239964 250726 239970
rect 250674 239906 250726 239912
rect 250628 239828 250680 239834
rect 250628 239770 250680 239776
rect 250180 239720 250254 239748
rect 250350 239728 250406 239737
rect 250074 239456 250130 239465
rect 250074 239391 250130 239400
rect 250180 239018 250208 239720
rect 250350 239663 250352 239672
rect 250404 239663 250406 239672
rect 250456 239720 250530 239748
rect 250352 239634 250404 239640
rect 250260 239624 250312 239630
rect 250260 239566 250312 239572
rect 250168 239012 250220 239018
rect 250168 238954 250220 238960
rect 250168 238060 250220 238066
rect 250168 238002 250220 238008
rect 249996 237884 250116 237912
rect 249984 237380 250036 237386
rect 249984 237322 250036 237328
rect 249892 236156 249944 236162
rect 249892 236098 249944 236104
rect 249800 233164 249852 233170
rect 249800 233106 249852 233112
rect 249904 229786 249932 236098
rect 249812 229758 249932 229786
rect 249812 220794 249840 229758
rect 249996 229650 250024 237322
rect 249904 229622 250024 229650
rect 249904 222154 249932 229622
rect 250088 228206 250116 237884
rect 250180 231810 250208 238002
rect 250168 231804 250220 231810
rect 250168 231746 250220 231752
rect 250076 228200 250128 228206
rect 250076 228142 250128 228148
rect 250272 224954 250300 239566
rect 250456 239290 250484 239720
rect 250536 239624 250588 239630
rect 250536 239566 250588 239572
rect 250444 239284 250496 239290
rect 250444 239226 250496 239232
rect 250444 239012 250496 239018
rect 250444 238954 250496 238960
rect 250352 238808 250404 238814
rect 250352 238750 250404 238756
rect 250364 236162 250392 238750
rect 250456 238678 250484 238954
rect 250444 238672 250496 238678
rect 250444 238614 250496 238620
rect 250444 238536 250496 238542
rect 250444 238478 250496 238484
rect 250352 236156 250404 236162
rect 250352 236098 250404 236104
rect 250456 227662 250484 238478
rect 250548 237969 250576 239566
rect 250640 238898 250668 239770
rect 250778 239748 250806 240108
rect 250870 239873 250898 240108
rect 250962 239902 250990 240108
rect 250950 239896 251002 239902
rect 250856 239864 250912 239873
rect 250950 239838 251002 239844
rect 250856 239799 250912 239808
rect 250904 239760 250956 239766
rect 250778 239720 250852 239748
rect 250720 239624 250772 239630
rect 250720 239566 250772 239572
rect 250732 239086 250760 239566
rect 250720 239080 250772 239086
rect 250720 239022 250772 239028
rect 250640 238870 250760 238898
rect 250628 238740 250680 238746
rect 250628 238682 250680 238688
rect 250534 237960 250590 237969
rect 250534 237895 250590 237904
rect 250548 235994 250576 237895
rect 250640 237289 250668 238682
rect 250732 237386 250760 238870
rect 250824 238746 250852 239720
rect 251054 239714 251082 240108
rect 251146 239970 251174 240108
rect 251238 239970 251266 240108
rect 251134 239964 251186 239970
rect 251134 239906 251186 239912
rect 251226 239964 251278 239970
rect 251226 239906 251278 239912
rect 251330 239902 251358 240108
rect 251318 239896 251370 239902
rect 251422 239873 251450 240108
rect 251318 239838 251370 239844
rect 251408 239864 251464 239873
rect 251408 239799 251464 239808
rect 250904 239702 250956 239708
rect 250916 238814 250944 239702
rect 251008 239686 251082 239714
rect 251180 239760 251232 239766
rect 251514 239748 251542 240108
rect 251606 239902 251634 240108
rect 251698 239902 251726 240108
rect 251790 239970 251818 240108
rect 251778 239964 251830 239970
rect 251778 239906 251830 239912
rect 251594 239896 251646 239902
rect 251594 239838 251646 239844
rect 251686 239896 251738 239902
rect 251686 239838 251738 239844
rect 251882 239816 251910 240108
rect 251974 239873 252002 240108
rect 252066 239902 252094 240108
rect 252158 239902 252186 240108
rect 252250 239970 252278 240108
rect 252342 239970 252370 240108
rect 252238 239964 252290 239970
rect 252238 239906 252290 239912
rect 252330 239964 252382 239970
rect 252330 239906 252382 239912
rect 252054 239896 252106 239902
rect 251790 239788 251910 239816
rect 251960 239864 252016 239873
rect 252054 239838 252106 239844
rect 252146 239896 252198 239902
rect 252146 239838 252198 239844
rect 252434 239834 252462 240108
rect 251960 239799 252016 239808
rect 252422 239828 252474 239834
rect 251790 239748 251818 239788
rect 252526 239816 252554 240108
rect 252618 239970 252646 240108
rect 252710 239970 252738 240108
rect 252606 239964 252658 239970
rect 252606 239906 252658 239912
rect 252698 239964 252750 239970
rect 252698 239906 252750 239912
rect 252802 239902 252830 240108
rect 252790 239896 252842 239902
rect 252790 239838 252842 239844
rect 252526 239788 252600 239816
rect 252422 239770 252474 239776
rect 251180 239702 251232 239708
rect 251468 239720 251542 239748
rect 251744 239720 251818 239748
rect 252008 239760 252060 239766
rect 250904 238808 250956 238814
rect 250904 238750 250956 238756
rect 250812 238740 250864 238746
rect 250812 238682 250864 238688
rect 250904 238672 250956 238678
rect 250904 238614 250956 238620
rect 250720 237380 250772 237386
rect 250720 237322 250772 237328
rect 250626 237280 250682 237289
rect 250626 237215 250682 237224
rect 250810 236192 250866 236201
rect 250810 236127 250866 236136
rect 250548 235966 250668 235994
rect 250444 227656 250496 227662
rect 250444 227598 250496 227604
rect 250640 227202 250668 235966
rect 250824 231854 250852 236127
rect 250916 235822 250944 238614
rect 251008 237046 251036 239686
rect 251088 239624 251140 239630
rect 251088 239566 251140 239572
rect 251100 238649 251128 239566
rect 251086 238640 251142 238649
rect 251086 238575 251142 238584
rect 250996 237040 251048 237046
rect 250996 236982 251048 236988
rect 250904 235816 250956 235822
rect 250904 235758 250956 235764
rect 251192 234938 251220 239702
rect 251364 239624 251416 239630
rect 251364 239566 251416 239572
rect 251272 239556 251324 239562
rect 251272 239498 251324 239504
rect 251284 238814 251312 239498
rect 251272 238808 251324 238814
rect 251272 238750 251324 238756
rect 251180 234932 251232 234938
rect 251180 234874 251232 234880
rect 251180 233028 251232 233034
rect 251180 232970 251232 232976
rect 251088 232552 251140 232558
rect 251088 232494 251140 232500
rect 250824 231826 251036 231854
rect 250640 227174 250944 227202
rect 250812 227112 250864 227118
rect 250812 227054 250864 227060
rect 249996 224926 250300 224954
rect 249996 224602 250024 224926
rect 249984 224596 250036 224602
rect 249984 224538 250036 224544
rect 249892 222148 249944 222154
rect 249892 222090 249944 222096
rect 249800 220788 249852 220794
rect 249800 220730 249852 220736
rect 250824 195294 250852 227054
rect 250812 195288 250864 195294
rect 250812 195230 250864 195236
rect 250916 164898 250944 227174
rect 251008 227118 251036 231826
rect 250996 227112 251048 227118
rect 250996 227054 251048 227060
rect 250994 226264 251050 226273
rect 250994 226199 251050 226208
rect 251008 223310 251036 226199
rect 250996 223304 251048 223310
rect 250996 223246 251048 223252
rect 250904 164892 250956 164898
rect 250904 164834 250956 164840
rect 251008 8974 251036 223246
rect 250996 8968 251048 8974
rect 250996 8910 251048 8916
rect 249984 4140 250036 4146
rect 249984 4082 250036 4088
rect 249708 3800 249760 3806
rect 249708 3742 249760 3748
rect 249524 3392 249576 3398
rect 249524 3334 249576 3340
rect 248788 3256 248840 3262
rect 248788 3198 248840 3204
rect 248800 480 248828 3198
rect 249996 480 250024 4082
rect 251100 4078 251128 232494
rect 251192 232490 251220 232970
rect 251180 232484 251232 232490
rect 251180 232426 251232 232432
rect 251376 231674 251404 239566
rect 251364 231668 251416 231674
rect 251364 231610 251416 231616
rect 251468 230314 251496 239720
rect 251640 239692 251692 239698
rect 251640 239634 251692 239640
rect 251652 239601 251680 239634
rect 251638 239592 251694 239601
rect 251548 239556 251600 239562
rect 251638 239527 251694 239536
rect 251548 239498 251600 239504
rect 251560 235958 251588 239498
rect 251640 239420 251692 239426
rect 251640 239362 251692 239368
rect 251652 238882 251680 239362
rect 251744 238898 251772 239720
rect 252008 239702 252060 239708
rect 251916 239556 251968 239562
rect 251916 239498 251968 239504
rect 251640 238876 251692 238882
rect 251744 238870 251864 238898
rect 251640 238818 251692 238824
rect 251732 238740 251784 238746
rect 251732 238682 251784 238688
rect 251744 235994 251772 238682
rect 251652 235966 251772 235994
rect 251548 235952 251600 235958
rect 251548 235894 251600 235900
rect 251652 231854 251680 235966
rect 251836 235385 251864 238870
rect 251928 238746 251956 239498
rect 251916 238740 251968 238746
rect 251916 238682 251968 238688
rect 251916 237788 251968 237794
rect 251916 237730 251968 237736
rect 251822 235376 251878 235385
rect 251822 235311 251878 235320
rect 251652 231826 251772 231854
rect 251456 230308 251508 230314
rect 251456 230250 251508 230256
rect 251744 227730 251772 231826
rect 251928 228410 251956 237730
rect 251916 228404 251968 228410
rect 251916 228346 251968 228352
rect 251732 227724 251784 227730
rect 251732 227666 251784 227672
rect 252020 224954 252048 239702
rect 252284 239692 252336 239698
rect 252284 239634 252336 239640
rect 252376 239692 252428 239698
rect 252376 239634 252428 239640
rect 252192 239624 252244 239630
rect 252192 239566 252244 239572
rect 252100 239284 252152 239290
rect 252100 239226 252152 239232
rect 252112 233753 252140 239226
rect 252098 233744 252154 233753
rect 252098 233679 252154 233688
rect 252204 232218 252232 239566
rect 252192 232212 252244 232218
rect 252192 232154 252244 232160
rect 252296 231854 252324 239634
rect 252388 236162 252416 239634
rect 252466 239592 252522 239601
rect 252466 239527 252522 239536
rect 252376 236156 252428 236162
rect 252376 236098 252428 236104
rect 252376 232484 252428 232490
rect 252376 232426 252428 232432
rect 251284 224926 252048 224954
rect 252204 231826 252324 231854
rect 251284 223446 251312 224926
rect 251272 223440 251324 223446
rect 251272 223382 251324 223388
rect 252204 215218 252232 231826
rect 252282 221640 252338 221649
rect 252282 221575 252338 221584
rect 252192 215212 252244 215218
rect 252192 215154 252244 215160
rect 251272 162172 251324 162178
rect 251272 162114 251324 162120
rect 251284 16574 251312 162114
rect 251284 16546 252232 16574
rect 251088 4072 251140 4078
rect 251088 4014 251140 4020
rect 252204 3482 252232 16546
rect 252296 3942 252324 221575
rect 252284 3936 252336 3942
rect 252284 3878 252336 3884
rect 252388 3738 252416 232426
rect 252480 3874 252508 239527
rect 252572 239358 252600 239788
rect 252744 239760 252796 239766
rect 252650 239728 252706 239737
rect 252894 239748 252922 240108
rect 252744 239702 252796 239708
rect 252848 239720 252922 239748
rect 252986 239748 253014 240108
rect 253078 239902 253106 240108
rect 253066 239896 253118 239902
rect 253066 239838 253118 239844
rect 253170 239850 253198 240108
rect 253262 239970 253290 240108
rect 253250 239964 253302 239970
rect 253250 239906 253302 239912
rect 253354 239873 253382 240108
rect 253340 239864 253396 239873
rect 253170 239822 253244 239850
rect 253112 239760 253164 239766
rect 252986 239720 253060 239748
rect 252650 239663 252652 239672
rect 252704 239663 252706 239672
rect 252652 239634 252704 239640
rect 252560 239352 252612 239358
rect 252560 239294 252612 239300
rect 252560 239216 252612 239222
rect 252560 239158 252612 239164
rect 252650 239184 252706 239193
rect 252572 237862 252600 239158
rect 252650 239119 252706 239128
rect 252560 237856 252612 237862
rect 252560 237798 252612 237804
rect 252664 6458 252692 239119
rect 252756 226166 252784 239702
rect 252848 228682 252876 239720
rect 252926 239592 252982 239601
rect 252926 239527 252982 239536
rect 252940 236026 252968 239527
rect 253032 236434 253060 239720
rect 253110 239728 253112 239737
rect 253164 239728 253166 239737
rect 253110 239663 253166 239672
rect 253216 239680 253244 239822
rect 253340 239799 253396 239808
rect 253446 239816 253474 240108
rect 253538 239970 253566 240108
rect 253630 239970 253658 240108
rect 253526 239964 253578 239970
rect 253526 239906 253578 239912
rect 253618 239964 253670 239970
rect 253618 239906 253670 239912
rect 253722 239816 253750 240108
rect 253814 239970 253842 240108
rect 253906 239970 253934 240108
rect 253802 239964 253854 239970
rect 253802 239906 253854 239912
rect 253894 239964 253946 239970
rect 253894 239906 253946 239912
rect 253446 239788 253612 239816
rect 253722 239788 253888 239816
rect 253388 239692 253440 239698
rect 253216 239652 253336 239680
rect 253112 239624 253164 239630
rect 253112 239566 253164 239572
rect 253124 238649 253152 239566
rect 253204 239488 253256 239494
rect 253204 239430 253256 239436
rect 253216 238678 253244 239430
rect 253308 238762 253336 239652
rect 253388 239634 253440 239640
rect 253400 239601 253428 239634
rect 253480 239624 253532 239630
rect 253386 239592 253442 239601
rect 253480 239566 253532 239572
rect 253386 239527 253442 239536
rect 253388 239352 253440 239358
rect 253388 239294 253440 239300
rect 253400 238882 253428 239294
rect 253492 239193 253520 239566
rect 253478 239184 253534 239193
rect 253478 239119 253534 239128
rect 253388 238876 253440 238882
rect 253388 238818 253440 238824
rect 253308 238734 253520 238762
rect 253204 238672 253256 238678
rect 253110 238640 253166 238649
rect 253204 238614 253256 238620
rect 253110 238575 253166 238584
rect 253388 238604 253440 238610
rect 253388 238546 253440 238552
rect 253020 236428 253072 236434
rect 253020 236370 253072 236376
rect 252928 236020 252980 236026
rect 252928 235962 252980 235968
rect 253204 235952 253256 235958
rect 253204 235894 253256 235900
rect 252836 228676 252888 228682
rect 252836 228618 252888 228624
rect 253216 227225 253244 235894
rect 253400 234614 253428 238546
rect 253308 234586 253428 234614
rect 253308 228478 253336 234586
rect 253296 228472 253348 228478
rect 253296 228414 253348 228420
rect 253202 227216 253258 227225
rect 253202 227151 253258 227160
rect 252744 226160 252796 226166
rect 252744 226102 252796 226108
rect 253492 218958 253520 238734
rect 253480 218952 253532 218958
rect 253480 218894 253532 218900
rect 253204 214600 253256 214606
rect 253204 214542 253256 214548
rect 252652 6452 252704 6458
rect 252652 6394 252704 6400
rect 252468 3868 252520 3874
rect 252468 3810 252520 3816
rect 252376 3732 252428 3738
rect 252376 3674 252428 3680
rect 252204 3454 252416 3482
rect 251180 3392 251232 3398
rect 251180 3334 251232 3340
rect 251192 480 251220 3334
rect 252388 480 252416 3454
rect 253216 3398 253244 214542
rect 253584 213926 253612 239788
rect 253754 239728 253810 239737
rect 253664 239692 253716 239698
rect 253754 239663 253756 239672
rect 253664 239634 253716 239640
rect 253808 239663 253810 239672
rect 253756 239634 253808 239640
rect 253676 236502 253704 239634
rect 253754 239592 253810 239601
rect 253754 239527 253810 239536
rect 253664 236496 253716 236502
rect 253664 236438 253716 236444
rect 253662 228712 253718 228721
rect 253662 228647 253718 228656
rect 253572 213920 253624 213926
rect 253572 213862 253624 213868
rect 253676 3738 253704 228647
rect 253768 224954 253796 239527
rect 253860 233209 253888 239788
rect 253998 239748 254026 240108
rect 254090 239902 254118 240108
rect 254078 239896 254130 239902
rect 254182 239873 254210 240108
rect 254078 239838 254130 239844
rect 254168 239864 254224 239873
rect 254168 239799 254224 239808
rect 254274 239816 254302 240108
rect 254366 239970 254394 240108
rect 254354 239964 254406 239970
rect 254354 239906 254406 239912
rect 254458 239902 254486 240108
rect 254446 239896 254498 239902
rect 254550 239873 254578 240108
rect 254642 239902 254670 240108
rect 254630 239896 254682 239902
rect 254446 239838 254498 239844
rect 254536 239864 254592 239873
rect 254274 239788 254348 239816
rect 254630 239838 254682 239844
rect 254734 239850 254762 240108
rect 254826 239970 254854 240108
rect 254918 239970 254946 240108
rect 254814 239964 254866 239970
rect 254814 239906 254866 239912
rect 254906 239964 254958 239970
rect 254906 239906 254958 239912
rect 254734 239822 254808 239850
rect 254536 239799 254592 239808
rect 253998 239720 254072 239748
rect 253940 239148 253992 239154
rect 253940 239090 253992 239096
rect 253952 237998 253980 239090
rect 253940 237992 253992 237998
rect 253940 237934 253992 237940
rect 253940 235952 253992 235958
rect 253940 235894 253992 235900
rect 253952 234938 253980 235894
rect 253940 234932 253992 234938
rect 253940 234874 253992 234880
rect 254044 234190 254072 239720
rect 254124 239692 254176 239698
rect 254124 239634 254176 239640
rect 254216 239692 254268 239698
rect 254216 239634 254268 239640
rect 254136 234614 254164 239634
rect 254228 239086 254256 239634
rect 254216 239080 254268 239086
rect 254216 239022 254268 239028
rect 254136 234586 254256 234614
rect 254032 234184 254084 234190
rect 254032 234126 254084 234132
rect 253846 233200 253902 233209
rect 253846 233135 253902 233144
rect 254124 229492 254176 229498
rect 254124 229434 254176 229440
rect 254032 229424 254084 229430
rect 254032 229366 254084 229372
rect 253940 229220 253992 229226
rect 253940 229162 253992 229168
rect 253768 224926 253888 224954
rect 253860 6390 253888 224926
rect 253952 211138 253980 229162
rect 254044 218006 254072 229366
rect 254136 221950 254164 229434
rect 254228 226030 254256 234586
rect 254320 230518 254348 239788
rect 254780 239714 254808 239822
rect 254860 239828 254912 239834
rect 255010 239816 255038 240108
rect 254860 239770 254912 239776
rect 254964 239788 255038 239816
rect 254492 239692 254544 239698
rect 254412 239652 254492 239680
rect 254308 230512 254360 230518
rect 254308 230454 254360 230460
rect 254216 226024 254268 226030
rect 254216 225966 254268 225972
rect 254412 222834 254440 239652
rect 254492 239634 254544 239640
rect 254688 239686 254808 239714
rect 254582 239592 254638 239601
rect 254582 239527 254638 239536
rect 254492 238808 254544 238814
rect 254492 238750 254544 238756
rect 254504 233034 254532 238750
rect 254492 233028 254544 233034
rect 254492 232970 254544 232976
rect 254596 229498 254624 239527
rect 254688 235929 254716 239686
rect 254768 239624 254820 239630
rect 254768 239566 254820 239572
rect 254780 237658 254808 239566
rect 254768 237652 254820 237658
rect 254768 237594 254820 237600
rect 254768 237516 254820 237522
rect 254768 237458 254820 237464
rect 254674 235920 254730 235929
rect 254674 235855 254730 235864
rect 254780 234614 254808 237458
rect 254688 234586 254808 234614
rect 254584 229492 254636 229498
rect 254584 229434 254636 229440
rect 254688 228342 254716 234586
rect 254768 230512 254820 230518
rect 254768 230454 254820 230460
rect 254676 228336 254728 228342
rect 254676 228278 254728 228284
rect 254780 224942 254808 230454
rect 254872 229430 254900 239770
rect 254964 236065 254992 239788
rect 255102 239748 255130 240108
rect 255194 239873 255222 240108
rect 255286 239970 255314 240108
rect 255274 239964 255326 239970
rect 255274 239906 255326 239912
rect 255378 239902 255406 240108
rect 255470 239970 255498 240108
rect 255458 239964 255510 239970
rect 255458 239906 255510 239912
rect 255562 239902 255590 240108
rect 255366 239896 255418 239902
rect 255180 239864 255236 239873
rect 255366 239838 255418 239844
rect 255550 239896 255602 239902
rect 255550 239838 255602 239844
rect 255180 239799 255236 239808
rect 255102 239720 255176 239748
rect 255044 239624 255096 239630
rect 255042 239592 255044 239601
rect 255096 239592 255098 239601
rect 255042 239527 255098 239536
rect 255042 239456 255098 239465
rect 255042 239391 255098 239400
rect 255056 239290 255084 239391
rect 255044 239284 255096 239290
rect 255044 239226 255096 239232
rect 254950 236056 255006 236065
rect 254950 235991 255006 236000
rect 254860 229424 254912 229430
rect 254860 229366 254912 229372
rect 255148 229226 255176 239720
rect 255226 239728 255282 239737
rect 255654 239714 255682 240108
rect 255746 239902 255774 240108
rect 255838 239970 255866 240108
rect 255930 239970 255958 240108
rect 256022 239970 256050 240108
rect 256114 239970 256142 240108
rect 255826 239964 255878 239970
rect 255826 239906 255878 239912
rect 255918 239964 255970 239970
rect 255918 239906 255970 239912
rect 256010 239964 256062 239970
rect 256010 239906 256062 239912
rect 256102 239964 256154 239970
rect 256102 239906 256154 239912
rect 255734 239896 255786 239902
rect 255734 239838 255786 239844
rect 256206 239816 256234 240108
rect 256298 239850 256326 240108
rect 256390 239970 256418 240108
rect 256378 239964 256430 239970
rect 256378 239906 256430 239912
rect 256298 239822 256372 239850
rect 256160 239788 256234 239816
rect 255654 239686 255728 239714
rect 255226 239663 255282 239672
rect 255240 238134 255268 239663
rect 255504 239624 255556 239630
rect 255596 239624 255648 239630
rect 255504 239566 255556 239572
rect 255594 239592 255596 239601
rect 255648 239592 255650 239601
rect 255320 239556 255372 239562
rect 255320 239498 255372 239504
rect 255228 238128 255280 238134
rect 255228 238070 255280 238076
rect 255226 237960 255282 237969
rect 255226 237895 255282 237904
rect 255136 229220 255188 229226
rect 255136 229162 255188 229168
rect 254768 224936 254820 224942
rect 254768 224878 254820 224884
rect 255134 223816 255190 223825
rect 255134 223751 255190 223760
rect 255148 223106 255176 223751
rect 255136 223100 255188 223106
rect 255136 223042 255188 223048
rect 255148 222986 255176 223042
rect 255056 222958 255176 222986
rect 254400 222828 254452 222834
rect 254400 222770 254452 222776
rect 254124 221944 254176 221950
rect 254124 221886 254176 221892
rect 254032 218000 254084 218006
rect 254032 217942 254084 217948
rect 253940 211132 253992 211138
rect 253940 211074 253992 211080
rect 255056 189786 255084 222958
rect 255136 222828 255188 222834
rect 255136 222770 255188 222776
rect 255044 189780 255096 189786
rect 255044 189722 255096 189728
rect 255148 171834 255176 222770
rect 255136 171828 255188 171834
rect 255136 171770 255188 171776
rect 255240 14482 255268 237895
rect 255332 237017 255360 239498
rect 255516 237969 255544 239566
rect 255594 239527 255650 239536
rect 255502 237960 255558 237969
rect 255502 237895 255558 237904
rect 255410 237688 255466 237697
rect 255410 237623 255466 237632
rect 255318 237008 255374 237017
rect 255318 236943 255374 236952
rect 255320 232212 255372 232218
rect 255320 232154 255372 232160
rect 255332 227322 255360 232154
rect 255320 227316 255372 227322
rect 255320 227258 255372 227264
rect 255424 220726 255452 237623
rect 255608 235994 255636 239527
rect 255700 236609 255728 239686
rect 255964 239692 256016 239698
rect 255964 239634 256016 239640
rect 255976 238066 256004 239634
rect 256056 239624 256108 239630
rect 256056 239566 256108 239572
rect 255964 238060 256016 238066
rect 255964 238002 256016 238008
rect 256068 237522 256096 239566
rect 256160 239465 256188 239788
rect 256344 239714 256372 239822
rect 256482 239816 256510 240108
rect 256574 239902 256602 240108
rect 256562 239896 256614 239902
rect 256666 239873 256694 240108
rect 256562 239838 256614 239844
rect 256652 239864 256708 239873
rect 256252 239686 256372 239714
rect 256436 239788 256510 239816
rect 256652 239799 256708 239808
rect 256146 239456 256202 239465
rect 256146 239391 256202 239400
rect 256252 239306 256280 239686
rect 256332 239624 256384 239630
rect 256330 239592 256332 239601
rect 256384 239592 256386 239601
rect 256330 239527 256386 239536
rect 256436 239306 256464 239788
rect 256758 239748 256786 240108
rect 256850 239850 256878 240108
rect 256942 239970 256970 240108
rect 257034 239970 257062 240108
rect 256930 239964 256982 239970
rect 256930 239906 256982 239912
rect 257022 239964 257074 239970
rect 257022 239906 257074 239912
rect 257126 239902 257154 240108
rect 257114 239896 257166 239902
rect 256850 239822 256924 239850
rect 257114 239838 257166 239844
rect 256514 239728 256570 239737
rect 256758 239720 256832 239748
rect 256514 239663 256570 239672
rect 256528 239562 256556 239663
rect 256516 239556 256568 239562
rect 256568 239516 256648 239544
rect 256516 239498 256568 239504
rect 256206 239278 256280 239306
rect 256344 239278 256464 239306
rect 256206 238626 256234 239278
rect 256344 239170 256372 239278
rect 256298 239142 256372 239170
rect 256424 239216 256476 239222
rect 256424 239158 256476 239164
rect 256298 238762 256326 239142
rect 256436 238950 256464 239158
rect 256424 238944 256476 238950
rect 256424 238886 256476 238892
rect 256298 238734 256372 238762
rect 256206 238598 256280 238626
rect 256252 238542 256280 238598
rect 256240 238536 256292 238542
rect 256240 238478 256292 238484
rect 256056 237516 256108 237522
rect 256056 237458 256108 237464
rect 255686 236600 255742 236609
rect 255686 236535 255742 236544
rect 255964 236564 256016 236570
rect 255964 236506 256016 236512
rect 255608 235966 255820 235994
rect 255792 229498 255820 235966
rect 255780 229492 255832 229498
rect 255780 229434 255832 229440
rect 255976 228546 256004 236506
rect 256148 236020 256200 236026
rect 256148 235962 256200 235968
rect 255964 228540 256016 228546
rect 255964 228482 256016 228488
rect 256160 225826 256188 235962
rect 256148 225820 256200 225826
rect 256148 225762 256200 225768
rect 256344 224954 256372 238734
rect 256424 238060 256476 238066
rect 256424 238002 256476 238008
rect 256516 238060 256568 238066
rect 256516 238002 256568 238008
rect 255516 224926 256372 224954
rect 255516 223582 255544 224926
rect 255504 223576 255556 223582
rect 255504 223518 255556 223524
rect 255412 220720 255464 220726
rect 255412 220662 255464 220668
rect 256436 220522 256464 238002
rect 256528 235890 256556 238002
rect 256516 235884 256568 235890
rect 256516 235826 256568 235832
rect 256516 229492 256568 229498
rect 256516 229434 256568 229440
rect 256424 220516 256476 220522
rect 256424 220458 256476 220464
rect 255320 33788 255372 33794
rect 255320 33730 255372 33736
rect 255332 16574 255360 33730
rect 255332 16546 255912 16574
rect 255228 14476 255280 14482
rect 255228 14418 255280 14424
rect 253848 6384 253900 6390
rect 253848 6326 253900 6332
rect 253480 3732 253532 3738
rect 253480 3674 253532 3680
rect 253664 3732 253716 3738
rect 253664 3674 253716 3680
rect 253204 3392 253256 3398
rect 253204 3334 253256 3340
rect 253492 480 253520 3674
rect 254676 3392 254728 3398
rect 254676 3334 254728 3340
rect 254688 480 254716 3334
rect 255884 480 255912 16546
rect 256528 6322 256556 229434
rect 256516 6316 256568 6322
rect 256516 6258 256568 6264
rect 256620 6254 256648 239516
rect 256700 239488 256752 239494
rect 256700 239430 256752 239436
rect 256712 236638 256740 239430
rect 256700 236632 256752 236638
rect 256700 236574 256752 236580
rect 256804 236570 256832 239720
rect 256896 237794 256924 239822
rect 256976 239828 257028 239834
rect 256976 239770 257028 239776
rect 256988 239737 257016 239770
rect 257068 239760 257120 239766
rect 256974 239728 257030 239737
rect 257218 239714 257246 240108
rect 257068 239702 257120 239708
rect 256974 239663 257030 239672
rect 256976 239624 257028 239630
rect 256976 239566 257028 239572
rect 256884 237788 256936 237794
rect 256884 237730 256936 237736
rect 256884 237652 256936 237658
rect 256884 237594 256936 237600
rect 256792 236564 256844 236570
rect 256792 236506 256844 236512
rect 256792 236428 256844 236434
rect 256792 236370 256844 236376
rect 256804 233889 256832 236370
rect 256790 233880 256846 233889
rect 256790 233815 256846 233824
rect 256792 233368 256844 233374
rect 256792 233310 256844 233316
rect 256700 229492 256752 229498
rect 256700 229434 256752 229440
rect 256712 213858 256740 229434
rect 256804 215286 256832 233310
rect 256896 229090 256924 237594
rect 256884 229084 256936 229090
rect 256884 229026 256936 229032
rect 256988 225962 257016 239566
rect 257080 238066 257108 239702
rect 257172 239686 257246 239714
rect 257068 238060 257120 238066
rect 257068 238002 257120 238008
rect 257068 237924 257120 237930
rect 257068 237866 257120 237872
rect 257080 231130 257108 237866
rect 257172 235249 257200 239686
rect 257310 239612 257338 240108
rect 257402 239902 257430 240108
rect 257494 239907 257522 240108
rect 257390 239896 257442 239902
rect 257390 239838 257442 239844
rect 257480 239898 257536 239907
rect 257480 239833 257536 239842
rect 257586 239680 257614 240108
rect 257540 239652 257614 239680
rect 257264 239584 257338 239612
rect 257436 239624 257488 239630
rect 257158 235240 257214 235249
rect 257158 235175 257214 235184
rect 257068 231124 257120 231130
rect 257068 231066 257120 231072
rect 256976 225956 257028 225962
rect 256976 225898 257028 225904
rect 257264 224954 257292 239584
rect 257436 239566 257488 239572
rect 257344 239420 257396 239426
rect 257344 239362 257396 239368
rect 257356 237998 257384 239362
rect 257344 237992 257396 237998
rect 257344 237934 257396 237940
rect 257448 234938 257476 239566
rect 257436 234932 257488 234938
rect 257436 234874 257488 234880
rect 257540 234682 257568 239652
rect 257678 239612 257706 240108
rect 257770 239970 257798 240108
rect 257862 239970 257890 240108
rect 257758 239964 257810 239970
rect 257758 239906 257810 239912
rect 257850 239964 257902 239970
rect 257850 239906 257902 239912
rect 257954 239907 257982 240108
rect 257940 239898 257996 239907
rect 258046 239902 258074 240108
rect 258138 239902 258166 240108
rect 258230 239907 258258 240108
rect 257940 239833 257996 239842
rect 258034 239896 258086 239902
rect 258034 239838 258086 239844
rect 258126 239896 258178 239902
rect 258126 239838 258178 239844
rect 258216 239898 258272 239907
rect 258322 239902 258350 240108
rect 258414 239902 258442 240108
rect 258216 239833 258272 239842
rect 258310 239896 258362 239902
rect 258310 239838 258362 239844
rect 258402 239896 258454 239902
rect 258402 239838 258454 239844
rect 257804 239760 257856 239766
rect 258356 239760 258408 239766
rect 257804 239702 257856 239708
rect 258078 239728 258134 239737
rect 257678 239584 257752 239612
rect 257620 239488 257672 239494
rect 257620 239430 257672 239436
rect 257448 234654 257568 234682
rect 257448 233374 257476 234654
rect 257632 234614 257660 239430
rect 257724 239086 257752 239584
rect 257712 239080 257764 239086
rect 257712 239022 257764 239028
rect 257540 234586 257660 234614
rect 257436 233368 257488 233374
rect 257436 233310 257488 233316
rect 257540 228585 257568 234586
rect 257816 230474 257844 239702
rect 257896 239692 257948 239698
rect 257896 239634 257948 239640
rect 257988 239692 258040 239698
rect 258078 239663 258134 239672
rect 258262 239728 258318 239737
rect 258506 239748 258534 240108
rect 258598 239873 258626 240108
rect 258690 239970 258718 240108
rect 258678 239964 258730 239970
rect 258678 239906 258730 239912
rect 258584 239864 258640 239873
rect 258584 239799 258640 239808
rect 258782 239816 258810 240108
rect 258874 239970 258902 240108
rect 258862 239964 258914 239970
rect 258862 239906 258914 239912
rect 258966 239850 258994 240108
rect 258920 239822 258994 239850
rect 258782 239788 258856 239816
rect 258460 239737 258534 239748
rect 258356 239702 258408 239708
rect 258446 239728 258534 239737
rect 258262 239663 258318 239672
rect 257988 239634 258040 239640
rect 257908 239601 257936 239634
rect 257894 239592 257950 239601
rect 257894 239527 257950 239536
rect 257724 230446 257844 230474
rect 257724 229498 257752 230446
rect 257712 229492 257764 229498
rect 257712 229434 257764 229440
rect 257526 228576 257582 228585
rect 257526 228511 257582 228520
rect 257908 224954 257936 239527
rect 258000 236745 258028 239634
rect 257986 236736 258042 236745
rect 257986 236671 258042 236680
rect 257988 236564 258040 236570
rect 257988 236506 258040 236512
rect 258000 229673 258028 236506
rect 258092 235793 258120 239663
rect 258078 235784 258134 235793
rect 258078 235719 258134 235728
rect 258172 235204 258224 235210
rect 258172 235146 258224 235152
rect 258184 229786 258212 235146
rect 258276 230466 258304 239663
rect 258368 235249 258396 239702
rect 258502 239720 258534 239728
rect 258446 239663 258502 239672
rect 258632 239692 258684 239698
rect 258632 239634 258684 239640
rect 258540 239624 258592 239630
rect 258540 239566 258592 239572
rect 258448 239556 258500 239562
rect 258448 239498 258500 239504
rect 258354 235240 258410 235249
rect 258460 235210 258488 239498
rect 258354 235175 258410 235184
rect 258448 235204 258500 235210
rect 258448 235146 258500 235152
rect 258276 230438 258488 230466
rect 258184 229758 258396 229786
rect 257986 229664 258042 229673
rect 257986 229599 258042 229608
rect 258264 229492 258316 229498
rect 258264 229434 258316 229440
rect 258080 229424 258132 229430
rect 258080 229366 258132 229372
rect 257264 224926 257844 224954
rect 257908 224926 258028 224954
rect 257816 223174 257844 224926
rect 257804 223168 257856 223174
rect 257804 223110 257856 223116
rect 256884 222964 256936 222970
rect 256884 222906 256936 222912
rect 256896 222834 256924 222906
rect 256884 222828 256936 222834
rect 256884 222770 256936 222776
rect 256792 215280 256844 215286
rect 256792 215222 256844 215228
rect 256700 213852 256752 213858
rect 256700 213794 256752 213800
rect 258000 149734 258028 224926
rect 258092 212430 258120 229366
rect 258172 229356 258224 229362
rect 258172 229298 258224 229304
rect 258080 212424 258132 212430
rect 258080 212366 258132 212372
rect 258078 204912 258134 204921
rect 258078 204847 258134 204856
rect 257988 149728 258040 149734
rect 257988 149670 258040 149676
rect 258092 16574 258120 204847
rect 258184 204270 258212 229298
rect 258276 205630 258304 229434
rect 258368 219366 258396 229758
rect 258460 226234 258488 230438
rect 258552 227390 258580 239566
rect 258644 229430 258672 239634
rect 258828 239494 258856 239788
rect 258816 239488 258868 239494
rect 258816 239430 258868 239436
rect 258814 239320 258870 239329
rect 258814 239255 258870 239264
rect 258828 238882 258856 239255
rect 258816 238876 258868 238882
rect 258816 238818 258868 238824
rect 258722 238096 258778 238105
rect 258722 238031 258778 238040
rect 258736 237862 258764 238031
rect 258724 237856 258776 237862
rect 258724 237798 258776 237804
rect 258724 236428 258776 236434
rect 258724 236370 258776 236376
rect 258736 236230 258764 236370
rect 258724 236224 258776 236230
rect 258724 236166 258776 236172
rect 258920 229498 258948 239822
rect 259058 239714 259086 240108
rect 259150 239873 259178 240108
rect 259136 239864 259192 239873
rect 259136 239799 259192 239808
rect 259242 239748 259270 240108
rect 259334 239816 259362 240108
rect 259426 239970 259454 240108
rect 259414 239964 259466 239970
rect 259414 239906 259466 239912
rect 259518 239850 259546 240108
rect 259610 239873 259638 240108
rect 259702 239970 259730 240108
rect 259690 239964 259742 239970
rect 259690 239906 259742 239912
rect 259794 239902 259822 240108
rect 259886 239970 259914 240108
rect 259874 239964 259926 239970
rect 259874 239906 259926 239912
rect 259978 239902 260006 240108
rect 259782 239896 259834 239902
rect 259472 239822 259546 239850
rect 259596 239864 259652 239873
rect 259334 239788 259408 239816
rect 259242 239720 259316 239748
rect 259012 239686 259086 239714
rect 259012 239193 259040 239686
rect 259092 239624 259144 239630
rect 259090 239592 259092 239601
rect 259184 239624 259236 239630
rect 259144 239592 259146 239601
rect 259184 239566 259236 239572
rect 259090 239527 259146 239536
rect 259196 239465 259224 239566
rect 259182 239456 259238 239465
rect 259182 239391 259238 239400
rect 258998 239184 259054 239193
rect 258998 239119 259054 239128
rect 259184 238808 259236 238814
rect 259184 238750 259236 238756
rect 259000 238536 259052 238542
rect 259000 238478 259052 238484
rect 259012 237402 259040 238478
rect 259012 237374 259132 237402
rect 259000 237040 259052 237046
rect 259000 236982 259052 236988
rect 259012 229945 259040 236982
rect 259104 230081 259132 237374
rect 259090 230072 259146 230081
rect 259090 230007 259146 230016
rect 258998 229936 259054 229945
rect 258998 229871 259054 229880
rect 258908 229492 258960 229498
rect 258908 229434 258960 229440
rect 258632 229424 258684 229430
rect 258632 229366 258684 229372
rect 259196 227594 259224 238750
rect 259288 229362 259316 239720
rect 259380 239698 259408 239788
rect 259472 239748 259500 239822
rect 259782 239838 259834 239844
rect 259966 239896 260018 239902
rect 259966 239838 260018 239844
rect 259596 239799 259652 239808
rect 259472 239720 259546 239748
rect 259518 239714 259546 239720
rect 259642 239728 259698 239737
rect 259368 239692 259420 239698
rect 259518 239686 259592 239714
rect 259368 239634 259420 239640
rect 259460 239556 259512 239562
rect 259460 239498 259512 239504
rect 259472 236881 259500 239498
rect 259458 236872 259514 236881
rect 259458 236807 259514 236816
rect 259276 229356 259328 229362
rect 259276 229298 259328 229304
rect 259184 227588 259236 227594
rect 259184 227530 259236 227536
rect 258540 227384 258592 227390
rect 258540 227326 258592 227332
rect 258448 226228 258500 226234
rect 258448 226170 258500 226176
rect 258356 219360 258408 219366
rect 258356 219302 258408 219308
rect 259366 218104 259422 218113
rect 259366 218039 259422 218048
rect 258264 205624 258316 205630
rect 258264 205566 258316 205572
rect 258172 204264 258224 204270
rect 258172 204206 258224 204212
rect 258092 16546 258304 16574
rect 256608 6248 256660 6254
rect 256608 6190 256660 6196
rect 257068 4004 257120 4010
rect 257068 3946 257120 3952
rect 257080 480 257108 3946
rect 258276 480 258304 16546
rect 259380 6186 259408 218039
rect 259564 211002 259592 239686
rect 259642 239663 259698 239672
rect 259736 239692 259788 239698
rect 259656 237153 259684 239663
rect 260070 239680 260098 240108
rect 260162 239714 260190 240108
rect 260254 239970 260282 240108
rect 260242 239964 260294 239970
rect 260242 239906 260294 239912
rect 260346 239902 260374 240108
rect 260334 239896 260386 239902
rect 260438 239873 260466 240108
rect 260334 239838 260386 239844
rect 260424 239864 260480 239873
rect 260530 239850 260558 240108
rect 260622 239970 260650 240108
rect 260610 239964 260662 239970
rect 260610 239906 260662 239912
rect 260714 239850 260742 240108
rect 260806 239970 260834 240108
rect 260794 239964 260846 239970
rect 260794 239906 260846 239912
rect 260898 239902 260926 240108
rect 260990 239902 261018 240108
rect 261082 239970 261110 240108
rect 261174 239970 261202 240108
rect 261266 239970 261294 240108
rect 261358 239970 261386 240108
rect 261450 239970 261478 240108
rect 261070 239964 261122 239970
rect 261070 239906 261122 239912
rect 261162 239964 261214 239970
rect 261162 239906 261214 239912
rect 261254 239964 261306 239970
rect 261254 239906 261306 239912
rect 261346 239964 261398 239970
rect 261346 239906 261398 239912
rect 261438 239964 261490 239970
rect 261438 239906 261490 239912
rect 260886 239896 260938 239902
rect 260530 239822 260604 239850
rect 260714 239822 260788 239850
rect 260886 239838 260938 239844
rect 260978 239896 261030 239902
rect 260978 239838 261030 239844
rect 260424 239799 260480 239808
rect 260162 239686 260236 239714
rect 259736 239634 259788 239640
rect 260024 239652 260098 239680
rect 259642 237144 259698 237153
rect 259642 237079 259698 237088
rect 259748 230474 259776 239634
rect 259828 239624 259880 239630
rect 259828 239566 259880 239572
rect 259840 237046 259868 239566
rect 259920 239556 259972 239562
rect 259920 239498 259972 239504
rect 259828 237040 259880 237046
rect 259828 236982 259880 236988
rect 259656 230446 259776 230474
rect 259656 222086 259684 230446
rect 259932 224670 259960 239498
rect 260024 234297 260052 239652
rect 260102 239592 260158 239601
rect 260102 239527 260104 239536
rect 260156 239527 260158 239536
rect 260104 239498 260156 239504
rect 260208 239034 260236 239686
rect 260288 239692 260340 239698
rect 260288 239634 260340 239640
rect 260116 239006 260236 239034
rect 260116 234433 260144 239006
rect 260300 238814 260328 239634
rect 260380 239624 260432 239630
rect 260576 239578 260604 239822
rect 260656 239760 260708 239766
rect 260656 239702 260708 239708
rect 260380 239566 260432 239572
rect 260288 238808 260340 238814
rect 260288 238750 260340 238756
rect 260392 237561 260420 239566
rect 260484 239550 260604 239578
rect 260484 239329 260512 239550
rect 260564 239488 260616 239494
rect 260564 239430 260616 239436
rect 260470 239320 260526 239329
rect 260470 239255 260526 239264
rect 260472 239080 260524 239086
rect 260472 239022 260524 239028
rect 260484 238882 260512 239022
rect 260472 238876 260524 238882
rect 260472 238818 260524 238824
rect 260472 238128 260524 238134
rect 260472 238070 260524 238076
rect 260378 237552 260434 237561
rect 260378 237487 260434 237496
rect 260380 237244 260432 237250
rect 260380 237186 260432 237192
rect 260392 236994 260420 237186
rect 260300 236966 260420 236994
rect 260196 234932 260248 234938
rect 260196 234874 260248 234880
rect 260102 234424 260158 234433
rect 260102 234359 260158 234368
rect 260010 234288 260066 234297
rect 260010 234223 260066 234232
rect 260208 226302 260236 234874
rect 260196 226296 260248 226302
rect 260196 226238 260248 226244
rect 259920 224664 259972 224670
rect 259920 224606 259972 224612
rect 259644 222080 259696 222086
rect 259644 222022 259696 222028
rect 259552 210996 259604 211002
rect 259552 210938 259604 210944
rect 260102 200696 260158 200705
rect 260102 200631 260158 200640
rect 259368 6180 259420 6186
rect 259368 6122 259420 6128
rect 259368 3800 259420 3806
rect 259368 3742 259420 3748
rect 259380 3398 259408 3742
rect 259840 3738 260052 3754
rect 259828 3732 260064 3738
rect 259880 3726 260012 3732
rect 259828 3674 259880 3680
rect 260012 3674 260064 3680
rect 260116 3670 260144 200631
rect 260300 6914 260328 236966
rect 260484 234614 260512 238070
rect 260576 237930 260604 239430
rect 260564 237924 260616 237930
rect 260564 237866 260616 237872
rect 260392 234586 260512 234614
rect 260392 225622 260420 234586
rect 260668 231849 260696 239702
rect 260760 237250 260788 239822
rect 261116 239828 261168 239834
rect 261116 239770 261168 239776
rect 260840 239760 260892 239766
rect 260840 239702 260892 239708
rect 261024 239760 261076 239766
rect 261024 239702 261076 239708
rect 260852 238678 260880 239702
rect 260932 239692 260984 239698
rect 260932 239634 260984 239640
rect 260944 239601 260972 239634
rect 260930 239592 260986 239601
rect 260930 239527 260986 239536
rect 260840 238672 260892 238678
rect 260840 238614 260892 238620
rect 260748 237244 260800 237250
rect 260748 237186 260800 237192
rect 260748 236156 260800 236162
rect 260748 236098 260800 236104
rect 260654 231840 260710 231849
rect 260654 231775 260710 231784
rect 260760 230874 260788 236098
rect 261036 231713 261064 239702
rect 261022 231704 261078 231713
rect 261022 231639 261078 231648
rect 260668 230846 260788 230874
rect 260668 227118 260696 230846
rect 261128 230474 261156 239770
rect 261346 239760 261398 239766
rect 261036 230446 261156 230474
rect 261220 239720 261346 239748
rect 260840 229492 260892 229498
rect 260840 229434 260892 229440
rect 260746 228984 260802 228993
rect 260746 228919 260802 228928
rect 260656 227112 260708 227118
rect 260656 227054 260708 227060
rect 260380 225616 260432 225622
rect 260380 225558 260432 225564
rect 260760 219162 260788 228919
rect 260852 219434 260880 229434
rect 260932 229424 260984 229430
rect 260932 229366 260984 229372
rect 260944 224806 260972 229366
rect 260932 224800 260984 224806
rect 260932 224742 260984 224748
rect 261036 224738 261064 230446
rect 261220 226098 261248 239720
rect 261542 239748 261570 240108
rect 261634 239970 261662 240108
rect 261726 239970 261754 240108
rect 261622 239964 261674 239970
rect 261622 239906 261674 239912
rect 261714 239964 261766 239970
rect 261714 239906 261766 239912
rect 261818 239902 261846 240108
rect 261910 239907 261938 240108
rect 262002 239970 262030 240108
rect 261990 239964 262042 239970
rect 261806 239896 261858 239902
rect 261806 239838 261858 239844
rect 261896 239898 261952 239907
rect 261990 239906 262042 239912
rect 262094 239907 262122 240108
rect 261896 239833 261952 239842
rect 262080 239898 262136 239907
rect 262080 239833 262136 239842
rect 261346 239702 261398 239708
rect 261496 239720 261570 239748
rect 261392 239556 261444 239562
rect 261392 239498 261444 239504
rect 261404 229498 261432 239498
rect 261496 237794 261524 239720
rect 261852 239692 261904 239698
rect 261852 239634 261904 239640
rect 261944 239692 261996 239698
rect 261944 239634 261996 239640
rect 261576 239556 261628 239562
rect 261576 239498 261628 239504
rect 261484 237788 261536 237794
rect 261484 237730 261536 237736
rect 261392 229492 261444 229498
rect 261392 229434 261444 229440
rect 261588 229430 261616 239498
rect 261666 239320 261722 239329
rect 261666 239255 261722 239264
rect 261680 238542 261708 239255
rect 261864 239154 261892 239634
rect 261852 239148 261904 239154
rect 261852 239090 261904 239096
rect 261668 238536 261720 238542
rect 261668 238478 261720 238484
rect 261850 236736 261906 236745
rect 261850 236671 261906 236680
rect 261668 236496 261720 236502
rect 261668 236438 261720 236444
rect 261576 229424 261628 229430
rect 261576 229366 261628 229372
rect 261208 226092 261260 226098
rect 261208 226034 261260 226040
rect 261680 225350 261708 236438
rect 261864 226137 261892 236671
rect 261956 233073 261984 239634
rect 262186 239476 262214 240108
rect 262278 239902 262306 240108
rect 262370 239970 262398 240108
rect 262358 239964 262410 239970
rect 262358 239906 262410 239912
rect 262266 239896 262318 239902
rect 262266 239838 262318 239844
rect 262462 239850 262490 240108
rect 262554 239970 262582 240108
rect 262646 239970 262674 240108
rect 262542 239964 262594 239970
rect 262542 239906 262594 239912
rect 262634 239964 262686 239970
rect 262634 239906 262686 239912
rect 262586 239864 262642 239873
rect 262462 239822 262536 239850
rect 262404 239760 262456 239766
rect 262508 239737 262536 239822
rect 262738 239816 262766 240108
rect 262586 239799 262588 239808
rect 262640 239799 262642 239808
rect 262588 239770 262640 239776
rect 262692 239788 262766 239816
rect 262404 239702 262456 239708
rect 262494 239728 262550 239737
rect 262312 239692 262364 239698
rect 262312 239634 262364 239640
rect 262140 239448 262214 239476
rect 261942 233064 261998 233073
rect 261942 232999 261998 233008
rect 262140 227497 262168 239448
rect 262220 235204 262272 235210
rect 262220 235146 262272 235152
rect 262126 227488 262182 227497
rect 262126 227423 262182 227432
rect 261850 226128 261906 226137
rect 261850 226063 261906 226072
rect 261668 225344 261720 225350
rect 261668 225286 261720 225292
rect 261024 224732 261076 224738
rect 261024 224674 261076 224680
rect 260840 219428 260892 219434
rect 260840 219370 260892 219376
rect 260748 219156 260800 219162
rect 260748 219098 260800 219104
rect 260760 145586 260788 219098
rect 262232 212498 262260 235146
rect 262324 234938 262352 239634
rect 262312 234932 262364 234938
rect 262312 234874 262364 234880
rect 262416 232801 262444 239702
rect 262692 239714 262720 239788
rect 262494 239663 262550 239672
rect 262600 239686 262720 239714
rect 262830 239714 262858 240108
rect 262922 239902 262950 240108
rect 263014 239907 263042 240108
rect 263106 239970 263134 240108
rect 263198 239970 263226 240108
rect 263094 239964 263146 239970
rect 262910 239896 262962 239902
rect 262910 239838 262962 239844
rect 263000 239898 263056 239907
rect 263094 239906 263146 239912
rect 263186 239964 263238 239970
rect 263186 239906 263238 239912
rect 263290 239850 263318 240108
rect 263000 239833 263056 239842
rect 263244 239834 263318 239850
rect 263140 239828 263192 239834
rect 263140 239770 263192 239776
rect 263232 239828 263318 239834
rect 263284 239822 263318 239828
rect 263232 239770 263284 239776
rect 262954 239728 263010 239737
rect 262830 239686 262904 239714
rect 262496 239624 262548 239630
rect 262496 239566 262548 239572
rect 262508 234025 262536 239566
rect 262600 235249 262628 239686
rect 262680 239624 262732 239630
rect 262680 239566 262732 239572
rect 262586 235240 262642 235249
rect 262586 235175 262642 235184
rect 262692 234161 262720 239566
rect 262772 239556 262824 239562
rect 262772 239498 262824 239504
rect 262678 234152 262734 234161
rect 262678 234087 262734 234096
rect 262494 234016 262550 234025
rect 262494 233951 262550 233960
rect 262402 232792 262458 232801
rect 262402 232727 262458 232736
rect 262784 231441 262812 239498
rect 262876 235210 262904 239686
rect 262954 239663 263010 239672
rect 262968 238134 262996 239663
rect 262956 238128 263008 238134
rect 262956 238070 263008 238076
rect 263152 236688 263180 239770
rect 263382 239714 263410 240108
rect 263474 239970 263502 240108
rect 263462 239964 263514 239970
rect 263462 239906 263514 239912
rect 263566 239902 263594 240108
rect 263554 239896 263606 239902
rect 263554 239838 263606 239844
rect 263060 236660 263180 236688
rect 263244 239686 263410 239714
rect 263506 239728 263562 239737
rect 262956 235340 263008 235346
rect 262956 235282 263008 235288
rect 262968 235210 262996 235282
rect 262864 235204 262916 235210
rect 262864 235146 262916 235152
rect 262956 235204 263008 235210
rect 262956 235146 263008 235152
rect 262770 231432 262826 231441
rect 262770 231367 262826 231376
rect 263060 228993 263088 236660
rect 263140 235884 263192 235890
rect 263140 235826 263192 235832
rect 263046 228984 263102 228993
rect 263046 228919 263102 228928
rect 263152 224466 263180 235826
rect 263244 225729 263272 239686
rect 263506 239663 263508 239672
rect 263560 239663 263562 239672
rect 263658 239680 263686 240108
rect 263750 239748 263778 240108
rect 263842 239873 263870 240108
rect 263934 239970 263962 240108
rect 263922 239964 263974 239970
rect 263922 239906 263974 239912
rect 263828 239864 263884 239873
rect 264026 239850 264054 240108
rect 264118 239970 264146 240108
rect 264210 239970 264238 240108
rect 264302 239970 264330 240108
rect 264106 239964 264158 239970
rect 264106 239906 264158 239912
rect 264198 239964 264250 239970
rect 264198 239906 264250 239912
rect 264290 239964 264342 239970
rect 264290 239906 264342 239912
rect 264394 239850 264422 240108
rect 264486 239873 264514 240108
rect 264026 239822 264284 239850
rect 263828 239799 263884 239808
rect 263968 239760 264020 239766
rect 263750 239720 263824 239748
rect 263658 239652 263732 239680
rect 263508 239634 263560 239640
rect 263324 239556 263376 239562
rect 263324 239498 263376 239504
rect 263230 225720 263286 225729
rect 263230 225655 263286 225664
rect 263140 224460 263192 224466
rect 263140 224402 263192 224408
rect 262220 212492 262272 212498
rect 262220 212434 262272 212440
rect 263336 186998 263364 239498
rect 263508 239420 263560 239426
rect 263508 239362 263560 239368
rect 263520 238746 263548 239362
rect 263598 239184 263654 239193
rect 263598 239119 263654 239128
rect 263508 238740 263560 238746
rect 263508 238682 263560 238688
rect 263416 234932 263468 234938
rect 263416 234874 263468 234880
rect 263428 230217 263456 234874
rect 263612 233234 263640 239119
rect 263704 237300 263732 239652
rect 263796 239329 263824 239720
rect 263968 239702 264020 239708
rect 264060 239760 264112 239766
rect 264060 239702 264112 239708
rect 264152 239760 264204 239766
rect 264152 239702 264204 239708
rect 263876 239624 263928 239630
rect 263876 239566 263928 239572
rect 263782 239320 263838 239329
rect 263782 239255 263838 239264
rect 263888 239193 263916 239566
rect 263874 239184 263930 239193
rect 263874 239119 263930 239128
rect 263874 237688 263930 237697
rect 263874 237623 263930 237632
rect 263888 237425 263916 237623
rect 263874 237416 263930 237425
rect 263874 237351 263930 237360
rect 263704 237272 263916 237300
rect 263784 236020 263836 236026
rect 263784 235962 263836 235968
rect 263520 233206 263640 233234
rect 263414 230208 263470 230217
rect 263414 230143 263470 230152
rect 263324 186992 263376 186998
rect 263324 186934 263376 186940
rect 260748 145580 260800 145586
rect 260748 145522 260800 145528
rect 263428 144226 263456 230143
rect 263416 144220 263468 144226
rect 263416 144162 263468 144168
rect 263520 141438 263548 233206
rect 263796 230353 263824 235962
rect 263888 235521 263916 237272
rect 263874 235512 263930 235521
rect 263874 235447 263930 235456
rect 263888 231854 263916 235447
rect 263980 234569 264008 239702
rect 264072 237969 264100 239702
rect 264058 237960 264114 237969
rect 264058 237895 264114 237904
rect 264164 236026 264192 239702
rect 264256 239601 264284 239822
rect 264348 239822 264422 239850
rect 264472 239864 264528 239873
rect 264348 239737 264376 239822
rect 264578 239834 264606 240108
rect 264670 239970 264698 240108
rect 264762 239970 264790 240108
rect 264658 239964 264710 239970
rect 264658 239906 264710 239912
rect 264750 239964 264802 239970
rect 264750 239906 264802 239912
rect 264472 239799 264528 239808
rect 264566 239828 264618 239834
rect 264566 239770 264618 239776
rect 264704 239828 264756 239834
rect 264704 239770 264756 239776
rect 264334 239728 264390 239737
rect 264610 239728 264666 239737
rect 264390 239686 264468 239714
rect 264334 239663 264390 239672
rect 264242 239592 264298 239601
rect 264242 239527 264298 239536
rect 264244 238604 264296 238610
rect 264244 238546 264296 238552
rect 264152 236020 264204 236026
rect 264152 235962 264204 235968
rect 263966 234560 264022 234569
rect 263966 234495 264022 234504
rect 263888 231826 264100 231854
rect 264072 230790 264100 231826
rect 264060 230784 264112 230790
rect 264060 230726 264112 230732
rect 263782 230344 263838 230353
rect 263782 230279 263838 230288
rect 264256 224954 264284 238546
rect 264334 236600 264390 236609
rect 264334 236535 264390 236544
rect 264348 225554 264376 236535
rect 264440 229634 264468 239686
rect 264532 239686 264610 239714
rect 264532 238610 264560 239686
rect 264610 239663 264666 239672
rect 264520 238604 264572 238610
rect 264520 238546 264572 238552
rect 264518 238504 264574 238513
rect 264518 238439 264574 238448
rect 264428 229628 264480 229634
rect 264428 229570 264480 229576
rect 264336 225548 264388 225554
rect 264336 225490 264388 225496
rect 263704 224926 264284 224954
rect 263704 224874 263732 224926
rect 263692 224868 263744 224874
rect 263692 224810 263744 224816
rect 264532 209098 264560 238439
rect 264716 231854 264744 239770
rect 264854 239748 264882 240108
rect 264946 239907 264974 240108
rect 265038 239970 265066 240108
rect 265130 239970 265158 240108
rect 265026 239964 265078 239970
rect 264932 239898 264988 239907
rect 265026 239906 265078 239912
rect 265118 239964 265170 239970
rect 265118 239906 265170 239912
rect 265222 239850 265250 240108
rect 265314 239970 265342 240108
rect 265406 239970 265434 240108
rect 265302 239964 265354 239970
rect 265302 239906 265354 239912
rect 265394 239964 265446 239970
rect 265394 239906 265446 239912
rect 265498 239850 265526 240108
rect 264932 239833 264988 239842
rect 265072 239828 265124 239834
rect 265072 239770 265124 239776
rect 265176 239822 265250 239850
rect 265452 239822 265526 239850
rect 264980 239760 265032 239766
rect 264854 239720 264928 239748
rect 264796 239624 264848 239630
rect 264796 239566 264848 239572
rect 264624 231826 264744 231854
rect 264624 223378 264652 231826
rect 264704 229628 264756 229634
rect 264704 229570 264756 229576
rect 264612 223372 264664 223378
rect 264612 223314 264664 223320
rect 264612 221468 264664 221474
rect 264612 221410 264664 221416
rect 264624 221241 264652 221410
rect 264610 221232 264666 221241
rect 264610 221167 264666 221176
rect 264520 209092 264572 209098
rect 264520 209034 264572 209040
rect 264624 185638 264652 221167
rect 264612 185632 264664 185638
rect 264612 185574 264664 185580
rect 264716 184210 264744 229570
rect 264704 184204 264756 184210
rect 264704 184146 264756 184152
rect 264808 181490 264836 239566
rect 264900 238513 264928 239720
rect 264978 239728 264980 239737
rect 265032 239728 265034 239737
rect 264978 239663 265034 239672
rect 264980 239556 265032 239562
rect 264980 239498 265032 239504
rect 264886 238504 264942 238513
rect 264886 238439 264942 238448
rect 264888 238128 264940 238134
rect 264888 238070 264940 238076
rect 264900 231577 264928 238070
rect 264992 236745 265020 239498
rect 265084 237386 265112 239770
rect 265072 237380 265124 237386
rect 265072 237322 265124 237328
rect 264978 236736 265034 236745
rect 264978 236671 265034 236680
rect 264886 231568 264942 231577
rect 264886 231503 264942 231512
rect 264888 230784 264940 230790
rect 264888 230726 264940 230732
rect 264796 181484 264848 181490
rect 264796 181426 264848 181432
rect 263508 141432 263560 141438
rect 262218 141400 262274 141409
rect 263508 141374 263560 141380
rect 262218 141335 262274 141344
rect 262232 16574 262260 141335
rect 264900 29646 264928 230726
rect 265176 224954 265204 239822
rect 265256 239760 265308 239766
rect 265256 239702 265308 239708
rect 265346 239728 265402 239737
rect 265268 238048 265296 239702
rect 265346 239663 265348 239672
rect 265400 239663 265402 239672
rect 265348 239634 265400 239640
rect 265348 239556 265400 239562
rect 265348 239498 265400 239504
rect 265360 239358 265388 239498
rect 265348 239352 265400 239358
rect 265348 239294 265400 239300
rect 265452 238116 265480 239822
rect 265590 239748 265618 240108
rect 265682 239970 265710 240108
rect 265774 239970 265802 240108
rect 265670 239964 265722 239970
rect 265670 239906 265722 239912
rect 265762 239964 265814 239970
rect 265762 239906 265814 239912
rect 265866 239850 265894 240108
rect 265958 239873 265986 240108
rect 265716 239828 265768 239834
rect 265716 239770 265768 239776
rect 265820 239822 265894 239850
rect 265944 239864 266000 239873
rect 265590 239720 265664 239748
rect 265452 238088 265572 238116
rect 265268 238020 265480 238048
rect 265256 236632 265308 236638
rect 265256 236574 265308 236580
rect 265268 231402 265296 236574
rect 265452 235890 265480 238020
rect 265440 235884 265492 235890
rect 265440 235826 265492 235832
rect 265256 231396 265308 231402
rect 265256 231338 265308 231344
rect 265544 229634 265572 238088
rect 265636 237318 265664 239720
rect 265728 237969 265756 239770
rect 265714 237960 265770 237969
rect 265714 237895 265770 237904
rect 265624 237312 265676 237318
rect 265624 237254 265676 237260
rect 265820 231854 265848 239822
rect 266050 239850 266078 240108
rect 266142 239970 266170 240108
rect 266234 239970 266262 240108
rect 266130 239964 266182 239970
rect 266130 239906 266182 239912
rect 266222 239964 266274 239970
rect 266222 239906 266274 239912
rect 266326 239902 266354 240108
rect 266418 239970 266446 240108
rect 266510 239970 266538 240108
rect 266406 239964 266458 239970
rect 266406 239906 266458 239912
rect 266498 239964 266550 239970
rect 266498 239906 266550 239912
rect 266314 239896 266366 239902
rect 266050 239822 266124 239850
rect 266602 239873 266630 240108
rect 266314 239838 266366 239844
rect 266588 239864 266644 239873
rect 265944 239799 266000 239808
rect 266096 239737 266124 239822
rect 266588 239799 266644 239808
rect 266452 239760 266504 239766
rect 266082 239728 266138 239737
rect 266452 239702 266504 239708
rect 266542 239728 266598 239737
rect 266082 239663 266138 239672
rect 266084 239624 266136 239630
rect 266084 239566 266136 239572
rect 266360 239624 266412 239630
rect 266360 239566 266412 239572
rect 266096 236178 266124 239566
rect 266268 239420 266320 239426
rect 266268 239362 266320 239368
rect 266280 238746 266308 239362
rect 266268 238740 266320 238746
rect 266268 238682 266320 238688
rect 266096 236150 266308 236178
rect 266176 236088 266228 236094
rect 266176 236030 266228 236036
rect 266084 232280 266136 232286
rect 266084 232222 266136 232228
rect 265636 231826 265848 231854
rect 265532 229628 265584 229634
rect 265532 229570 265584 229576
rect 265636 228857 265664 231826
rect 265714 231024 265770 231033
rect 265714 230959 265770 230968
rect 265622 228848 265678 228857
rect 265622 228783 265678 228792
rect 264992 224926 265204 224954
rect 264992 215150 265020 224926
rect 264980 215144 265032 215150
rect 264980 215086 265032 215092
rect 265728 180130 265756 230959
rect 265992 229628 266044 229634
rect 265992 229570 266044 229576
rect 266004 205562 266032 229570
rect 266096 224954 266124 232222
rect 266188 229786 266216 236030
rect 266280 232393 266308 236150
rect 266372 235278 266400 239566
rect 266464 236858 266492 239702
rect 266694 239714 266722 240108
rect 266786 239902 266814 240108
rect 266878 239970 266906 240108
rect 266866 239964 266918 239970
rect 266866 239906 266918 239912
rect 266774 239896 266826 239902
rect 266970 239850 266998 240108
rect 267062 239970 267090 240108
rect 267154 239970 267182 240108
rect 267050 239964 267102 239970
rect 267050 239906 267102 239912
rect 267142 239964 267194 239970
rect 267142 239906 267194 239912
rect 266774 239838 266826 239844
rect 266924 239822 266998 239850
rect 267094 239864 267150 239873
rect 266820 239760 266872 239766
rect 266818 239728 266820 239737
rect 266872 239728 266874 239737
rect 266694 239686 266768 239714
rect 266542 239663 266598 239672
rect 266556 239358 266584 239663
rect 266636 239624 266688 239630
rect 266636 239566 266688 239572
rect 266544 239352 266596 239358
rect 266544 239294 266596 239300
rect 266648 238105 266676 239566
rect 266634 238096 266690 238105
rect 266634 238031 266690 238040
rect 266464 236830 266584 236858
rect 266452 236700 266504 236706
rect 266452 236642 266504 236648
rect 266360 235272 266412 235278
rect 266360 235214 266412 235220
rect 266266 232384 266322 232393
rect 266266 232319 266322 232328
rect 266188 229758 266308 229786
rect 266096 224926 266216 224954
rect 265992 205556 266044 205562
rect 265992 205498 266044 205504
rect 265716 180124 265768 180130
rect 265716 180066 265768 180072
rect 266188 177342 266216 224926
rect 266176 177336 266228 177342
rect 266176 177278 266228 177284
rect 266280 137290 266308 229758
rect 266464 216578 266492 236642
rect 266556 226953 266584 236830
rect 266542 226944 266598 226953
rect 266542 226879 266598 226888
rect 266740 224954 266768 239686
rect 266818 239663 266874 239672
rect 266820 235272 266872 235278
rect 266820 235214 266872 235220
rect 266832 232529 266860 235214
rect 266818 232520 266874 232529
rect 266818 232455 266874 232464
rect 266924 229094 266952 239822
rect 267246 239816 267274 240108
rect 267338 239952 267366 240108
rect 267398 240094 267780 240122
rect 267556 240032 267608 240038
rect 267554 240000 267556 240009
rect 267608 240000 267610 240009
rect 267464 239964 267516 239970
rect 267338 239924 267464 239952
rect 267554 239935 267610 239944
rect 267464 239906 267516 239912
rect 267646 239864 267702 239873
rect 267094 239799 267150 239808
rect 267004 239760 267056 239766
rect 267108 239748 267136 239799
rect 267056 239720 267136 239748
rect 267200 239788 267274 239816
rect 267556 239828 267608 239834
rect 267004 239702 267056 239708
rect 267200 236706 267228 239788
rect 267646 239799 267702 239808
rect 267556 239770 267608 239776
rect 267372 239556 267424 239562
rect 267372 239498 267424 239504
rect 267384 239358 267412 239498
rect 267372 239352 267424 239358
rect 267372 239294 267424 239300
rect 267280 238740 267332 238746
rect 267280 238682 267332 238688
rect 267188 236700 267240 236706
rect 267188 236642 267240 236648
rect 266556 224926 266768 224954
rect 266832 229066 266952 229094
rect 266556 220658 266584 224926
rect 266544 220652 266596 220658
rect 266544 220594 266596 220600
rect 266832 217938 266860 229066
rect 266820 217932 266872 217938
rect 266820 217874 266872 217880
rect 266452 216572 266504 216578
rect 266452 216514 266504 216520
rect 266360 215960 266412 215966
rect 266360 215902 266412 215908
rect 266268 137284 266320 137290
rect 266268 137226 266320 137232
rect 264888 29640 264940 29646
rect 264888 29582 264940 29588
rect 266372 16574 266400 215902
rect 267292 173194 267320 238682
rect 267384 175982 267412 239294
rect 267568 238950 267596 239770
rect 267660 239766 267688 239799
rect 267648 239760 267700 239766
rect 267648 239702 267700 239708
rect 267556 238944 267608 238950
rect 267556 238886 267608 238892
rect 267554 238368 267610 238377
rect 267554 238303 267610 238312
rect 267372 175976 267424 175982
rect 267372 175918 267424 175924
rect 267568 174554 267596 238303
rect 267556 174548 267608 174554
rect 267556 174490 267608 174496
rect 267280 173188 267332 173194
rect 267280 173130 267332 173136
rect 267660 170406 267688 239702
rect 267752 238746 267780 240094
rect 267844 239970 267872 243471
rect 267936 240106 267964 246191
rect 268108 241324 268160 241330
rect 268108 241266 268160 241272
rect 268014 241088 268070 241097
rect 268014 241023 268070 241032
rect 268028 240242 268056 241023
rect 268120 240922 268148 241266
rect 268200 241256 268252 241262
rect 268200 241198 268252 241204
rect 268108 240916 268160 240922
rect 268108 240858 268160 240864
rect 268016 240236 268068 240242
rect 268016 240178 268068 240184
rect 267924 240100 267976 240106
rect 267924 240042 267976 240048
rect 267832 239964 267884 239970
rect 267832 239906 267884 239912
rect 268212 239562 268240 241198
rect 268292 240576 268344 240582
rect 268292 240518 268344 240524
rect 268304 240174 268332 240518
rect 268292 240168 268344 240174
rect 268292 240110 268344 240116
rect 268200 239556 268252 239562
rect 268200 239498 268252 239504
rect 268200 239352 268252 239358
rect 268200 239294 268252 239300
rect 267924 238944 267976 238950
rect 267924 238886 267976 238892
rect 267936 238814 267964 238886
rect 268212 238882 268240 239294
rect 268200 238876 268252 238882
rect 268200 238818 268252 238824
rect 267924 238808 267976 238814
rect 267924 238750 267976 238756
rect 267740 238740 267792 238746
rect 267740 238682 267792 238688
rect 267832 238060 267884 238066
rect 267832 238002 267884 238008
rect 267740 237448 267792 237454
rect 267740 237390 267792 237396
rect 267752 235822 267780 237390
rect 267740 235816 267792 235822
rect 267740 235758 267792 235764
rect 267844 235210 267872 238002
rect 267832 235204 267884 235210
rect 267832 235146 267884 235152
rect 267648 170400 267700 170406
rect 267648 170342 267700 170348
rect 267844 16574 267872 235146
rect 268396 232422 268424 315522
rect 268474 314664 268530 314673
rect 268474 314599 268530 314608
rect 268488 233753 268516 314599
rect 268568 313336 268620 313342
rect 268568 313278 268620 313284
rect 268580 237017 268608 313278
rect 268660 305652 268712 305658
rect 268660 305594 268712 305600
rect 268672 240145 268700 305594
rect 269672 260160 269724 260166
rect 269672 260102 269724 260108
rect 269580 251864 269632 251870
rect 269580 251806 269632 251812
rect 269302 247616 269358 247625
rect 269302 247551 269358 247560
rect 269120 246356 269172 246362
rect 269120 246298 269172 246304
rect 268936 244996 268988 245002
rect 268936 244938 268988 244944
rect 268842 243672 268898 243681
rect 268842 243607 268898 243616
rect 268750 240816 268806 240825
rect 268750 240751 268806 240760
rect 268764 240446 268792 240751
rect 268752 240440 268804 240446
rect 268752 240382 268804 240388
rect 268856 240281 268884 243607
rect 268842 240272 268898 240281
rect 268842 240207 268898 240216
rect 268658 240136 268714 240145
rect 268658 240071 268714 240080
rect 268948 238649 268976 244938
rect 269028 243568 269080 243574
rect 269028 243510 269080 243516
rect 269040 240106 269068 243510
rect 269132 242321 269160 246298
rect 269212 244928 269264 244934
rect 269212 244870 269264 244876
rect 269118 242312 269174 242321
rect 269118 242247 269174 242256
rect 269118 241224 269174 241233
rect 269118 241159 269174 241168
rect 269028 240100 269080 240106
rect 269028 240042 269080 240048
rect 268934 238640 268990 238649
rect 268934 238575 268990 238584
rect 268660 238060 268712 238066
rect 268660 238002 268712 238008
rect 268672 237289 268700 238002
rect 268658 237280 268714 237289
rect 268658 237215 268714 237224
rect 268566 237008 268622 237017
rect 268566 236943 268622 236952
rect 269040 236094 269068 240042
rect 269132 239601 269160 241159
rect 269224 240310 269252 244870
rect 269316 240378 269344 247551
rect 269486 243808 269542 243817
rect 269486 243743 269542 243752
rect 269500 242894 269528 243743
rect 269408 242866 269528 242894
rect 269304 240372 269356 240378
rect 269304 240314 269356 240320
rect 269212 240304 269264 240310
rect 269212 240246 269264 240252
rect 269408 239698 269436 242866
rect 269396 239692 269448 239698
rect 269396 239634 269448 239640
rect 269118 239592 269174 239601
rect 269118 239527 269174 239536
rect 269120 237788 269172 237794
rect 269120 237730 269172 237736
rect 269028 236088 269080 236094
rect 269028 236030 269080 236036
rect 269132 235657 269160 237730
rect 269118 235648 269174 235657
rect 269118 235583 269174 235592
rect 268474 233744 268530 233753
rect 268474 233679 268530 233688
rect 268384 232416 268436 232422
rect 268384 232358 268436 232364
rect 269408 232286 269436 239634
rect 269488 239556 269540 239562
rect 269488 239498 269540 239504
rect 269500 238241 269528 239498
rect 269486 238232 269542 238241
rect 269592 238202 269620 251806
rect 269684 238270 269712 260102
rect 269672 238264 269724 238270
rect 269672 238206 269724 238212
rect 269486 238167 269542 238176
rect 269580 238196 269632 238202
rect 269580 238138 269632 238144
rect 269776 236434 269804 319602
rect 271142 317248 271198 317257
rect 271142 317183 271198 317192
rect 269856 314560 269908 314566
rect 269856 314502 269908 314508
rect 269764 236428 269816 236434
rect 269764 236370 269816 236376
rect 269396 232280 269448 232286
rect 269396 232222 269448 232228
rect 269118 228304 269174 228313
rect 269118 228239 269174 228248
rect 269132 16574 269160 228239
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 267844 16546 268424 16574
rect 269132 16546 269712 16574
rect 260208 6886 260328 6914
rect 260104 3664 260156 3670
rect 260104 3606 260156 3612
rect 260208 3482 260236 6886
rect 260656 4072 260708 4078
rect 260656 4014 260708 4020
rect 259472 3454 260236 3482
rect 259368 3392 259420 3398
rect 259368 3334 259420 3340
rect 259472 480 259500 3454
rect 260668 480 260696 4014
rect 261760 3664 261812 3670
rect 261760 3606 261812 3612
rect 261772 480 261800 3606
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 265348 3800 265400 3806
rect 265348 3742 265400 3748
rect 264152 3392 264204 3398
rect 264152 3334 264204 3340
rect 264164 480 264192 3334
rect 265360 480 265388 3742
rect 266556 480 266584 16546
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 267752 480 267780 3470
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 269684 3482 269712 16546
rect 269776 3670 269804 236370
rect 269868 228274 269896 314502
rect 270040 314288 270092 314294
rect 270040 314230 270092 314236
rect 269948 290080 270000 290086
rect 269948 290022 270000 290028
rect 269856 228268 269908 228274
rect 269856 228210 269908 228216
rect 269960 206990 269988 290022
rect 270052 237153 270080 314230
rect 270130 286512 270186 286521
rect 270130 286447 270186 286456
rect 270144 237930 270172 286447
rect 270224 284980 270276 284986
rect 270224 284922 270276 284928
rect 270236 238406 270264 284922
rect 271052 282192 271104 282198
rect 271052 282134 271104 282140
rect 270316 275324 270368 275330
rect 270316 275266 270368 275272
rect 270328 238474 270356 275266
rect 270960 273964 271012 273970
rect 270960 273906 271012 273912
rect 270408 264240 270460 264246
rect 270408 264182 270460 264188
rect 270316 238468 270368 238474
rect 270316 238410 270368 238416
rect 270224 238400 270276 238406
rect 270224 238342 270276 238348
rect 270420 238338 270448 264182
rect 270408 238332 270460 238338
rect 270408 238274 270460 238280
rect 270132 237924 270184 237930
rect 270132 237866 270184 237872
rect 270972 237561 271000 273906
rect 271064 237726 271092 282134
rect 271156 239737 271184 317183
rect 271420 317144 271472 317150
rect 271420 317086 271472 317092
rect 271328 316464 271380 316470
rect 271328 316406 271380 316412
rect 271236 315648 271288 315654
rect 271236 315590 271288 315596
rect 271142 239728 271198 239737
rect 271142 239663 271198 239672
rect 271052 237720 271104 237726
rect 271052 237662 271104 237668
rect 270958 237552 271014 237561
rect 270958 237487 271014 237496
rect 270038 237144 270094 237153
rect 270038 237079 270094 237088
rect 271144 236700 271196 236706
rect 271144 236642 271196 236648
rect 269948 206984 270000 206990
rect 269948 206926 270000 206932
rect 269764 3664 269816 3670
rect 269764 3606 269816 3612
rect 271156 3602 271184 236642
rect 271248 233782 271276 315590
rect 271236 233776 271288 233782
rect 271236 233718 271288 233724
rect 270868 3596 270920 3602
rect 270868 3538 270920 3544
rect 271144 3596 271196 3602
rect 271144 3538 271196 3544
rect 269684 3454 270080 3482
rect 270052 480 270080 3454
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270880 354 270908 3538
rect 271248 3534 271276 233718
rect 271340 226982 271368 316406
rect 271432 229498 271460 317086
rect 271512 316940 271564 316946
rect 271512 316882 271564 316888
rect 271524 229809 271552 316882
rect 271602 315888 271658 315897
rect 271602 315823 271658 315832
rect 271616 230926 271644 315823
rect 272524 315512 272576 315518
rect 272524 315454 272576 315460
rect 271696 313132 271748 313138
rect 271696 313074 271748 313080
rect 271708 236706 271736 313074
rect 271788 283620 271840 283626
rect 271788 283562 271840 283568
rect 271800 237697 271828 283562
rect 271786 237688 271842 237697
rect 271786 237623 271842 237632
rect 271696 236700 271748 236706
rect 271696 236642 271748 236648
rect 271880 232620 271932 232626
rect 271880 232562 271932 232568
rect 271892 232218 271920 232562
rect 271880 232212 271932 232218
rect 271880 232154 271932 232160
rect 271604 230920 271656 230926
rect 271604 230862 271656 230868
rect 271510 229800 271566 229809
rect 271510 229735 271566 229744
rect 271420 229492 271472 229498
rect 271420 229434 271472 229440
rect 271328 226976 271380 226982
rect 271328 226918 271380 226924
rect 272536 224097 272564 315454
rect 272628 233714 272656 320486
rect 272984 318980 273036 318986
rect 272984 318922 273036 318928
rect 272892 318572 272944 318578
rect 272892 318514 272944 318520
rect 272800 317484 272852 317490
rect 272800 317426 272852 317432
rect 272708 315784 272760 315790
rect 272708 315726 272760 315732
rect 272616 233708 272668 233714
rect 272616 233650 272668 233656
rect 272720 229430 272748 315726
rect 272812 232762 272840 317426
rect 272800 232756 272852 232762
rect 272800 232698 272852 232704
rect 272904 232354 272932 318514
rect 272996 235142 273024 318922
rect 274180 317348 274232 317354
rect 274180 317290 274232 317296
rect 273996 317076 274048 317082
rect 273996 317018 274048 317024
rect 273168 317008 273220 317014
rect 273168 316950 273220 316956
rect 272984 235136 273036 235142
rect 272984 235078 273036 235084
rect 272892 232348 272944 232354
rect 272892 232290 272944 232296
rect 273180 232218 273208 316950
rect 273902 316840 273958 316849
rect 273902 316775 273958 316784
rect 273916 239465 273944 316775
rect 273902 239456 273958 239465
rect 273902 239391 273958 239400
rect 273168 232212 273220 232218
rect 273168 232154 273220 232160
rect 273904 232212 273956 232218
rect 273904 232154 273956 232160
rect 272708 229424 272760 229430
rect 272708 229366 272760 229372
rect 273260 225480 273312 225486
rect 273260 225422 273312 225428
rect 273272 225010 273300 225422
rect 273260 225004 273312 225010
rect 273260 224946 273312 224952
rect 272522 224088 272578 224097
rect 272522 224023 272578 224032
rect 273168 223032 273220 223038
rect 273168 222974 273220 222980
rect 273180 221610 273208 222974
rect 273168 221604 273220 221610
rect 273168 221546 273220 221552
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 272444 480 272472 3470
rect 273180 3126 273208 221546
rect 273168 3120 273220 3126
rect 273168 3062 273220 3068
rect 271206 354 271318 480
rect 270880 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 224946
rect 273916 3534 273944 232154
rect 274008 225010 274036 317018
rect 274088 315716 274140 315722
rect 274088 315658 274140 315664
rect 274100 226846 274128 315658
rect 274192 229838 274220 317290
rect 274272 317280 274324 317286
rect 274272 317222 274324 317228
rect 274180 229832 274232 229838
rect 274180 229774 274232 229780
rect 274284 229770 274312 317222
rect 274364 315852 274416 315858
rect 274364 315794 274416 315800
rect 274376 230994 274404 315794
rect 274548 314492 274600 314498
rect 274548 314434 274600 314440
rect 274456 302932 274508 302938
rect 274456 302874 274508 302880
rect 274468 239358 274496 302874
rect 274456 239352 274508 239358
rect 274456 239294 274508 239300
rect 274560 233850 274588 314434
rect 275112 304502 275140 375838
rect 278596 374876 278648 374882
rect 278596 374818 278648 374824
rect 277952 374808 278004 374814
rect 277952 374750 278004 374756
rect 275744 374740 275796 374746
rect 275744 374682 275796 374688
rect 275192 374536 275244 374542
rect 275192 374478 275244 374484
rect 275100 304496 275152 304502
rect 275100 304438 275152 304444
rect 275204 300830 275232 374478
rect 275652 320272 275704 320278
rect 275652 320214 275704 320220
rect 275284 319048 275336 319054
rect 275284 318990 275336 318996
rect 275192 300824 275244 300830
rect 275192 300766 275244 300772
rect 275296 235482 275324 318990
rect 275560 315988 275612 315994
rect 275560 315930 275612 315936
rect 275466 315072 275522 315081
rect 275466 315007 275522 315016
rect 275376 312996 275428 313002
rect 275376 312938 275428 312944
rect 275284 235476 275336 235482
rect 275284 235418 275336 235424
rect 274548 233844 274600 233850
rect 274548 233786 274600 233792
rect 275284 233844 275336 233850
rect 275284 233786 275336 233792
rect 274364 230988 274416 230994
rect 274364 230930 274416 230936
rect 274272 229764 274324 229770
rect 274272 229706 274324 229712
rect 274088 226840 274140 226846
rect 274088 226782 274140 226788
rect 273996 225004 274048 225010
rect 273996 224946 274048 224952
rect 274824 3664 274876 3670
rect 274824 3606 274876 3612
rect 273904 3528 273956 3534
rect 273904 3470 273956 3476
rect 274836 480 274864 3606
rect 275296 3602 275324 233786
rect 275388 221377 275416 312938
rect 275480 224330 275508 315007
rect 275572 231062 275600 315930
rect 275664 236910 275692 320214
rect 275756 290494 275784 374682
rect 275928 372700 275980 372706
rect 275928 372642 275980 372648
rect 275836 307556 275888 307562
rect 275836 307498 275888 307504
rect 275744 290488 275796 290494
rect 275744 290430 275796 290436
rect 275652 236904 275704 236910
rect 275652 236846 275704 236852
rect 275560 231056 275612 231062
rect 275560 230998 275612 231004
rect 275848 225418 275876 307498
rect 275940 292058 275968 372642
rect 277860 370116 277912 370122
rect 277860 370058 277912 370064
rect 277584 318640 277636 318646
rect 277582 318608 277584 318617
rect 277636 318608 277638 318617
rect 277582 318543 277638 318552
rect 277766 318200 277822 318209
rect 277766 318135 277822 318144
rect 277780 317801 277808 318135
rect 277766 317792 277822 317801
rect 277766 317727 277822 317736
rect 276940 317688 276992 317694
rect 276940 317630 276992 317636
rect 276848 316600 276900 316606
rect 276848 316542 276900 316548
rect 276756 315920 276808 315926
rect 276756 315862 276808 315868
rect 276664 314628 276716 314634
rect 276664 314570 276716 314576
rect 276020 310344 276072 310350
rect 276020 310286 276072 310292
rect 276032 307358 276060 310286
rect 276020 307352 276072 307358
rect 276020 307294 276072 307300
rect 275928 292052 275980 292058
rect 275928 291994 275980 292000
rect 275928 235272 275980 235278
rect 275928 235214 275980 235220
rect 275836 225412 275888 225418
rect 275836 225354 275888 225360
rect 275468 224324 275520 224330
rect 275468 224266 275520 224272
rect 275374 221368 275430 221377
rect 275374 221303 275430 221312
rect 275940 4078 275968 235214
rect 276676 220153 276704 314570
rect 276768 226914 276796 315862
rect 276860 229906 276888 316542
rect 276952 232694 276980 317630
rect 277308 316872 277360 316878
rect 277308 316814 277360 316820
rect 277216 311568 277268 311574
rect 277216 311510 277268 311516
rect 277228 233918 277256 311510
rect 277216 233912 277268 233918
rect 277216 233854 277268 233860
rect 277320 233209 277348 316814
rect 277872 297430 277900 370058
rect 277860 297424 277912 297430
rect 277860 297366 277912 297372
rect 277964 296070 277992 374750
rect 278504 374672 278556 374678
rect 278504 374614 278556 374620
rect 278044 318844 278096 318850
rect 278044 318786 278096 318792
rect 277952 296064 278004 296070
rect 277952 296006 278004 296012
rect 278056 235521 278084 318786
rect 278412 318640 278464 318646
rect 278410 318608 278412 318617
rect 278464 318608 278466 318617
rect 278410 318543 278466 318552
rect 278410 318472 278466 318481
rect 278410 318407 278466 318416
rect 278424 318073 278452 318407
rect 278410 318064 278466 318073
rect 278410 317999 278466 318008
rect 278136 317960 278188 317966
rect 278136 317902 278188 317908
rect 278148 236298 278176 317902
rect 278318 317384 278374 317393
rect 278318 317319 278374 317328
rect 278228 310276 278280 310282
rect 278228 310218 278280 310224
rect 278136 236292 278188 236298
rect 278136 236234 278188 236240
rect 278042 235512 278098 235521
rect 278042 235447 278098 235456
rect 278044 233912 278096 233918
rect 278044 233854 278096 233860
rect 277306 233200 277362 233209
rect 277306 233135 277362 233144
rect 276940 232688 276992 232694
rect 276940 232630 276992 232636
rect 276848 229900 276900 229906
rect 276848 229842 276900 229848
rect 276756 226908 276808 226914
rect 276756 226850 276808 226856
rect 276662 220144 276718 220153
rect 276662 220079 276718 220088
rect 275928 4072 275980 4078
rect 275928 4014 275980 4020
rect 278056 3602 278084 233854
rect 278134 233200 278190 233209
rect 278134 233135 278190 233144
rect 278148 3806 278176 233135
rect 278240 221678 278268 310218
rect 278332 229974 278360 317319
rect 278412 313064 278464 313070
rect 278412 313006 278464 313012
rect 278320 229968 278372 229974
rect 278320 229910 278372 229916
rect 278424 228721 278452 313006
rect 278516 293418 278544 374614
rect 278608 294642 278636 374818
rect 281080 374060 281132 374066
rect 281080 374002 281132 374008
rect 279516 372020 279568 372026
rect 279516 371962 279568 371968
rect 279424 371748 279476 371754
rect 279424 371690 279476 371696
rect 279436 326398 279464 371690
rect 279528 327758 279556 371962
rect 280804 371952 280856 371958
rect 280804 371894 280856 371900
rect 280436 371816 280488 371822
rect 280436 371758 280488 371764
rect 280252 371612 280304 371618
rect 280252 371554 280304 371560
rect 279974 369880 280030 369889
rect 279974 369815 280030 369824
rect 279516 327752 279568 327758
rect 279516 327694 279568 327700
rect 279424 326392 279476 326398
rect 279424 326334 279476 326340
rect 279988 322250 280016 369815
rect 280264 366382 280292 371554
rect 280252 366376 280304 366382
rect 280252 366318 280304 366324
rect 280448 364410 280476 371758
rect 280436 364404 280488 364410
rect 280436 364346 280488 364352
rect 280712 360256 280764 360262
rect 280710 360224 280712 360233
rect 280764 360224 280766 360233
rect 280710 360159 280766 360168
rect 280710 358864 280766 358873
rect 280068 358828 280120 358834
rect 280710 358799 280712 358808
rect 280068 358770 280120 358776
rect 280764 358799 280766 358808
rect 280712 358770 280764 358776
rect 279976 322244 280028 322250
rect 279976 322186 280028 322192
rect 279884 318912 279936 318918
rect 279884 318854 279936 318860
rect 279608 318708 279660 318714
rect 279608 318650 279660 318656
rect 278688 315172 278740 315178
rect 278688 315114 278740 315120
rect 278596 294636 278648 294642
rect 278596 294578 278648 294584
rect 278504 293412 278556 293418
rect 278504 293354 278556 293360
rect 278700 236774 278728 315114
rect 279424 314424 279476 314430
rect 279424 314366 279476 314372
rect 279436 236842 279464 314366
rect 279516 311636 279568 311642
rect 279516 311578 279568 311584
rect 279424 236836 279476 236842
rect 279424 236778 279476 236784
rect 278688 236768 278740 236774
rect 278688 236710 278740 236716
rect 278780 229696 278832 229702
rect 278780 229638 278832 229644
rect 278410 228712 278466 228721
rect 278410 228647 278466 228656
rect 278792 228274 278820 229638
rect 278780 228268 278832 228274
rect 278780 228210 278832 228216
rect 278228 221672 278280 221678
rect 278228 221614 278280 221620
rect 278792 16574 278820 228210
rect 278792 16546 279096 16574
rect 278320 4072 278372 4078
rect 278320 4014 278372 4020
rect 278136 3800 278188 3806
rect 278136 3742 278188 3748
rect 275284 3596 275336 3602
rect 275284 3538 275336 3544
rect 278044 3596 278096 3602
rect 278044 3538 278096 3544
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 276032 480 276060 3470
rect 277124 3120 277176 3126
rect 277124 3062 277176 3068
rect 277136 480 277164 3062
rect 278332 480 278360 4014
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279436 4010 279464 236778
rect 279528 218793 279556 311578
rect 279620 232830 279648 318650
rect 279792 317416 279844 317422
rect 279792 317358 279844 317364
rect 279700 315240 279752 315246
rect 279700 315182 279752 315188
rect 279608 232824 279660 232830
rect 279608 232766 279660 232772
rect 279712 231198 279740 315182
rect 279804 232490 279832 317358
rect 279896 235006 279924 318854
rect 279884 235000 279936 235006
rect 279884 234942 279936 234948
rect 279792 232484 279844 232490
rect 279792 232426 279844 232432
rect 279700 231192 279752 231198
rect 279700 231134 279752 231140
rect 279514 218784 279570 218793
rect 279514 218719 279570 218728
rect 280080 100706 280108 358770
rect 280816 323610 280844 371894
rect 280896 371884 280948 371890
rect 280896 371826 280948 371832
rect 280908 324970 280936 371826
rect 280988 371680 281040 371686
rect 280988 371622 281040 371628
rect 281000 356726 281028 371622
rect 280988 356720 281040 356726
rect 280988 356662 281040 356668
rect 280896 324964 280948 324970
rect 280896 324906 280948 324912
rect 280804 323604 280856 323610
rect 280804 323546 280856 323552
rect 280804 322244 280856 322250
rect 280804 322186 280856 322192
rect 280158 320376 280214 320385
rect 280158 320311 280214 320320
rect 280172 315382 280200 320311
rect 280712 320136 280764 320142
rect 280712 320078 280764 320084
rect 280620 317620 280672 317626
rect 280620 317562 280672 317568
rect 280160 315376 280212 315382
rect 280160 315318 280212 315324
rect 280632 304434 280660 317562
rect 280620 304428 280672 304434
rect 280620 304370 280672 304376
rect 280724 293350 280752 320078
rect 280712 293344 280764 293350
rect 280712 293286 280764 293292
rect 280158 214568 280214 214577
rect 280158 214503 280214 214512
rect 280068 100700 280120 100706
rect 280068 100642 280120 100648
rect 280172 16574 280200 214503
rect 280816 60722 280844 322186
rect 280988 316532 281040 316538
rect 280988 316474 281040 316480
rect 280896 314356 280948 314362
rect 280896 314298 280948 314304
rect 280908 310298 280936 314298
rect 281000 311166 281028 316474
rect 280988 311160 281040 311166
rect 280988 311102 281040 311108
rect 280908 310270 281028 310298
rect 280896 306400 280948 306406
rect 280896 306342 280948 306348
rect 280908 219026 280936 306342
rect 281000 228585 281028 310270
rect 281092 291990 281120 374002
rect 289096 373289 289124 632062
rect 298744 630692 298796 630698
rect 298744 630634 298796 630640
rect 291844 605872 291896 605878
rect 291844 605814 291896 605820
rect 291856 380254 291884 605814
rect 295984 447840 296036 447846
rect 295984 447782 296036 447788
rect 294604 430636 294656 430642
rect 294604 430578 294656 430584
rect 291844 380248 291896 380254
rect 291844 380190 291896 380196
rect 292580 378208 292632 378214
rect 292580 378150 292632 378156
rect 292592 375374 292620 378150
rect 292316 375346 292620 375374
rect 291568 373380 291620 373386
rect 291568 373322 291620 373328
rect 289082 373280 289138 373289
rect 289082 373215 289138 373224
rect 288992 373040 289044 373046
rect 288992 372982 289044 372988
rect 281172 372632 281224 372638
rect 281172 372574 281224 372580
rect 281080 291984 281132 291990
rect 281080 291926 281132 291932
rect 281184 291922 281212 372574
rect 288256 372088 288308 372094
rect 288256 372030 288308 372036
rect 286782 371784 286838 371793
rect 286782 371719 286838 371728
rect 281262 371512 281318 371521
rect 281262 371447 281318 371456
rect 281276 358873 281304 371447
rect 282090 371376 282146 371385
rect 282000 371340 282052 371346
rect 282090 371311 282146 371320
rect 286046 371376 286102 371385
rect 286046 371311 286102 371320
rect 282000 371282 282052 371288
rect 281356 369980 281408 369986
rect 281356 369922 281408 369928
rect 281262 358864 281318 358873
rect 281262 358799 281318 358808
rect 281264 311160 281316 311166
rect 281264 311102 281316 311108
rect 281172 291916 281224 291922
rect 281172 291858 281224 291864
rect 281276 236978 281304 311102
rect 281368 291174 281396 369922
rect 281448 369912 281500 369918
rect 281448 369854 281500 369860
rect 281356 291168 281408 291174
rect 281356 291110 281408 291116
rect 281368 290494 281396 291110
rect 281356 290488 281408 290494
rect 281356 290430 281408 290436
rect 281460 287065 281488 369854
rect 282012 364334 282040 371282
rect 282104 369050 282132 371311
rect 286060 370297 286088 371311
rect 286046 370288 286102 370297
rect 286046 370223 286102 370232
rect 282276 370048 282328 370054
rect 282276 369990 282328 369996
rect 282184 369368 282236 369374
rect 282184 369310 282236 369316
rect 282196 369170 282224 369310
rect 282184 369164 282236 369170
rect 282184 369106 282236 369112
rect 282104 369022 282224 369050
rect 282012 364306 282132 364334
rect 281998 322008 282054 322017
rect 281998 321943 282054 321952
rect 281908 321020 281960 321026
rect 281908 320962 281960 320968
rect 281920 320550 281948 320962
rect 281908 320544 281960 320550
rect 281908 320486 281960 320492
rect 281906 320240 281962 320249
rect 281906 320175 281962 320184
rect 281724 319864 281776 319870
rect 281724 319806 281776 319812
rect 281736 310010 281764 319806
rect 281920 318209 281948 320175
rect 282012 319938 282040 321943
rect 282000 319932 282052 319938
rect 282000 319874 282052 319880
rect 281906 318200 281962 318209
rect 281906 318135 281962 318144
rect 281998 315208 282054 315217
rect 281998 315143 282054 315152
rect 281724 310004 281776 310010
rect 281724 309946 281776 309952
rect 282012 309398 282040 315143
rect 282000 309392 282052 309398
rect 282000 309334 282052 309340
rect 282104 306338 282132 364306
rect 282196 329089 282224 369022
rect 282288 345681 282316 369990
rect 286060 369866 286088 370223
rect 285844 369838 286088 369866
rect 286184 369880 286240 369889
rect 286184 369815 286240 369824
rect 286796 369730 286824 371719
rect 288268 371657 288296 372030
rect 288254 371648 288310 371657
rect 288254 371583 288310 371592
rect 287058 371512 287114 371521
rect 287058 371447 287114 371456
rect 287072 369866 287100 371447
rect 288024 369880 288080 369889
rect 287072 369838 287316 369866
rect 288024 369815 288080 369824
rect 288268 369730 288296 371583
rect 288532 369912 288584 369918
rect 288584 369860 288788 369866
rect 288532 369854 288788 369860
rect 288544 369838 288788 369854
rect 286796 369702 286948 369730
rect 288268 369702 288420 369730
rect 285218 369608 285274 369617
rect 289004 369594 289032 372982
rect 289268 372088 289320 372094
rect 289268 372030 289320 372036
rect 289280 371278 289308 372030
rect 290556 372020 290608 372026
rect 290556 371962 290608 371968
rect 290568 371414 290596 371962
rect 290556 371408 290608 371414
rect 290556 371350 290608 371356
rect 289268 371272 289320 371278
rect 289268 371214 289320 371220
rect 289280 369866 289308 371214
rect 290004 370660 290056 370666
rect 290004 370602 290056 370608
rect 289280 369838 289524 369866
rect 290016 369854 290044 370602
rect 290568 370138 290596 371350
rect 290568 370110 290642 370138
rect 289878 369826 290044 369854
rect 290614 369852 290642 370110
rect 291580 369986 291608 373322
rect 292212 372156 292264 372162
rect 292212 372098 292264 372104
rect 291844 371340 291896 371346
rect 291844 371282 291896 371288
rect 291568 369980 291620 369986
rect 291568 369922 291620 369928
rect 290740 369912 290792 369918
rect 290792 369860 290996 369866
rect 290740 369854 290996 369860
rect 290752 369838 290996 369854
rect 291580 369730 291608 369922
rect 291856 369866 291884 371282
rect 291856 369838 292100 369866
rect 290016 369714 290504 369730
rect 290016 369708 290516 369714
rect 290016 369702 290464 369708
rect 285274 369566 285476 369594
rect 289004 369566 289156 369594
rect 285218 369543 285274 369552
rect 283654 369472 283710 369481
rect 282368 369436 282420 369442
rect 284482 369472 284538 369481
rect 283710 369430 284004 369458
rect 284128 369442 284372 369458
rect 284116 369436 284372 369442
rect 283654 369407 283710 369416
rect 282368 369378 282420 369384
rect 284168 369430 284372 369436
rect 284942 369472 284998 369481
rect 284538 369430 284740 369458
rect 284482 369407 284538 369416
rect 287426 369472 287482 369481
rect 284998 369430 285108 369458
rect 284942 369407 284998 369416
rect 287482 369430 287684 369458
rect 290016 369442 290044 369702
rect 291364 369702 291608 369730
rect 290464 369650 290516 369656
rect 292224 369646 292252 372098
rect 291936 369640 291988 369646
rect 291732 369588 291936 369594
rect 291732 369582 291988 369588
rect 292212 369640 292264 369646
rect 292212 369582 292264 369588
rect 291732 369566 291976 369582
rect 292316 369442 292344 375346
rect 294616 374202 294644 430578
rect 294696 418192 294748 418198
rect 294696 418134 294748 418140
rect 294708 375834 294736 418134
rect 294788 404388 294840 404394
rect 294788 404330 294840 404336
rect 294696 375828 294748 375834
rect 294696 375770 294748 375776
rect 294800 374610 294828 404330
rect 295996 383654 296024 447782
rect 297364 396772 297416 396778
rect 297364 396714 297416 396720
rect 296076 387184 296128 387190
rect 296076 387126 296128 387132
rect 295904 383626 296024 383654
rect 294880 375828 294932 375834
rect 294880 375770 294932 375776
rect 294788 374604 294840 374610
rect 294788 374546 294840 374552
rect 294604 374196 294656 374202
rect 294604 374138 294656 374144
rect 294328 373584 294380 373590
rect 294328 373526 294380 373532
rect 293788 371606 294000 371634
rect 293684 371544 293736 371550
rect 293684 371486 293736 371492
rect 293696 370666 293724 371486
rect 293684 370660 293736 370666
rect 293684 370602 293736 370608
rect 292948 370524 293000 370530
rect 292948 370466 293000 370472
rect 292672 370388 292724 370394
rect 292672 370330 292724 370336
rect 292684 369594 292712 370330
rect 292960 369730 292988 370466
rect 293178 370116 293230 370122
rect 293178 370058 293230 370064
rect 293190 369852 293218 370058
rect 292836 369702 292988 369730
rect 293696 369730 293724 370602
rect 293788 370530 293816 371606
rect 293972 371550 294000 371606
rect 293960 371544 294012 371550
rect 293960 371486 294012 371492
rect 293776 370524 293828 370530
rect 293776 370466 293828 370472
rect 294340 370138 294368 373526
rect 294294 370110 294368 370138
rect 294616 370138 294644 374138
rect 294800 373590 294828 374546
rect 294788 373584 294840 373590
rect 294788 373526 294840 373532
rect 294616 370110 294690 370138
rect 294294 369852 294322 370110
rect 294662 369852 294690 370110
rect 294892 369866 294920 375770
rect 295904 374678 295932 383626
rect 296088 374882 296116 387126
rect 296720 385688 296772 385694
rect 296720 385630 296772 385636
rect 296628 376168 296680 376174
rect 296628 376110 296680 376116
rect 296076 374876 296128 374882
rect 296076 374818 296128 374824
rect 295892 374672 295944 374678
rect 295892 374614 295944 374620
rect 295524 374604 295576 374610
rect 295524 374546 295576 374552
rect 295536 372638 295564 374546
rect 295800 373652 295852 373658
rect 295800 373594 295852 373600
rect 295524 372632 295576 372638
rect 295524 372574 295576 372580
rect 294892 369838 295044 369866
rect 295536 369730 295564 372574
rect 295614 370424 295670 370433
rect 295614 370359 295670 370368
rect 295628 370161 295656 370359
rect 295614 370152 295670 370161
rect 295812 370138 295840 373594
rect 295614 370087 295670 370096
rect 295766 370110 295840 370138
rect 295766 369852 295794 370110
rect 295904 369866 295932 374614
rect 296088 373658 296116 374818
rect 296076 373652 296128 373658
rect 296076 373594 296128 373600
rect 296640 370462 296668 376110
rect 296628 370456 296680 370462
rect 296628 370398 296680 370404
rect 295904 369838 296148 369866
rect 296640 369730 296668 370398
rect 296732 370161 296760 385630
rect 297088 377528 297140 377534
rect 297088 377470 297140 377476
rect 297100 370598 297128 377470
rect 297376 375426 297404 396714
rect 298756 375562 298784 630634
rect 298836 399492 298888 399498
rect 298836 399434 298888 399440
rect 298848 375698 298876 399434
rect 298928 388544 298980 388550
rect 298928 388486 298980 388492
rect 298940 383654 298968 388486
rect 299584 386345 299612 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 305000 700324 305052 700330
rect 305000 700266 305052 700272
rect 299664 696992 299716 696998
rect 299664 696934 299716 696940
rect 299570 386336 299626 386345
rect 299570 386271 299626 386280
rect 298940 383626 299152 383654
rect 298928 377460 298980 377466
rect 298928 377402 298980 377408
rect 298836 375692 298888 375698
rect 298836 375634 298888 375640
rect 298744 375556 298796 375562
rect 298744 375498 298796 375504
rect 298756 375426 298784 375498
rect 297364 375420 297416 375426
rect 297364 375362 297416 375368
rect 298744 375420 298796 375426
rect 298744 375362 298796 375368
rect 297088 370592 297140 370598
rect 297088 370534 297140 370540
rect 296718 370152 296774 370161
rect 296718 370087 296774 370096
rect 297100 369866 297128 370534
rect 297376 369866 297404 375362
rect 298848 375034 298876 375634
rect 298572 375006 298876 375034
rect 297824 374876 297876 374882
rect 297824 374818 297876 374824
rect 297836 374066 297864 374818
rect 297824 374060 297876 374066
rect 297824 374002 297876 374008
rect 296884 369838 297128 369866
rect 297252 369838 297404 369866
rect 297836 369730 297864 374002
rect 297960 370152 298016 370161
rect 297960 370087 298016 370096
rect 297974 369852 298002 370087
rect 298572 369866 298600 375006
rect 298940 371385 298968 377402
rect 299124 374241 299152 383626
rect 299388 375420 299440 375426
rect 299388 375362 299440 375368
rect 299110 374232 299166 374241
rect 299110 374167 299166 374176
rect 298926 371376 298982 371385
rect 298926 371311 298982 371320
rect 298940 369866 298968 371311
rect 299124 370138 299152 374167
rect 299296 371340 299348 371346
rect 299296 371282 299348 371288
rect 298356 369838 298600 369866
rect 298724 369838 298968 369866
rect 299078 370110 299152 370138
rect 299078 369852 299106 370110
rect 293696 369702 293940 369730
rect 295412 369702 295564 369730
rect 296516 369702 296668 369730
rect 297620 369702 297864 369730
rect 292468 369566 292712 369594
rect 299308 369481 299336 371282
rect 299400 370138 299428 375362
rect 299480 371408 299532 371414
rect 299480 371350 299532 371356
rect 299492 370598 299520 371350
rect 299480 370592 299532 370598
rect 299480 370534 299532 370540
rect 299676 370433 299704 696934
rect 300124 683256 300176 683262
rect 300124 683198 300176 683204
rect 299756 380180 299808 380186
rect 299756 380122 299808 380128
rect 299768 374474 299796 380122
rect 300136 379514 300164 683198
rect 302884 618316 302936 618322
rect 302884 618258 302936 618264
rect 302896 395418 302924 618258
rect 304264 402280 304316 402286
rect 304264 402222 304316 402228
rect 302976 400920 303028 400926
rect 302976 400862 303028 400868
rect 302884 395412 302936 395418
rect 302884 395354 302936 395360
rect 301504 393984 301556 393990
rect 301504 393926 301556 393932
rect 301044 384328 301096 384334
rect 301044 384270 301096 384276
rect 300136 379486 300348 379514
rect 300320 375494 300348 379486
rect 300308 375488 300360 375494
rect 300308 375430 300360 375436
rect 299756 374468 299808 374474
rect 299756 374410 299808 374416
rect 299662 370424 299718 370433
rect 299662 370359 299718 370368
rect 299676 370161 299704 370359
rect 299662 370152 299718 370161
rect 299400 370110 299474 370138
rect 299446 369852 299474 370110
rect 299768 370138 299796 374410
rect 300168 370152 300224 370161
rect 299768 370110 299842 370138
rect 299662 370087 299718 370096
rect 299814 369852 299842 370110
rect 300168 370087 300224 370096
rect 300182 369852 300210 370087
rect 300320 369866 300348 375430
rect 300768 374400 300820 374406
rect 300768 374342 300820 374348
rect 300320 369838 300564 369866
rect 300780 369594 300808 374342
rect 301056 370569 301084 384270
rect 301516 375737 301544 393926
rect 302884 391264 302936 391270
rect 302884 391206 302936 391212
rect 301780 381540 301832 381546
rect 301780 381482 301832 381488
rect 301502 375728 301558 375737
rect 301502 375663 301558 375672
rect 301042 370560 301098 370569
rect 301042 370495 301098 370504
rect 301056 369866 301084 370495
rect 301516 369866 301544 375663
rect 301056 369838 301300 369866
rect 301516 369838 301668 369866
rect 300780 369566 300932 369594
rect 301792 369481 301820 381482
rect 302606 375592 302662 375601
rect 302606 375527 302662 375536
rect 302330 371648 302386 371657
rect 302330 371583 302386 371592
rect 302240 370796 302292 370802
rect 302240 370738 302292 370744
rect 302252 369866 302280 370738
rect 302344 370666 302372 371583
rect 302332 370660 302384 370666
rect 302332 370602 302384 370608
rect 302620 369866 302648 375527
rect 302896 370326 302924 391206
rect 302988 375601 303016 400862
rect 303252 389836 303304 389842
rect 303252 389778 303304 389784
rect 303160 376100 303212 376106
rect 303160 376042 303212 376048
rect 302974 375592 303030 375601
rect 302974 375527 303030 375536
rect 303172 374406 303200 376042
rect 303160 374400 303212 374406
rect 303160 374342 303212 374348
rect 303264 370802 303292 389778
rect 303344 383036 303396 383042
rect 303344 382978 303396 382984
rect 303252 370796 303304 370802
rect 303252 370738 303304 370744
rect 302884 370320 302936 370326
rect 302884 370262 302936 370268
rect 302252 369838 302404 369866
rect 302620 369838 302772 369866
rect 302896 369753 302924 370262
rect 302882 369744 302938 369753
rect 302882 369679 302938 369688
rect 299294 369472 299350 369481
rect 293328 369442 293572 369458
rect 290004 369436 290056 369442
rect 287426 369407 287482 369416
rect 284116 369378 284168 369384
rect 290004 369378 290056 369384
rect 292304 369436 292356 369442
rect 292304 369378 292356 369384
rect 293316 369436 293572 369442
rect 293368 369430 293572 369436
rect 299294 369407 299350 369416
rect 301778 369472 301834 369481
rect 302882 369472 302938 369481
rect 301834 369430 302036 369458
rect 301778 369407 301834 369416
rect 303356 369458 303384 382978
rect 304276 375630 304304 402222
rect 304356 398132 304408 398138
rect 304356 398074 304408 398080
rect 304264 375624 304316 375630
rect 304264 375566 304316 375572
rect 304368 374746 304396 398074
rect 304448 392692 304500 392698
rect 304448 392634 304500 392640
rect 304460 379514 304488 392634
rect 304460 379486 304580 379514
rect 304552 374814 304580 379486
rect 304724 375624 304776 375630
rect 304724 375566 304776 375572
rect 304540 374808 304592 374814
rect 304540 374750 304592 374756
rect 304356 374740 304408 374746
rect 304356 374682 304408 374688
rect 304368 373538 304396 374682
rect 304092 373510 304396 373538
rect 304092 369866 304120 373510
rect 304448 373380 304500 373386
rect 304448 373322 304500 373328
rect 303876 369838 304120 369866
rect 303480 369744 303536 369753
rect 303480 369679 303536 369688
rect 302938 369430 303384 369458
rect 303986 369472 304042 369481
rect 302882 369407 302938 369416
rect 304460 369458 304488 373322
rect 304552 370138 304580 374750
rect 304552 370110 304626 370138
rect 304598 369852 304626 370110
rect 304736 369866 304764 375566
rect 305012 372230 305040 700266
rect 306380 698964 306432 698970
rect 306380 698906 306432 698912
rect 305644 397520 305696 397526
rect 305644 397462 305696 397468
rect 305656 385665 305684 397462
rect 305642 385656 305698 385665
rect 305642 385591 305698 385600
rect 305552 383104 305604 383110
rect 305552 383046 305604 383052
rect 305000 372224 305052 372230
rect 305000 372166 305052 372172
rect 305564 369866 305592 383046
rect 306392 375902 306420 698906
rect 310520 683188 310572 683194
rect 310520 683130 310572 683136
rect 309600 409896 309652 409902
rect 309600 409838 309652 409844
rect 309140 407788 309192 407794
rect 309140 407730 309192 407736
rect 306472 394052 306524 394058
rect 306472 393994 306524 394000
rect 306484 383654 306512 393994
rect 307760 392624 307812 392630
rect 307760 392566 307812 392572
rect 306484 383626 306604 383654
rect 306380 375896 306432 375902
rect 306380 375838 306432 375844
rect 306392 375426 306420 375838
rect 306380 375420 306432 375426
rect 306380 375362 306432 375368
rect 305828 372224 305880 372230
rect 305828 372166 305880 372172
rect 305840 369866 305868 372166
rect 306576 370258 306604 383626
rect 306932 375420 306984 375426
rect 306932 375362 306984 375368
rect 306564 370252 306616 370258
rect 306564 370194 306616 370200
rect 306576 369866 306604 370194
rect 306944 369866 306972 375362
rect 307772 372570 307800 392566
rect 307852 387116 307904 387122
rect 307852 387058 307904 387064
rect 307760 372564 307812 372570
rect 307760 372506 307812 372512
rect 307864 372042 307892 387058
rect 307944 382968 307996 382974
rect 307944 382910 307996 382916
rect 307956 372609 307984 382910
rect 309152 375766 309180 407730
rect 309612 403646 309640 409838
rect 309600 403640 309652 403646
rect 309600 403582 309652 403588
rect 309232 388476 309284 388482
rect 309232 388418 309284 388424
rect 309244 383654 309272 388418
rect 309244 383626 310008 383654
rect 309140 375760 309192 375766
rect 309140 375702 309192 375708
rect 309152 375426 309180 375702
rect 309140 375420 309192 375426
rect 309140 375362 309192 375368
rect 307942 372600 307998 372609
rect 309598 372600 309654 372609
rect 307942 372535 307998 372544
rect 308036 372564 308088 372570
rect 309598 372535 309654 372544
rect 308036 372506 308088 372512
rect 307680 372014 307892 372042
rect 307680 370190 307708 372014
rect 308048 371482 308076 372506
rect 308036 371476 308088 371482
rect 308036 371418 308088 371424
rect 308864 371476 308916 371482
rect 308864 371418 308916 371424
rect 307668 370184 307720 370190
rect 307668 370126 307720 370132
rect 304736 369838 304980 369866
rect 305564 369838 305716 369866
rect 305840 369838 306084 369866
rect 306576 369838 306820 369866
rect 306944 369838 307188 369866
rect 307680 369594 307708 370126
rect 308048 369866 308076 371418
rect 308048 369838 308292 369866
rect 308402 369744 308458 369753
rect 308458 369702 308660 369730
rect 308402 369679 308458 369688
rect 307680 369566 307924 369594
rect 308876 369510 308904 371418
rect 309368 369744 309424 369753
rect 309368 369679 309424 369688
rect 308864 369504 308916 369510
rect 305458 369472 305514 369481
rect 304042 369430 304488 369458
rect 305348 369430 305458 369458
rect 303986 369407 304042 369416
rect 307298 369472 307354 369481
rect 306300 369442 306452 369458
rect 305458 369407 305514 369416
rect 306288 369436 306452 369442
rect 293316 369378 293368 369384
rect 306340 369430 306452 369436
rect 307354 369430 307556 369458
rect 308864 369446 308916 369452
rect 309612 369458 309640 372535
rect 309874 369472 309930 369481
rect 309612 369430 309874 369458
rect 307298 369407 307354 369416
rect 309980 369458 310008 383626
rect 310244 375420 310296 375426
rect 310244 375362 310296 375368
rect 310256 369866 310284 375362
rect 310532 374626 310560 683130
rect 310612 670744 310664 670750
rect 310612 670686 310664 670692
rect 330484 670744 330536 670750
rect 330484 670686 330536 670692
rect 310624 374762 310652 670686
rect 310704 656940 310756 656946
rect 310704 656882 310756 656888
rect 310716 379514 310744 656882
rect 323584 643136 323636 643142
rect 323584 643078 323636 643084
rect 313280 565888 313332 565894
rect 313280 565830 313332 565836
rect 311900 395412 311952 395418
rect 311900 395354 311952 395360
rect 310716 379486 311020 379514
rect 310624 374734 310744 374762
rect 310532 374598 310652 374626
rect 310256 369838 310500 369866
rect 310104 369472 310160 369481
rect 309980 369430 310104 369458
rect 309874 369407 309930 369416
rect 310624 369458 310652 374598
rect 310716 372609 310744 374734
rect 310992 374105 311020 379486
rect 311912 375465 311940 395354
rect 312084 380248 312136 380254
rect 312084 380190 312136 380196
rect 311898 375456 311954 375465
rect 311898 375391 311954 375400
rect 310978 374096 311034 374105
rect 310978 374031 311034 374040
rect 310702 372600 310758 372609
rect 310702 372535 310758 372544
rect 310992 369866 311020 374031
rect 311714 373280 311770 373289
rect 311714 373215 311770 373224
rect 311346 372600 311402 372609
rect 311346 372535 311402 372544
rect 311360 371929 311388 372535
rect 311346 371920 311402 371929
rect 311346 371855 311402 371864
rect 311360 369866 311388 371855
rect 311728 369866 311756 373215
rect 310992 369838 311236 369866
rect 311360 369838 311604 369866
rect 311728 369838 311972 369866
rect 311728 369753 311756 369838
rect 311714 369744 311770 369753
rect 311714 369679 311770 369688
rect 312096 369481 312124 380190
rect 312820 376032 312872 376038
rect 312820 375974 312872 375980
rect 312450 375456 312506 375465
rect 312450 375391 312506 375400
rect 312464 369866 312492 375391
rect 312464 369838 312708 369866
rect 312832 369617 312860 375974
rect 313292 374406 313320 565830
rect 319444 563100 319496 563106
rect 319444 563042 319496 563048
rect 318064 510672 318116 510678
rect 318064 510614 318116 510620
rect 314752 462392 314804 462398
rect 314752 462334 314804 462340
rect 313372 395344 313424 395350
rect 313372 395286 313424 395292
rect 313280 374400 313332 374406
rect 313280 374342 313332 374348
rect 313384 374218 313412 395286
rect 313464 374400 313516 374406
rect 313464 374342 313516 374348
rect 313292 374190 313412 374218
rect 313292 369617 313320 374190
rect 313476 371686 313504 374342
rect 313740 373244 313792 373250
rect 313740 373186 313792 373192
rect 313752 372026 313780 373186
rect 313740 372020 313792 372026
rect 313740 371962 313792 371968
rect 314764 371958 314792 462334
rect 314844 406428 314896 406434
rect 314844 406370 314896 406376
rect 314752 371952 314804 371958
rect 314752 371894 314804 371900
rect 313464 371680 313516 371686
rect 313464 371622 313516 371628
rect 313476 370138 313504 371622
rect 314856 371414 314884 406370
rect 316040 403640 316092 403646
rect 316040 403582 316092 403588
rect 314936 390584 314988 390590
rect 314936 390526 314988 390532
rect 314948 383654 314976 390526
rect 314948 383626 315436 383654
rect 314844 371408 314896 371414
rect 314844 371350 314896 371356
rect 314568 371272 314620 371278
rect 314568 371214 314620 371220
rect 314580 370734 314608 371214
rect 314568 370728 314620 370734
rect 314568 370670 314620 370676
rect 314856 370138 314884 371350
rect 313476 370110 313596 370138
rect 314856 370110 314930 370138
rect 313568 369866 313596 370110
rect 313568 369838 313812 369866
rect 314902 369852 314930 370110
rect 315408 369866 315436 383626
rect 315764 371952 315816 371958
rect 315764 371894 315816 371900
rect 315776 369866 315804 371894
rect 316052 371890 316080 403582
rect 316132 384396 316184 384402
rect 316132 384338 316184 384344
rect 316040 371884 316092 371890
rect 316040 371826 316092 371832
rect 316144 371482 316172 384338
rect 318076 376174 318104 510614
rect 318064 376168 318116 376174
rect 318064 376110 318116 376116
rect 319456 374882 319484 563042
rect 320824 536852 320876 536858
rect 320824 536794 320876 536800
rect 320836 377534 320864 536794
rect 322204 484424 322256 484430
rect 322204 484366 322256 484372
rect 322216 387190 322244 484366
rect 323596 388550 323624 643078
rect 324964 590708 325016 590714
rect 324964 590650 325016 590656
rect 323584 388544 323636 388550
rect 323584 388486 323636 388492
rect 322204 387184 322256 387190
rect 322204 387126 322256 387132
rect 324976 385694 325004 590650
rect 329104 524476 329156 524482
rect 329104 524418 329156 524424
rect 329116 396778 329144 524418
rect 329104 396772 329156 396778
rect 329104 396714 329156 396720
rect 324964 385688 325016 385694
rect 324964 385630 325016 385636
rect 330496 380186 330524 670686
rect 331232 392698 331260 702986
rect 348804 700330 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 340144 700324 340196 700330
rect 340144 700266 340196 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 334624 576904 334676 576910
rect 334624 576846 334676 576852
rect 334636 399498 334664 576846
rect 340156 402286 340184 700266
rect 363604 616888 363656 616894
rect 363604 616830 363656 616836
rect 340144 402280 340196 402286
rect 340144 402222 340196 402228
rect 334624 399492 334676 399498
rect 334624 399434 334676 399440
rect 331220 392692 331272 392698
rect 331220 392634 331272 392640
rect 330484 380180 330536 380186
rect 330484 380122 330536 380128
rect 320824 377528 320876 377534
rect 320824 377470 320876 377476
rect 363616 377466 363644 616830
rect 363604 377460 363656 377466
rect 363604 377402 363656 377408
rect 322388 376780 322440 376786
rect 322388 376722 322440 376728
rect 319444 374876 319496 374882
rect 319444 374818 319496 374824
rect 319076 374536 319128 374542
rect 319076 374478 319128 374484
rect 317328 373176 317380 373182
rect 317328 373118 317380 373124
rect 317236 373108 317288 373114
rect 317236 373050 317288 373056
rect 316868 371884 316920 371890
rect 316868 371826 316920 371832
rect 316132 371476 316184 371482
rect 316132 371418 316184 371424
rect 316144 369866 316172 371418
rect 316880 369866 316908 371826
rect 317248 369866 317276 373050
rect 317340 371482 317368 373118
rect 318800 372972 318852 372978
rect 318800 372914 318852 372920
rect 317972 371816 318024 371822
rect 317972 371758 318024 371764
rect 317328 371476 317380 371482
rect 317328 371418 317380 371424
rect 317604 370048 317656 370054
rect 317604 369990 317656 369996
rect 317616 369866 317644 369990
rect 317984 369866 318012 371758
rect 318340 371476 318392 371482
rect 318340 371418 318392 371424
rect 318352 369866 318380 371418
rect 318812 369866 318840 372914
rect 319088 369866 319116 374478
rect 319812 374332 319864 374338
rect 319812 374274 319864 374280
rect 319534 372872 319590 372881
rect 319534 372807 319590 372816
rect 319548 371278 319576 372807
rect 319444 371272 319496 371278
rect 319444 371214 319496 371220
rect 319536 371272 319588 371278
rect 319536 371214 319588 371220
rect 319456 369866 319484 371214
rect 319824 369866 319852 374274
rect 320180 374128 320232 374134
rect 320180 374070 320232 374076
rect 320192 369866 320220 374070
rect 320548 372836 320600 372842
rect 320548 372778 320600 372784
rect 320560 369866 320588 372778
rect 321652 372768 321704 372774
rect 321652 372710 321704 372716
rect 321284 371748 321336 371754
rect 321284 371690 321336 371696
rect 321296 369866 321324 371690
rect 321664 369866 321692 372710
rect 322020 372020 322072 372026
rect 322020 371962 322072 371968
rect 322032 369866 322060 371962
rect 322400 369866 322428 376722
rect 323124 374944 323176 374950
rect 323124 374886 323176 374892
rect 322940 372904 322992 372910
rect 322940 372846 322992 372852
rect 322952 370138 322980 372846
rect 322952 370110 323026 370138
rect 315408 369838 315652 369866
rect 315776 369838 316020 369866
rect 316144 369838 316388 369866
rect 316880 369838 317124 369866
rect 317248 369838 317492 369866
rect 317616 369838 317860 369866
rect 317984 369838 318228 369866
rect 318352 369838 318596 369866
rect 318812 369838 318964 369866
rect 319088 369838 319332 369866
rect 319456 369838 319700 369866
rect 319824 369838 320068 369866
rect 320192 369838 320436 369866
rect 320560 369838 320804 369866
rect 321296 369838 321540 369866
rect 321664 369838 321908 369866
rect 322032 369838 322276 369866
rect 322400 369838 322644 369866
rect 322998 369852 323026 370110
rect 323136 369866 323164 374886
rect 325332 374264 325384 374270
rect 325332 374206 325384 374212
rect 324962 372736 325018 372745
rect 323492 372700 323544 372706
rect 324962 372671 325018 372680
rect 323492 372642 323544 372648
rect 323504 369866 323532 372642
rect 324596 371612 324648 371618
rect 324596 371554 324648 371560
rect 323860 371272 323912 371278
rect 323860 371214 323912 371220
rect 323872 369866 323900 371214
rect 324608 369866 324636 371554
rect 324976 369866 325004 372671
rect 325344 369866 325372 374206
rect 364352 373386 364380 702406
rect 397472 699718 397500 703520
rect 413664 700330 413692 703520
rect 403624 700324 403676 700330
rect 403624 700266 403676 700272
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 414664 700324 414716 700330
rect 414664 700266 414716 700272
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 396736 391270 396764 699654
rect 399484 470620 399536 470626
rect 399484 470562 399536 470568
rect 399496 447846 399524 470562
rect 399484 447840 399536 447846
rect 399484 447782 399536 447788
rect 403636 398138 403664 700266
rect 414676 400926 414704 700266
rect 414664 400920 414716 400926
rect 414664 400862 414716 400868
rect 403624 398132 403676 398138
rect 403624 398074 403676 398080
rect 396724 391264 396776 391270
rect 396724 391206 396776 391212
rect 429212 383042 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 389842 462360 703520
rect 478524 700330 478552 703520
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 462320 389836 462372 389842
rect 462320 389778 462372 389784
rect 429200 383036 429252 383042
rect 429200 382978 429252 382984
rect 494072 381546 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 699718 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 526444 699712 526496 699718
rect 526444 699654 526496 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 526456 384334 526484 699654
rect 542372 393990 542400 702406
rect 542360 393984 542412 393990
rect 542360 393926 542412 393932
rect 526444 384328 526496 384334
rect 526444 384270 526496 384276
rect 494060 381540 494112 381546
rect 494060 381482 494112 381488
rect 558932 376106 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 558920 376100 558972 376106
rect 558920 376042 558972 376048
rect 580276 374678 580304 458079
rect 580264 374672 580316 374678
rect 580264 374614 580316 374620
rect 364340 373380 364392 373386
rect 364340 373322 364392 373328
rect 577596 373040 577648 373046
rect 577596 372982 577648 372988
rect 363604 372156 363656 372162
rect 363604 372098 363656 372104
rect 336004 371544 336056 371550
rect 336004 371486 336056 371492
rect 329104 370388 329156 370394
rect 329104 370330 329156 370336
rect 323136 369838 323380 369866
rect 323504 369838 323748 369866
rect 323872 369838 324116 369866
rect 324608 369838 324852 369866
rect 324976 369838 325220 369866
rect 325344 369838 325588 369866
rect 312818 369608 312874 369617
rect 313278 369608 313334 369617
rect 312874 369566 313076 369594
rect 312818 369543 312874 369552
rect 313278 369543 313334 369552
rect 314520 369608 314576 369617
rect 314520 369543 314576 369552
rect 310978 369472 311034 369481
rect 310624 369430 310978 369458
rect 310104 369407 310160 369416
rect 310978 369407 311034 369416
rect 312082 369472 312138 369481
rect 312082 369407 312138 369416
rect 313922 369472 313978 369481
rect 315026 369472 315082 369481
rect 313978 369430 314180 369458
rect 313922 369407 313978 369416
rect 320914 369472 320970 369481
rect 315082 369430 315284 369458
rect 315026 369407 315082 369416
rect 324226 369472 324282 369481
rect 320970 369430 321172 369458
rect 320914 369407 320970 369416
rect 324282 369430 324484 369458
rect 325956 369442 326292 369458
rect 325956 369436 326304 369442
rect 325956 369430 326252 369436
rect 324226 369407 324282 369416
rect 306288 369378 306340 369384
rect 326252 369378 326304 369384
rect 329012 369436 329064 369442
rect 329012 369378 329064 369384
rect 282380 363633 282408 369378
rect 286552 369336 286608 369345
rect 286552 369271 286608 369280
rect 309000 369336 309056 369345
rect 309000 369271 309056 369280
rect 310104 369336 310160 369345
rect 310104 369271 310160 369280
rect 312312 369336 312368 369345
rect 312312 369271 312368 369280
rect 313416 369336 313472 369345
rect 313416 369271 313472 369280
rect 316728 369336 316784 369345
rect 316728 369271 316784 369280
rect 282460 369232 282512 369238
rect 282460 369174 282512 369180
rect 282472 368830 282500 369174
rect 282460 368824 282512 368830
rect 282460 368766 282512 368772
rect 282366 363624 282422 363633
rect 282366 363559 282422 363568
rect 282274 345672 282330 345681
rect 282274 345607 282330 345616
rect 282182 329080 282238 329089
rect 282182 329015 282238 329024
rect 282274 322144 282330 322153
rect 282274 322079 282330 322088
rect 282288 320754 282316 322079
rect 327722 321328 327778 321337
rect 327722 321263 327778 321272
rect 327538 320920 327594 320929
rect 327538 320855 327594 320864
rect 288024 320784 288080 320793
rect 283714 320754 283742 320756
rect 282276 320748 282328 320754
rect 282276 320690 282328 320696
rect 283702 320748 283754 320754
rect 288024 320719 288080 320728
rect 290140 320784 290196 320793
rect 290140 320719 290196 320728
rect 293452 320784 293508 320793
rect 293452 320719 293508 320728
rect 294096 320784 294152 320793
rect 294096 320719 294152 320728
rect 295384 320784 295440 320793
rect 295384 320719 295440 320728
rect 299432 320784 299488 320793
rect 311208 320784 311264 320793
rect 299432 320719 299488 320728
rect 283702 320690 283754 320696
rect 302942 320686 302970 320756
rect 311208 320719 311264 320728
rect 323352 320784 323408 320793
rect 323352 320719 323408 320728
rect 324456 320784 324512 320793
rect 324456 320719 324512 320728
rect 282184 320680 282236 320686
rect 282184 320622 282236 320628
rect 302930 320680 302982 320686
rect 302930 320622 302982 320628
rect 311944 320648 312000 320657
rect 282196 320414 282224 320622
rect 285830 320618 285858 320620
rect 285818 320612 285870 320618
rect 311944 320583 312000 320592
rect 313140 320648 313196 320657
rect 313140 320583 313196 320592
rect 322800 320648 322856 320657
rect 322800 320583 322856 320592
rect 325008 320648 325064 320657
rect 325008 320583 325064 320592
rect 285818 320554 285870 320560
rect 315072 320512 315128 320521
rect 315072 320447 315128 320456
rect 317648 320512 317704 320521
rect 317648 320447 317704 320456
rect 318844 320512 318900 320521
rect 318844 320447 318900 320456
rect 323904 320512 323960 320521
rect 323904 320447 323960 320456
rect 325560 320512 325616 320521
rect 325560 320447 325616 320456
rect 282184 320408 282236 320414
rect 282184 320350 282236 320356
rect 282964 320376 283020 320385
rect 282964 320311 283020 320320
rect 283240 320376 283296 320385
rect 283240 320311 283296 320320
rect 283792 320376 283848 320385
rect 283792 320311 283848 320320
rect 289680 320376 289736 320385
rect 289680 320311 289736 320320
rect 291060 320376 291116 320385
rect 297684 320376 297740 320385
rect 292454 320346 292482 320348
rect 291060 320311 291116 320320
rect 292442 320340 292494 320346
rect 297684 320311 297740 320320
rect 298052 320376 298108 320385
rect 298052 320311 298108 320320
rect 298604 320376 298660 320385
rect 298604 320311 298660 320320
rect 300628 320376 300684 320385
rect 300628 320311 300684 320320
rect 308908 320376 308964 320385
rect 308908 320311 308964 320320
rect 312220 320376 312276 320385
rect 312220 320311 312276 320320
rect 313232 320376 313288 320385
rect 313232 320311 313288 320320
rect 317096 320376 317152 320385
rect 317096 320311 317152 320320
rect 318752 320376 318808 320385
rect 318752 320311 318808 320320
rect 318936 320376 318992 320385
rect 318936 320311 318992 320320
rect 323168 320376 323224 320385
rect 323168 320311 323224 320320
rect 326664 320376 326720 320385
rect 326664 320311 326720 320320
rect 292442 320282 292494 320288
rect 285172 320240 285228 320249
rect 285172 320175 285228 320184
rect 286460 320240 286516 320249
rect 286460 320175 286516 320184
rect 286644 320240 286700 320249
rect 286644 320175 286700 320184
rect 287380 320240 287436 320249
rect 287380 320175 287436 320184
rect 288116 320240 288172 320249
rect 288116 320175 288172 320184
rect 289036 320240 289092 320249
rect 289036 320175 289092 320184
rect 290324 320240 290380 320249
rect 290324 320175 290380 320184
rect 290968 320240 291024 320249
rect 290968 320175 291024 320184
rect 291336 320240 291392 320249
rect 291336 320175 291392 320184
rect 293544 320240 293600 320249
rect 293544 320175 293600 320184
rect 294188 320240 294244 320249
rect 294188 320175 294244 320184
rect 296856 320240 296912 320249
rect 296856 320175 296912 320184
rect 297776 320240 297832 320249
rect 297776 320175 297832 320184
rect 299340 320240 299396 320249
rect 299340 320175 299396 320184
rect 300996 320240 301052 320249
rect 300996 320175 301052 320184
rect 304216 320240 304272 320249
rect 304216 320175 304272 320184
rect 308448 320240 308504 320249
rect 308448 320175 308504 320184
rect 309920 320240 309976 320249
rect 309920 320175 309976 320184
rect 310840 320240 310896 320249
rect 310840 320175 310896 320184
rect 311668 320240 311724 320249
rect 311668 320175 311724 320184
rect 312404 320240 312460 320249
rect 312404 320175 312460 320184
rect 312956 320240 313012 320249
rect 312956 320175 313012 320184
rect 314336 320240 314392 320249
rect 314336 320175 314392 320184
rect 316268 320240 316324 320249
rect 316268 320175 316324 320184
rect 316544 320240 316600 320249
rect 316544 320175 316600 320184
rect 317280 320240 317336 320249
rect 317280 320175 317336 320184
rect 318384 320240 318440 320249
rect 318384 320175 318440 320184
rect 320132 320240 320188 320249
rect 320132 320175 320188 320184
rect 321420 320240 321476 320249
rect 321420 320175 321476 320184
rect 322064 320240 322120 320249
rect 322064 320175 322120 320184
rect 323076 320240 323132 320249
rect 323076 320175 323132 320184
rect 324272 320240 324328 320249
rect 324272 320175 324328 320184
rect 326112 320240 326168 320249
rect 327552 320210 327580 320855
rect 327632 320816 327684 320822
rect 327632 320758 327684 320764
rect 327644 320278 327672 320758
rect 327736 320482 327764 321263
rect 328550 320784 328606 320793
rect 328550 320719 328606 320728
rect 328184 320680 328236 320686
rect 328184 320622 328236 320628
rect 327724 320476 327776 320482
rect 327724 320418 327776 320424
rect 327632 320272 327684 320278
rect 327632 320214 327684 320220
rect 326112 320175 326168 320184
rect 327540 320204 327592 320210
rect 327540 320146 327592 320152
rect 321698 320136 321750 320142
rect 282274 320104 282330 320113
rect 282872 320104 282928 320113
rect 282274 320039 282330 320048
rect 282184 318640 282236 318646
rect 282184 318582 282236 318588
rect 282092 306332 282144 306338
rect 282092 306274 282144 306280
rect 282104 305726 282132 306274
rect 282092 305720 282144 305726
rect 282092 305662 282144 305668
rect 281446 287056 281502 287065
rect 281446 286991 281502 287000
rect 281460 286385 281488 286991
rect 281446 286376 281502 286385
rect 281446 286311 281502 286320
rect 281264 236972 281316 236978
rect 281264 236914 281316 236920
rect 281540 235408 281592 235414
rect 281540 235350 281592 235356
rect 280986 228576 281042 228585
rect 280986 228511 281042 228520
rect 280896 219020 280948 219026
rect 280896 218962 280948 218968
rect 281170 214568 281226 214577
rect 281170 214503 281226 214512
rect 281184 213897 281212 214503
rect 281170 213888 281226 213897
rect 281170 213823 281226 213832
rect 280804 60716 280856 60722
rect 280804 60658 280856 60664
rect 280172 16546 280752 16574
rect 279424 4004 279476 4010
rect 279424 3946 279476 3952
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 235350
rect 282196 216510 282224 318582
rect 282288 318442 282316 320039
rect 282518 319818 282546 320076
rect 282472 319790 282546 319818
rect 282366 319288 282422 319297
rect 282366 319223 282422 319232
rect 282276 318436 282328 318442
rect 282276 318378 282328 318384
rect 282380 318016 282408 319223
rect 282472 318753 282500 319790
rect 282610 319716 282638 320076
rect 282702 319870 282730 320076
rect 282690 319864 282742 319870
rect 282690 319806 282742 319812
rect 282794 319818 282822 320076
rect 282872 320039 282928 320048
rect 283056 320104 283112 320113
rect 284160 320104 284216 320113
rect 283056 320039 283112 320048
rect 283162 319818 283190 320076
rect 283346 319938 283374 320076
rect 283334 319932 283386 319938
rect 283334 319874 283386 319880
rect 283438 319818 283466 320076
rect 283530 319938 283558 320076
rect 283518 319932 283570 319938
rect 283518 319874 283570 319880
rect 282794 319790 282868 319818
rect 283162 319790 283328 319818
rect 282564 319688 282638 319716
rect 282458 318744 282514 318753
rect 282458 318679 282514 318688
rect 282564 318617 282592 319688
rect 282550 318608 282606 318617
rect 282550 318543 282606 318552
rect 282840 318510 282868 319790
rect 283196 319728 283248 319734
rect 283196 319670 283248 319676
rect 282828 318504 282880 318510
rect 282828 318446 282880 318452
rect 282644 318436 282696 318442
rect 282644 318378 282696 318384
rect 282550 318200 282606 318209
rect 282550 318135 282606 318144
rect 282380 317988 282500 318016
rect 282366 317928 282422 317937
rect 282366 317863 282422 317872
rect 282274 310448 282330 310457
rect 282274 310383 282330 310392
rect 282288 309913 282316 310383
rect 282274 309904 282330 309913
rect 282274 309839 282330 309848
rect 282276 309528 282328 309534
rect 282276 309470 282328 309476
rect 282288 226001 282316 309470
rect 282274 225992 282330 226001
rect 282274 225927 282330 225936
rect 282380 221814 282408 317863
rect 282472 233986 282500 317988
rect 282564 312730 282592 318135
rect 282552 312724 282604 312730
rect 282552 312666 282604 312672
rect 282552 312588 282604 312594
rect 282552 312530 282604 312536
rect 282564 309534 282592 312530
rect 282656 311250 282684 318378
rect 282828 316668 282880 316674
rect 282828 316610 282880 316616
rect 282656 311222 282776 311250
rect 282644 311160 282696 311166
rect 282644 311102 282696 311108
rect 282552 309528 282604 309534
rect 282552 309470 282604 309476
rect 282552 309392 282604 309398
rect 282552 309334 282604 309340
rect 282460 233980 282512 233986
rect 282460 233922 282512 233928
rect 282564 231334 282592 309334
rect 282656 235550 282684 311102
rect 282748 236366 282776 311222
rect 282736 236360 282788 236366
rect 282736 236302 282788 236308
rect 282644 235544 282696 235550
rect 282644 235486 282696 235492
rect 282840 235414 282868 316610
rect 283104 316124 283156 316130
rect 283104 316066 283156 316072
rect 283012 316056 283064 316062
rect 283012 315998 283064 316004
rect 282920 315444 282972 315450
rect 282920 315386 282972 315392
rect 282932 315110 282960 315386
rect 282920 315104 282972 315110
rect 282920 315046 282972 315052
rect 283024 311506 283052 315998
rect 283012 311500 283064 311506
rect 283012 311442 283064 311448
rect 283116 297673 283144 316066
rect 283208 307290 283236 319670
rect 283300 307465 283328 319790
rect 283392 319790 283466 319818
rect 283286 307456 283342 307465
rect 283286 307391 283342 307400
rect 283196 307284 283248 307290
rect 283196 307226 283248 307232
rect 283102 297664 283158 297673
rect 283102 297599 283158 297608
rect 283392 296002 283420 319790
rect 283622 319784 283650 320076
rect 283748 319932 283800 319938
rect 283748 319874 283800 319880
rect 283576 319756 283650 319784
rect 283470 319288 283526 319297
rect 283470 319223 283526 319232
rect 283484 319122 283512 319223
rect 283472 319116 283524 319122
rect 283472 319058 283524 319064
rect 283576 316010 283604 319756
rect 283760 318374 283788 319874
rect 283898 319716 283926 320076
rect 283990 319938 284018 320076
rect 284082 319954 284110 320076
rect 284712 320104 284768 320113
rect 284160 320039 284216 320048
rect 283978 319932 284030 319938
rect 284082 319926 284156 319954
rect 283978 319874 284030 319880
rect 284128 319818 284156 319926
rect 284266 319920 284294 320076
rect 284358 319938 284386 320076
rect 283852 319688 283926 319716
rect 284036 319790 284156 319818
rect 284220 319892 284294 319920
rect 284346 319932 284398 319938
rect 283748 318368 283800 318374
rect 283748 318310 283800 318316
rect 283748 317824 283800 317830
rect 283748 317766 283800 317772
rect 283760 317626 283788 317766
rect 283748 317620 283800 317626
rect 283748 317562 283800 317568
rect 283656 317552 283708 317558
rect 283656 317494 283708 317500
rect 283484 315982 283604 316010
rect 283380 295996 283432 296002
rect 283380 295938 283432 295944
rect 283484 273970 283512 315982
rect 283564 315444 283616 315450
rect 283564 315386 283616 315392
rect 283472 273964 283524 273970
rect 283472 273906 283524 273912
rect 282828 235408 282880 235414
rect 282828 235350 282880 235356
rect 282552 231328 282604 231334
rect 282552 231270 282604 231276
rect 283012 227044 283064 227050
rect 283012 226986 283064 226992
rect 283024 226438 283052 226986
rect 283012 226432 283064 226438
rect 283012 226374 283064 226380
rect 282368 221808 282420 221814
rect 282368 221750 282420 221756
rect 282918 220280 282974 220289
rect 282918 220215 282920 220224
rect 282972 220215 282974 220224
rect 282920 220186 282972 220192
rect 283024 219434 283052 226374
rect 282932 219406 283052 219434
rect 282184 216504 282236 216510
rect 282184 216446 282236 216452
rect 282932 16574 282960 219406
rect 283576 219298 283604 315386
rect 283668 311250 283696 317494
rect 283852 316062 283880 319688
rect 284036 319297 284064 319790
rect 284022 319288 284078 319297
rect 284220 319274 284248 319892
rect 284346 319874 284398 319880
rect 284450 319818 284478 320076
rect 284022 319223 284078 319232
rect 284128 319246 284248 319274
rect 284312 319790 284478 319818
rect 284542 319818 284570 320076
rect 284634 320074 284662 320076
rect 284622 320068 284674 320074
rect 285540 320104 285596 320113
rect 284712 320039 284768 320048
rect 284622 320010 284674 320016
rect 284818 319938 284846 320076
rect 284910 319938 284938 320076
rect 284806 319932 284858 319938
rect 284806 319874 284858 319880
rect 284898 319932 284950 319938
rect 284898 319874 284950 319880
rect 285002 319818 285030 320076
rect 284542 319790 284662 319818
rect 284022 318336 284078 318345
rect 284022 318271 284078 318280
rect 283932 317620 283984 317626
rect 283932 317562 283984 317568
rect 283840 316056 283892 316062
rect 283840 315998 283892 316004
rect 283668 311222 283788 311250
rect 283654 309632 283710 309641
rect 283654 309567 283710 309576
rect 283564 219292 283616 219298
rect 283564 219234 283616 219240
rect 283668 219094 283696 309567
rect 283760 306374 283788 311222
rect 283760 306346 283880 306374
rect 283748 305720 283800 305726
rect 283748 305662 283800 305668
rect 283760 226438 283788 305662
rect 283852 294681 283880 306346
rect 283944 297809 283972 317562
rect 284036 312662 284064 318271
rect 284128 316130 284156 319246
rect 284206 319152 284262 319161
rect 284206 319087 284262 319096
rect 284220 318850 284248 319087
rect 284208 318844 284260 318850
rect 284208 318786 284260 318792
rect 284206 318200 284262 318209
rect 284206 318135 284262 318144
rect 284220 316577 284248 318135
rect 284312 317414 284340 319790
rect 284484 319728 284536 319734
rect 284484 319670 284536 319676
rect 284634 319682 284662 319790
rect 284760 319796 284812 319802
rect 284956 319790 285030 319818
rect 285094 319818 285122 320076
rect 285278 319954 285306 320076
rect 285232 319926 285306 319954
rect 285094 319790 285168 319818
rect 284812 319756 284892 319784
rect 284760 319738 284812 319744
rect 284312 317386 284432 317414
rect 284206 316568 284262 316577
rect 284206 316503 284262 316512
rect 284300 316260 284352 316266
rect 284300 316202 284352 316208
rect 284116 316124 284168 316130
rect 284116 316066 284168 316072
rect 284312 315314 284340 316202
rect 284404 315450 284432 317386
rect 284392 315444 284444 315450
rect 284392 315386 284444 315392
rect 284300 315308 284352 315314
rect 284300 315250 284352 315256
rect 284392 315308 284444 315314
rect 284392 315250 284444 315256
rect 284024 312656 284076 312662
rect 284024 312598 284076 312604
rect 284404 309942 284432 315250
rect 284392 309936 284444 309942
rect 284392 309878 284444 309884
rect 284208 307352 284260 307358
rect 284208 307294 284260 307300
rect 283930 297800 283986 297809
rect 283930 297735 283986 297744
rect 283838 294672 283894 294681
rect 283838 294607 283894 294616
rect 284220 231266 284248 307294
rect 284496 245002 284524 319670
rect 284634 319654 284708 319682
rect 284574 319288 284630 319297
rect 284574 319223 284630 319232
rect 284588 283626 284616 319223
rect 284680 317414 284708 319654
rect 284864 318374 284892 319756
rect 284852 318368 284904 318374
rect 284852 318310 284904 318316
rect 284956 318050 284984 319790
rect 285036 319728 285088 319734
rect 285036 319670 285088 319676
rect 285048 319297 285076 319670
rect 285034 319288 285090 319297
rect 285034 319223 285090 319232
rect 285036 318776 285088 318782
rect 285036 318718 285088 318724
rect 284864 318022 284984 318050
rect 284680 317386 284800 317414
rect 284772 316985 284800 317386
rect 284758 316976 284814 316985
rect 284758 316911 284814 316920
rect 284864 316266 284892 318022
rect 284942 317928 284998 317937
rect 284942 317863 284998 317872
rect 284852 316260 284904 316266
rect 284852 316202 284904 316208
rect 284760 316192 284812 316198
rect 284760 316134 284812 316140
rect 284668 316124 284720 316130
rect 284668 316066 284720 316072
rect 284680 311098 284708 316066
rect 284668 311092 284720 311098
rect 284668 311034 284720 311040
rect 284576 283620 284628 283626
rect 284576 283562 284628 283568
rect 284484 244996 284536 245002
rect 284484 244938 284536 244944
rect 284772 239057 284800 316134
rect 284852 316056 284904 316062
rect 284852 315998 284904 316004
rect 284864 241369 284892 315998
rect 284850 241360 284906 241369
rect 284850 241295 284906 241304
rect 284758 239048 284814 239057
rect 284758 238983 284814 238992
rect 284208 231260 284260 231266
rect 284208 231202 284260 231208
rect 284220 231146 284248 231202
rect 284220 231118 284432 231146
rect 283748 226432 283800 226438
rect 283748 226374 283800 226380
rect 283656 219088 283708 219094
rect 283656 219030 283708 219036
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284404 6914 284432 231118
rect 284956 220386 284984 317863
rect 285048 315314 285076 318718
rect 285140 318458 285168 319790
rect 285232 318782 285260 319926
rect 285370 319852 285398 320076
rect 285324 319824 285398 319852
rect 285220 318776 285272 318782
rect 285220 318718 285272 318724
rect 285140 318430 285260 318458
rect 285128 318368 285180 318374
rect 285128 318310 285180 318316
rect 285036 315308 285088 315314
rect 285036 315250 285088 315256
rect 285036 310004 285088 310010
rect 285036 309946 285088 309952
rect 284944 220380 284996 220386
rect 284944 220322 284996 220328
rect 285048 218657 285076 309946
rect 285140 307222 285168 318310
rect 285232 317665 285260 318430
rect 285218 317656 285274 317665
rect 285218 317591 285274 317600
rect 285324 316062 285352 319824
rect 285462 319784 285490 320076
rect 286092 320104 286148 320113
rect 285540 320039 285596 320048
rect 285646 319920 285674 320076
rect 285600 319892 285674 319920
rect 285600 319852 285628 319892
rect 285416 319756 285490 319784
rect 285554 319824 285628 319852
rect 285738 319852 285766 320076
rect 285738 319824 285812 319852
rect 285554 319784 285582 319824
rect 285554 319756 285628 319784
rect 285416 318646 285444 319756
rect 285494 319288 285550 319297
rect 285494 319223 285550 319232
rect 285404 318640 285456 318646
rect 285404 318582 285456 318588
rect 285508 316198 285536 319223
rect 285496 316192 285548 316198
rect 285496 316134 285548 316140
rect 285600 316130 285628 319756
rect 285784 317801 285812 319824
rect 285922 319818 285950 320076
rect 285876 319790 285950 319818
rect 286014 319818 286042 320076
rect 287656 320104 287712 320113
rect 286092 320039 286148 320048
rect 286198 319920 286226 320076
rect 286152 319892 286226 319920
rect 286014 319790 286088 319818
rect 285770 317792 285826 317801
rect 285770 317727 285826 317736
rect 285588 316124 285640 316130
rect 285588 316066 285640 316072
rect 285312 316056 285364 316062
rect 285312 315998 285364 316004
rect 285680 316056 285732 316062
rect 285680 315998 285732 316004
rect 285692 310350 285720 315998
rect 285680 310344 285732 310350
rect 285680 310286 285732 310292
rect 285678 309904 285734 309913
rect 285678 309839 285734 309848
rect 285692 309194 285720 309839
rect 285680 309188 285732 309194
rect 285680 309130 285732 309136
rect 285588 307420 285640 307426
rect 285588 307362 285640 307368
rect 285128 307216 285180 307222
rect 285128 307158 285180 307164
rect 285600 220182 285628 307362
rect 285876 307154 285904 319790
rect 285956 319728 286008 319734
rect 285956 319670 286008 319676
rect 285968 308446 285996 319670
rect 285956 308440 286008 308446
rect 285956 308382 286008 308388
rect 285864 307148 285916 307154
rect 285864 307090 285916 307096
rect 286060 282198 286088 319790
rect 286152 317529 286180 319892
rect 286290 319818 286318 320076
rect 286382 319870 286410 320076
rect 286566 319920 286594 320076
rect 286566 319892 286640 319920
rect 286244 319790 286318 319818
rect 286370 319864 286422 319870
rect 286370 319806 286422 319812
rect 286508 319796 286560 319802
rect 286244 318306 286272 319790
rect 286508 319738 286560 319744
rect 286324 318776 286376 318782
rect 286324 318718 286376 318724
rect 286232 318300 286284 318306
rect 286232 318242 286284 318248
rect 286232 318164 286284 318170
rect 286232 318106 286284 318112
rect 286138 317520 286194 317529
rect 286138 317455 286194 317464
rect 286244 296177 286272 318106
rect 286230 296168 286286 296177
rect 286230 296103 286286 296112
rect 286048 282192 286100 282198
rect 286048 282134 286100 282140
rect 286336 220454 286364 318718
rect 286416 315036 286468 315042
rect 286416 314978 286468 314984
rect 286324 220448 286376 220454
rect 286324 220390 286376 220396
rect 286428 220318 286456 314978
rect 286520 312526 286548 319738
rect 286612 317121 286640 319892
rect 286750 319852 286778 320076
rect 286704 319824 286778 319852
rect 286704 318850 286732 319824
rect 286842 319784 286870 320076
rect 286934 319920 286962 320076
rect 287026 320074 287054 320076
rect 287014 320068 287066 320074
rect 287014 320010 287066 320016
rect 286934 319892 287008 319920
rect 286796 319756 286870 319784
rect 286692 318844 286744 318850
rect 286692 318786 286744 318792
rect 286690 318744 286746 318753
rect 286690 318679 286746 318688
rect 286598 317112 286654 317121
rect 286598 317047 286654 317056
rect 286704 313886 286732 318679
rect 286796 318170 286824 319756
rect 286876 318844 286928 318850
rect 286876 318786 286928 318792
rect 286784 318164 286836 318170
rect 286784 318106 286836 318112
rect 286784 317892 286836 317898
rect 286784 317834 286836 317840
rect 286692 313880 286744 313886
rect 286692 313822 286744 313828
rect 286508 312520 286560 312526
rect 286508 312462 286560 312468
rect 286508 309936 286560 309942
rect 286508 309878 286560 309884
rect 286416 220312 286468 220318
rect 286416 220254 286468 220260
rect 285588 220176 285640 220182
rect 285588 220118 285640 220124
rect 285600 219434 285628 220118
rect 285600 219406 285720 219434
rect 285034 218648 285090 218657
rect 285034 218583 285090 218592
rect 285692 16574 285720 219406
rect 286520 218521 286548 309878
rect 286598 307184 286654 307193
rect 286598 307119 286654 307128
rect 286692 307148 286744 307154
rect 286612 224398 286640 307119
rect 286692 307090 286744 307096
rect 286704 225865 286732 307090
rect 286796 239562 286824 317834
rect 286888 316062 286916 318786
rect 286980 317665 287008 319892
rect 287118 319818 287146 320076
rect 287072 319790 287146 319818
rect 286966 317656 287022 317665
rect 286966 317591 287022 317600
rect 287072 317529 287100 319790
rect 287210 319716 287238 320076
rect 287302 319818 287330 320076
rect 287486 319938 287514 320076
rect 287578 319954 287606 320076
rect 288392 320104 288448 320113
rect 287656 320039 287712 320048
rect 287474 319932 287526 319938
rect 287578 319926 287652 319954
rect 287474 319874 287526 319880
rect 287302 319790 287422 319818
rect 287394 319784 287422 319790
rect 287520 319796 287572 319802
rect 287394 319756 287468 319784
rect 287164 319688 287238 319716
rect 287164 318209 287192 319688
rect 287244 318232 287296 318238
rect 287150 318200 287206 318209
rect 287244 318174 287296 318180
rect 287150 318135 287206 318144
rect 287150 318064 287206 318073
rect 287256 318034 287284 318174
rect 287150 317999 287206 318008
rect 287244 318028 287296 318034
rect 287058 317520 287114 317529
rect 287058 317455 287114 317464
rect 286876 316056 286928 316062
rect 286876 315998 286928 316004
rect 287164 315314 287192 317999
rect 287244 317970 287296 317976
rect 287336 316124 287388 316130
rect 287336 316066 287388 316072
rect 287244 316056 287296 316062
rect 287244 315998 287296 316004
rect 287152 315308 287204 315314
rect 287152 315250 287204 315256
rect 286876 314220 286928 314226
rect 286876 314162 286928 314168
rect 286784 239556 286836 239562
rect 286784 239498 286836 239504
rect 286888 235618 286916 314162
rect 287150 309360 287206 309369
rect 287150 309295 287206 309304
rect 287164 309262 287192 309295
rect 287152 309256 287204 309262
rect 287152 309198 287204 309204
rect 287256 291961 287284 315998
rect 287348 296041 287376 316066
rect 287440 298761 287468 319756
rect 287520 319738 287572 319744
rect 287532 318782 287560 319738
rect 287520 318776 287572 318782
rect 287520 318718 287572 318724
rect 287624 315602 287652 319926
rect 287762 319920 287790 320076
rect 287716 319892 287790 319920
rect 287716 317529 287744 319892
rect 287854 319818 287882 320076
rect 287808 319790 287882 319818
rect 287808 318753 287836 319790
rect 287946 319716 287974 320076
rect 288222 319920 288250 320076
rect 287900 319688 287974 319716
rect 288176 319892 288250 319920
rect 287794 318744 287850 318753
rect 287794 318679 287850 318688
rect 287796 318640 287848 318646
rect 287796 318582 287848 318588
rect 287808 318102 287836 318582
rect 287796 318096 287848 318102
rect 287796 318038 287848 318044
rect 287794 317792 287850 317801
rect 287794 317727 287850 317736
rect 287702 317520 287758 317529
rect 287702 317455 287758 317464
rect 287624 315574 287744 315602
rect 287612 315444 287664 315450
rect 287612 315386 287664 315392
rect 287426 298752 287482 298761
rect 287426 298687 287482 298696
rect 287334 296032 287390 296041
rect 287334 295967 287390 295976
rect 287242 291952 287298 291961
rect 287242 291887 287298 291896
rect 286876 235612 286928 235618
rect 286876 235554 286928 235560
rect 286690 225856 286746 225865
rect 286690 225791 286746 225800
rect 286600 224392 286652 224398
rect 286600 224334 286652 224340
rect 287426 223544 287482 223553
rect 287426 223479 287482 223488
rect 287440 222902 287468 223479
rect 287624 223242 287652 315386
rect 287716 315382 287744 315574
rect 287704 315376 287756 315382
rect 287704 315318 287756 315324
rect 287808 311894 287836 317727
rect 287900 316130 287928 319688
rect 288070 319288 288126 319297
rect 288070 319223 288126 319232
rect 287978 318744 288034 318753
rect 287978 318679 288034 318688
rect 287888 316124 287940 316130
rect 287888 316066 287940 316072
rect 287992 315466 288020 318679
rect 287900 315438 288020 315466
rect 287900 315042 287928 315438
rect 287980 315376 288032 315382
rect 287980 315318 288032 315324
rect 287888 315036 287940 315042
rect 287888 314978 287940 314984
rect 287716 311866 287836 311894
rect 287612 223236 287664 223242
rect 287612 223178 287664 223184
rect 287428 222896 287480 222902
rect 287428 222838 287480 222844
rect 287716 219230 287744 311866
rect 287888 307624 287940 307630
rect 287888 307566 287940 307572
rect 287796 307012 287848 307018
rect 287796 306954 287848 306960
rect 287704 219224 287756 219230
rect 287704 219166 287756 219172
rect 287808 218929 287836 306954
rect 287900 221746 287928 307566
rect 287992 290737 288020 315318
rect 288084 302841 288112 319223
rect 288176 316062 288204 319892
rect 288314 319852 288342 320076
rect 288852 320104 288908 320113
rect 288392 320039 288448 320048
rect 288498 319954 288526 320076
rect 288268 319824 288342 319852
rect 288452 319926 288526 319954
rect 288164 316056 288216 316062
rect 288164 315998 288216 316004
rect 288268 315450 288296 319824
rect 288346 318744 288402 318753
rect 288346 318679 288402 318688
rect 288256 315444 288308 315450
rect 288256 315386 288308 315392
rect 288360 315382 288388 318679
rect 288348 315376 288400 315382
rect 288348 315318 288400 315324
rect 288452 315314 288480 319926
rect 288590 319852 288618 320076
rect 288544 319824 288618 319852
rect 288544 317529 288572 319824
rect 288682 319784 288710 320076
rect 288774 319954 288802 320076
rect 289404 320104 289460 320113
rect 288852 320039 288908 320048
rect 288958 319954 288986 320076
rect 288774 319926 288848 319954
rect 288636 319756 288710 319784
rect 288636 318209 288664 319756
rect 288716 318844 288768 318850
rect 288716 318786 288768 318792
rect 288622 318200 288678 318209
rect 288622 318135 288678 318144
rect 288530 317520 288586 317529
rect 288530 317455 288586 317464
rect 288532 316124 288584 316130
rect 288532 316066 288584 316072
rect 288256 315308 288308 315314
rect 288256 315250 288308 315256
rect 288440 315308 288492 315314
rect 288440 315250 288492 315256
rect 288268 311642 288296 315250
rect 288438 312080 288494 312089
rect 288438 312015 288440 312024
rect 288492 312015 288494 312024
rect 288440 311986 288492 311992
rect 288256 311636 288308 311642
rect 288256 311578 288308 311584
rect 288348 307488 288400 307494
rect 288348 307430 288400 307436
rect 288070 302832 288126 302841
rect 288070 302767 288126 302776
rect 287978 290728 288034 290737
rect 287978 290663 288034 290672
rect 287888 221740 287940 221746
rect 287888 221682 287940 221688
rect 287794 218920 287850 218929
rect 288360 218890 288388 307430
rect 288544 247761 288572 316066
rect 288624 316056 288676 316062
rect 288624 315998 288676 316004
rect 288636 310282 288664 315998
rect 288624 310276 288676 310282
rect 288624 310218 288676 310224
rect 288728 307562 288756 318786
rect 288820 318238 288848 319926
rect 288912 319926 288986 319954
rect 288912 319784 288940 319926
rect 288912 319756 289032 319784
rect 288898 318744 288954 318753
rect 288898 318679 288954 318688
rect 288808 318232 288860 318238
rect 288808 318174 288860 318180
rect 288808 318028 288860 318034
rect 288808 317970 288860 317976
rect 288820 308514 288848 317970
rect 288912 315110 288940 318679
rect 288900 315104 288952 315110
rect 288900 315046 288952 315052
rect 288808 308508 288860 308514
rect 288808 308450 288860 308456
rect 288716 307556 288768 307562
rect 288716 307498 288768 307504
rect 288530 247752 288586 247761
rect 288530 247687 288586 247696
rect 289004 238921 289032 319756
rect 289142 319716 289170 320076
rect 289234 319818 289262 320076
rect 289326 319920 289354 320076
rect 289864 320104 289920 320113
rect 289404 320039 289460 320048
rect 289510 319938 289538 320076
rect 289498 319932 289550 319938
rect 289326 319892 289400 319920
rect 289234 319790 289308 319818
rect 289096 319688 289170 319716
rect 289096 318034 289124 319688
rect 289280 318322 289308 319790
rect 289188 318294 289308 318322
rect 289084 318028 289136 318034
rect 289084 317970 289136 317976
rect 289082 317656 289138 317665
rect 289082 317591 289138 317600
rect 288990 238912 289046 238921
rect 288990 238847 289046 238856
rect 289096 220153 289124 317591
rect 289188 316062 289216 318294
rect 289268 318232 289320 318238
rect 289268 318174 289320 318180
rect 289176 316056 289228 316062
rect 289176 315998 289228 316004
rect 289280 311894 289308 318174
rect 289372 316130 289400 319892
rect 289498 319874 289550 319880
rect 289602 319818 289630 320076
rect 289786 319920 289814 320076
rect 290416 320104 290472 320113
rect 289864 320039 289920 320048
rect 289970 319920 289998 320076
rect 290062 319938 290090 320076
rect 290246 319954 290274 320076
rect 290876 320104 290932 320113
rect 290416 320039 290472 320048
rect 289740 319892 289814 319920
rect 289924 319892 289998 319920
rect 290050 319932 290102 319938
rect 289740 319852 289768 319892
rect 289452 319796 289504 319802
rect 289452 319738 289504 319744
rect 289556 319790 289630 319818
rect 289694 319824 289768 319852
rect 289464 318782 289492 319738
rect 289452 318776 289504 318782
rect 289452 318718 289504 318724
rect 289556 318481 289584 319790
rect 289694 319784 289722 319824
rect 289694 319756 289768 319784
rect 289740 318850 289768 319756
rect 289924 319410 289952 319892
rect 290050 319874 290102 319880
rect 290154 319926 290274 319954
rect 290154 319818 290182 319926
rect 290522 319920 290550 320076
rect 290476 319892 290550 319920
rect 290004 319796 290056 319802
rect 290154 319790 290228 319818
rect 290004 319738 290056 319744
rect 289832 319382 289952 319410
rect 289728 318844 289780 318850
rect 289728 318786 289780 318792
rect 289636 318776 289688 318782
rect 289636 318718 289688 318724
rect 289542 318472 289598 318481
rect 289452 318436 289504 318442
rect 289542 318407 289598 318416
rect 289452 318378 289504 318384
rect 289360 316124 289412 316130
rect 289360 316066 289412 316072
rect 289280 311866 289400 311894
rect 289176 310480 289228 310486
rect 289176 310422 289228 310428
rect 289188 227089 289216 310422
rect 289268 310412 289320 310418
rect 289268 310354 289320 310360
rect 289280 230110 289308 310354
rect 289372 308689 289400 311866
rect 289464 311166 289492 318378
rect 289542 317928 289598 317937
rect 289542 317863 289598 317872
rect 289556 317558 289584 317863
rect 289544 317552 289596 317558
rect 289544 317494 289596 317500
rect 289544 315308 289596 315314
rect 289544 315250 289596 315256
rect 289452 311160 289504 311166
rect 289452 311102 289504 311108
rect 289358 308680 289414 308689
rect 289358 308615 289414 308624
rect 289452 308508 289504 308514
rect 289452 308450 289504 308456
rect 289360 307216 289412 307222
rect 289360 307158 289412 307164
rect 289268 230104 289320 230110
rect 289268 230046 289320 230052
rect 289372 229090 289400 307158
rect 289464 238513 289492 308450
rect 289556 304201 289584 315250
rect 289648 306406 289676 318718
rect 289832 316713 289860 319382
rect 289910 319288 289966 319297
rect 289910 319223 289966 319232
rect 289818 316704 289874 316713
rect 289818 316639 289874 316648
rect 289924 316062 289952 319223
rect 289912 316056 289964 316062
rect 289912 315998 289964 316004
rect 290016 315450 290044 319738
rect 290094 318744 290150 318753
rect 290094 318679 290150 318688
rect 290004 315444 290056 315450
rect 290004 315386 290056 315392
rect 290108 307329 290136 318679
rect 290200 317801 290228 319790
rect 290370 319288 290426 319297
rect 290370 319223 290426 319232
rect 290186 317792 290242 317801
rect 290186 317727 290242 317736
rect 290188 316124 290240 316130
rect 290188 316066 290240 316072
rect 290200 309806 290228 316066
rect 290384 315602 290412 319223
rect 290476 316130 290504 319892
rect 290614 319852 290642 320076
rect 290568 319824 290642 319852
rect 290464 316124 290516 316130
rect 290464 316066 290516 316072
rect 290384 315574 290504 315602
rect 290372 315444 290424 315450
rect 290372 315386 290424 315392
rect 290280 315376 290332 315382
rect 290280 315318 290332 315324
rect 290188 309800 290240 309806
rect 290188 309742 290240 309748
rect 290094 307320 290150 307329
rect 290094 307255 290150 307264
rect 289636 306400 289688 306406
rect 289636 306342 289688 306348
rect 289542 304192 289598 304201
rect 289542 304127 289598 304136
rect 289450 238504 289506 238513
rect 289450 238439 289506 238448
rect 289360 229084 289412 229090
rect 289360 229026 289412 229032
rect 289174 227080 289230 227089
rect 289174 227015 289230 227024
rect 290292 220590 290320 315318
rect 290384 307601 290412 315386
rect 290476 314566 290504 315574
rect 290568 314634 290596 319824
rect 290706 319784 290734 320076
rect 290660 319756 290734 319784
rect 290798 319784 290826 320076
rect 291520 320104 291576 320113
rect 290876 320039 290932 320048
rect 291166 319784 291194 320076
rect 290798 319756 290964 319784
rect 290660 317626 290688 319756
rect 290830 319288 290886 319297
rect 290830 319223 290886 319232
rect 290740 318232 290792 318238
rect 290740 318174 290792 318180
rect 290648 317620 290700 317626
rect 290648 317562 290700 317568
rect 290752 316146 290780 318174
rect 290660 316118 290780 316146
rect 290660 315994 290688 316118
rect 290740 316056 290792 316062
rect 290740 315998 290792 316004
rect 290648 315988 290700 315994
rect 290648 315930 290700 315936
rect 290556 314628 290608 314634
rect 290556 314570 290608 314576
rect 290464 314560 290516 314566
rect 290464 314502 290516 314508
rect 290648 313676 290700 313682
rect 290648 313618 290700 313624
rect 290370 307592 290426 307601
rect 290370 307527 290426 307536
rect 290556 307556 290608 307562
rect 290556 307498 290608 307504
rect 290464 307284 290516 307290
rect 290464 307226 290516 307232
rect 290476 221513 290504 307226
rect 290568 224534 290596 307498
rect 290660 237590 290688 313618
rect 290752 275330 290780 315998
rect 290740 275324 290792 275330
rect 290740 275266 290792 275272
rect 290844 260166 290872 319223
rect 290936 318850 290964 319756
rect 291028 319756 291194 319784
rect 290924 318844 290976 318850
rect 290924 318786 290976 318792
rect 290922 318744 290978 318753
rect 290922 318679 290978 318688
rect 290936 284986 290964 318679
rect 291028 315761 291056 319756
rect 291258 319716 291286 320076
rect 291442 319784 291470 320076
rect 291704 320104 291760 320113
rect 291520 320039 291576 320048
rect 291626 319938 291654 320076
rect 292348 320104 292404 320113
rect 291704 320039 291760 320048
rect 291810 319954 291838 320076
rect 291614 319932 291666 319938
rect 291614 319874 291666 319880
rect 291764 319926 291838 319954
rect 291442 319756 291516 319784
rect 291212 319688 291286 319716
rect 291212 319410 291240 319688
rect 291212 319382 291332 319410
rect 291198 319288 291254 319297
rect 291198 319223 291254 319232
rect 291108 318844 291160 318850
rect 291108 318786 291160 318792
rect 291014 315752 291070 315761
rect 291014 315687 291070 315696
rect 291120 309874 291148 318786
rect 291212 313682 291240 319223
rect 291304 317529 291332 319382
rect 291290 317520 291346 317529
rect 291290 317455 291346 317464
rect 291488 317414 291516 319756
rect 291568 319728 291620 319734
rect 291568 319670 291620 319676
rect 291580 317529 291608 319670
rect 291764 319648 291792 319926
rect 291902 319852 291930 320076
rect 291672 319620 291792 319648
rect 291856 319824 291930 319852
rect 291566 317520 291622 317529
rect 291566 317455 291622 317464
rect 291396 317386 291516 317414
rect 291200 313676 291252 313682
rect 291200 313618 291252 313624
rect 291108 309868 291160 309874
rect 291108 309810 291160 309816
rect 290924 284980 290976 284986
rect 290924 284922 290976 284928
rect 290832 260160 290884 260166
rect 290832 260102 290884 260108
rect 291396 238785 291424 317386
rect 291476 316056 291528 316062
rect 291672 316010 291700 319620
rect 291856 317414 291884 319824
rect 291994 319784 292022 320076
rect 291948 319756 292022 319784
rect 291948 318889 291976 319756
rect 292086 319716 292114 320076
rect 292178 319852 292206 320076
rect 292270 319954 292298 320076
rect 293176 320104 293232 320113
rect 292348 320039 292404 320048
rect 292270 319926 292436 319954
rect 292178 319824 292344 319852
rect 292040 319688 292114 319716
rect 291934 318880 291990 318889
rect 291934 318815 291990 318824
rect 291936 318368 291988 318374
rect 291936 318310 291988 318316
rect 291476 315998 291528 316004
rect 291488 251870 291516 315998
rect 291580 315982 291700 316010
rect 291764 317386 291884 317414
rect 291580 264246 291608 315982
rect 291660 313948 291712 313954
rect 291660 313890 291712 313896
rect 291568 264240 291620 264246
rect 291568 264182 291620 264188
rect 291476 251864 291528 251870
rect 291476 251806 291528 251812
rect 291382 238776 291438 238785
rect 291382 238711 291438 238720
rect 290648 237584 290700 237590
rect 290648 237526 290700 237532
rect 291672 230246 291700 313890
rect 291764 239834 291792 317386
rect 291844 315308 291896 315314
rect 291844 315250 291896 315256
rect 291752 239828 291804 239834
rect 291752 239770 291804 239776
rect 291660 230240 291712 230246
rect 291660 230182 291712 230188
rect 291856 230042 291884 315250
rect 291948 314090 291976 318310
rect 292040 316062 292068 319688
rect 292120 319116 292172 319122
rect 292120 319058 292172 319064
rect 292132 318850 292160 319058
rect 292210 318880 292266 318889
rect 292120 318844 292172 318850
rect 292210 318815 292266 318824
rect 292120 318786 292172 318792
rect 292120 318300 292172 318306
rect 292120 318242 292172 318248
rect 292028 316056 292080 316062
rect 292028 315998 292080 316004
rect 291936 314084 291988 314090
rect 291936 314026 291988 314032
rect 291936 311908 291988 311914
rect 292132 311894 292160 318242
rect 292224 314158 292252 318815
rect 292316 317830 292344 319824
rect 292304 317824 292356 317830
rect 292304 317766 292356 317772
rect 292408 316538 292436 319926
rect 292546 319818 292574 320076
rect 292500 319790 292574 319818
rect 292396 316532 292448 316538
rect 292396 316474 292448 316480
rect 292394 315752 292450 315761
rect 292394 315687 292396 315696
rect 292448 315687 292450 315696
rect 292396 315658 292448 315664
rect 292304 315648 292356 315654
rect 292304 315590 292356 315596
rect 292316 315382 292344 315590
rect 292304 315376 292356 315382
rect 292304 315318 292356 315324
rect 292212 314152 292264 314158
rect 292212 314094 292264 314100
rect 292500 313954 292528 319790
rect 292638 319784 292666 320076
rect 292730 319938 292758 320076
rect 292718 319932 292770 319938
rect 292718 319874 292770 319880
rect 292822 319784 292850 320076
rect 292638 319756 292712 319784
rect 292684 317529 292712 319756
rect 292776 319756 292850 319784
rect 292670 317520 292726 317529
rect 292670 317455 292726 317464
rect 292776 315976 292804 319756
rect 292914 319716 292942 320076
rect 293006 319784 293034 320076
rect 293098 319852 293126 320076
rect 293728 320104 293784 320113
rect 293176 320039 293232 320048
rect 293282 319954 293310 320076
rect 293236 319926 293310 319954
rect 293098 319824 293172 319852
rect 293006 319756 293080 319784
rect 292868 319688 292942 319716
rect 292868 317665 292896 319688
rect 292948 318844 293000 318850
rect 292948 318786 293000 318792
rect 292854 317656 292910 317665
rect 292854 317591 292910 317600
rect 292684 315948 292804 315976
rect 292856 315988 292908 315994
rect 292580 315784 292632 315790
rect 292580 315726 292632 315732
rect 292592 315110 292620 315726
rect 292580 315104 292632 315110
rect 292580 315046 292632 315052
rect 292488 313948 292540 313954
rect 292488 313890 292540 313896
rect 292578 312080 292634 312089
rect 292578 312015 292634 312024
rect 292592 311982 292620 312015
rect 292580 311976 292632 311982
rect 292580 311918 292632 311924
rect 291936 311850 291988 311856
rect 292040 311866 292160 311894
rect 291844 230036 291896 230042
rect 291844 229978 291896 229984
rect 290556 224528 290608 224534
rect 290556 224470 290608 224476
rect 290462 221504 290518 221513
rect 290462 221439 290518 221448
rect 290280 220584 290332 220590
rect 290280 220526 290332 220532
rect 289082 220144 289138 220153
rect 289082 220079 289138 220088
rect 287794 218855 287850 218864
rect 288348 218884 288400 218890
rect 288348 218826 288400 218832
rect 286506 218512 286562 218521
rect 286506 218447 286562 218456
rect 288360 218074 288388 218826
rect 288348 218068 288400 218074
rect 288348 218010 288400 218016
rect 289084 218068 289136 218074
rect 289084 218010 289136 218016
rect 285692 16546 286640 16574
rect 284312 6886 284432 6914
rect 284312 480 284340 6886
rect 285404 3664 285456 3670
rect 285404 3606 285456 3612
rect 285416 480 285444 3606
rect 286612 480 286640 16546
rect 288992 4004 289044 4010
rect 288992 3946 289044 3952
rect 287796 3460 287848 3466
rect 287796 3402 287848 3408
rect 287808 480 287836 3402
rect 289004 480 289032 3946
rect 289096 3534 289124 218010
rect 289174 211848 289230 211857
rect 289174 211783 289230 211792
rect 289084 3528 289136 3534
rect 289084 3470 289136 3476
rect 289188 3466 289216 211783
rect 291856 3670 291884 229978
rect 291948 222737 291976 311850
rect 292040 232966 292068 311866
rect 292028 232960 292080 232966
rect 292028 232902 292080 232908
rect 292684 230382 292712 315948
rect 292856 315930 292908 315936
rect 292764 315852 292816 315858
rect 292764 315794 292816 315800
rect 292776 234530 292804 315794
rect 292764 234524 292816 234530
rect 292764 234466 292816 234472
rect 292868 234326 292896 315930
rect 292960 240038 292988 318786
rect 293052 318782 293080 319756
rect 293040 318776 293092 318782
rect 293040 318718 293092 318724
rect 293038 315752 293094 315761
rect 293038 315687 293040 315696
rect 293092 315687 293094 315696
rect 293040 315658 293092 315664
rect 292948 240032 293000 240038
rect 292948 239974 293000 239980
rect 292856 234320 292908 234326
rect 292856 234262 292908 234268
rect 292672 230376 292724 230382
rect 292672 230318 292724 230324
rect 293144 227458 293172 319824
rect 293236 319433 293264 319926
rect 293374 319784 293402 320076
rect 293650 319852 293678 320076
rect 294280 320104 294336 320113
rect 293728 320039 293784 320048
rect 293834 319938 293862 320076
rect 293822 319932 293874 319938
rect 293822 319874 293874 319880
rect 293926 319870 293954 320076
rect 293914 319864 293966 319870
rect 293650 319824 293724 319852
rect 293374 319756 293448 319784
rect 293222 319424 293278 319433
rect 293420 319410 293448 319756
rect 293420 319382 293540 319410
rect 293222 319359 293278 319368
rect 293222 318880 293278 318889
rect 293222 318815 293278 318824
rect 293236 315858 293264 318815
rect 293316 318776 293368 318782
rect 293316 318718 293368 318724
rect 293224 315852 293276 315858
rect 293224 315794 293276 315800
rect 293224 313268 293276 313274
rect 293224 313210 293276 313216
rect 293236 234122 293264 313210
rect 293328 310486 293356 318718
rect 293512 318288 293540 319382
rect 293696 318782 293724 319824
rect 293914 319806 293966 319812
rect 293776 319796 293828 319802
rect 294018 319784 294046 320076
rect 295016 320104 295072 320113
rect 294280 320039 294336 320048
rect 294386 319954 294414 320076
rect 294248 319926 294414 319954
rect 294018 319756 294092 319784
rect 293776 319738 293828 319744
rect 293684 318776 293736 318782
rect 293684 318718 293736 318724
rect 293590 318472 293646 318481
rect 293590 318407 293646 318416
rect 293420 318260 293540 318288
rect 293420 317898 293448 318260
rect 293498 318200 293554 318209
rect 293498 318135 293554 318144
rect 293408 317892 293460 317898
rect 293408 317834 293460 317840
rect 293408 317620 293460 317626
rect 293408 317562 293460 317568
rect 293316 310480 293368 310486
rect 293316 310422 293368 310428
rect 293420 307562 293448 317562
rect 293512 311001 293540 318135
rect 293604 311914 293632 318407
rect 293788 315994 293816 319738
rect 293868 319660 293920 319666
rect 293868 319602 293920 319608
rect 293960 319660 294012 319666
rect 293960 319602 294012 319608
rect 293880 318850 293908 319602
rect 293868 318844 293920 318850
rect 293868 318786 293920 318792
rect 293868 317892 293920 317898
rect 293868 317834 293920 317840
rect 293880 316742 293908 317834
rect 293868 316736 293920 316742
rect 293868 316678 293920 316684
rect 293972 316606 294000 319602
rect 294064 318714 294092 319756
rect 294248 318968 294276 319926
rect 294328 319864 294380 319870
rect 294328 319806 294380 319812
rect 294156 318940 294276 318968
rect 294052 318708 294104 318714
rect 294052 318650 294104 318656
rect 294052 318572 294104 318578
rect 294052 318514 294104 318520
rect 294064 318102 294092 318514
rect 294052 318096 294104 318102
rect 294052 318038 294104 318044
rect 293960 316600 294012 316606
rect 293960 316542 294012 316548
rect 293776 315988 293828 315994
rect 293776 315930 293828 315936
rect 294052 315784 294104 315790
rect 294052 315726 294104 315732
rect 294064 315586 294092 315726
rect 293960 315580 294012 315586
rect 293960 315522 294012 315528
rect 294052 315580 294104 315586
rect 294052 315522 294104 315528
rect 293972 315450 294000 315522
rect 293960 315444 294012 315450
rect 293960 315386 294012 315392
rect 293592 311908 293644 311914
rect 293592 311850 293644 311856
rect 293498 310992 293554 311001
rect 293498 310927 293554 310936
rect 293408 307556 293460 307562
rect 293408 307498 293460 307504
rect 294156 234598 294184 318940
rect 294234 318880 294290 318889
rect 294234 318815 294290 318824
rect 294248 316062 294276 318815
rect 294340 316470 294368 319806
rect 294478 319784 294506 320076
rect 294570 319938 294598 320076
rect 294558 319932 294610 319938
rect 294558 319874 294610 319880
rect 294662 319784 294690 320076
rect 294432 319756 294506 319784
rect 294616 319756 294690 319784
rect 294432 318374 294460 319756
rect 294616 319716 294644 319756
rect 294754 319716 294782 320076
rect 294524 319688 294644 319716
rect 294708 319688 294782 319716
rect 294420 318368 294472 318374
rect 294420 318310 294472 318316
rect 294328 316464 294380 316470
rect 294328 316406 294380 316412
rect 294524 316146 294552 319688
rect 294602 319424 294658 319433
rect 294602 319359 294658 319368
rect 294616 319054 294644 319359
rect 294604 319048 294656 319054
rect 294604 318990 294656 318996
rect 294602 318880 294658 318889
rect 294602 318815 294658 318824
rect 294616 316810 294644 318815
rect 294604 316804 294656 316810
rect 294604 316746 294656 316752
rect 294340 316118 294552 316146
rect 294236 316056 294288 316062
rect 294236 315998 294288 316004
rect 294340 315874 294368 316118
rect 294512 316056 294564 316062
rect 294512 315998 294564 316004
rect 294604 316056 294656 316062
rect 294604 315998 294656 316004
rect 294248 315846 294368 315874
rect 294420 315852 294472 315858
rect 294248 239222 294276 315846
rect 294420 315794 294472 315800
rect 294328 315784 294380 315790
rect 294328 315726 294380 315732
rect 294236 239216 294288 239222
rect 294236 239158 294288 239164
rect 294144 234592 294196 234598
rect 294144 234534 294196 234540
rect 293224 234116 293276 234122
rect 293224 234058 293276 234064
rect 293132 227452 293184 227458
rect 293132 227394 293184 227400
rect 294340 224777 294368 315726
rect 294432 307018 294460 315794
rect 294420 307012 294472 307018
rect 294420 306954 294472 306960
rect 294524 233238 294552 315998
rect 294616 311894 294644 315998
rect 294708 315790 294736 319688
rect 294846 319648 294874 320076
rect 294938 319716 294966 320076
rect 295568 320104 295624 320113
rect 295016 320039 295072 320048
rect 295122 319920 295150 320076
rect 295214 319938 295242 320076
rect 295306 319938 295334 320076
rect 295076 319892 295150 319920
rect 295202 319932 295254 319938
rect 294938 319688 295012 319716
rect 294846 319620 294920 319648
rect 294788 318708 294840 318714
rect 294788 318650 294840 318656
rect 294800 317937 294828 318650
rect 294786 317928 294842 317937
rect 294786 317863 294842 317872
rect 294788 317824 294840 317830
rect 294788 317766 294840 317772
rect 294696 315784 294748 315790
rect 294696 315726 294748 315732
rect 294696 315648 294748 315654
rect 294696 315590 294748 315596
rect 294708 315382 294736 315590
rect 294696 315376 294748 315382
rect 294696 315318 294748 315324
rect 294616 311866 294736 311894
rect 294604 311160 294656 311166
rect 294604 311102 294656 311108
rect 294616 235754 294644 311102
rect 294604 235748 294656 235754
rect 294604 235690 294656 235696
rect 294708 235278 294736 311866
rect 294800 311166 294828 317766
rect 294892 315858 294920 319620
rect 294984 318646 295012 319688
rect 294972 318640 295024 318646
rect 294972 318582 295024 318588
rect 295076 317626 295104 319892
rect 295202 319874 295254 319880
rect 295294 319932 295346 319938
rect 295294 319874 295346 319880
rect 295490 319852 295518 320076
rect 295936 320104 295992 320113
rect 295568 320039 295624 320048
rect 295398 319824 295518 319852
rect 295156 319728 295208 319734
rect 295398 319716 295426 319824
rect 295674 319784 295702 320076
rect 295766 319938 295794 320076
rect 295754 319932 295806 319938
rect 295754 319874 295806 319880
rect 295858 319784 295886 320076
rect 296212 320104 296268 320113
rect 295936 320039 295992 320048
rect 296042 319784 296070 320076
rect 295674 319756 295748 319784
rect 295524 319728 295576 319734
rect 295398 319688 295472 319716
rect 295156 319670 295208 319676
rect 295168 318578 295196 319670
rect 295340 319456 295392 319462
rect 295338 319424 295340 319433
rect 295392 319424 295394 319433
rect 295338 319359 295394 319368
rect 295156 318572 295208 318578
rect 295156 318514 295208 318520
rect 295156 318436 295208 318442
rect 295156 318378 295208 318384
rect 295064 317620 295116 317626
rect 295064 317562 295116 317568
rect 294970 317384 295026 317393
rect 294970 317319 295026 317328
rect 294880 315852 294932 315858
rect 294880 315794 294932 315800
rect 294984 311894 295012 317319
rect 295168 315178 295196 318378
rect 295340 318028 295392 318034
rect 295340 317970 295392 317976
rect 295352 317694 295380 317970
rect 295444 317966 295472 319688
rect 295524 319670 295576 319676
rect 295536 318918 295564 319670
rect 295720 319462 295748 319756
rect 295812 319756 295886 319784
rect 295996 319756 296070 319784
rect 295708 319456 295760 319462
rect 295708 319398 295760 319404
rect 295708 319048 295760 319054
rect 295708 318990 295760 318996
rect 295524 318912 295576 318918
rect 295524 318854 295576 318860
rect 295616 318572 295668 318578
rect 295616 318514 295668 318520
rect 295432 317960 295484 317966
rect 295432 317902 295484 317908
rect 295340 317688 295392 317694
rect 295340 317630 295392 317636
rect 295340 317484 295392 317490
rect 295340 317426 295392 317432
rect 295248 316804 295300 316810
rect 295248 316746 295300 316752
rect 295156 315172 295208 315178
rect 295156 315114 295208 315120
rect 295260 314498 295288 316746
rect 295248 314492 295300 314498
rect 295248 314434 295300 314440
rect 294892 311866 295012 311894
rect 294788 311160 294840 311166
rect 294788 311102 294840 311108
rect 294892 307086 294920 311866
rect 295352 310418 295380 317426
rect 295628 316130 295656 318514
rect 295616 316124 295668 316130
rect 295616 316066 295668 316072
rect 295340 310412 295392 310418
rect 295340 310354 295392 310360
rect 294880 307080 294932 307086
rect 294880 307022 294932 307028
rect 294696 235272 294748 235278
rect 294696 235214 294748 235220
rect 294512 233232 294564 233238
rect 294512 233174 294564 233180
rect 294326 224768 294382 224777
rect 294326 224703 294382 224712
rect 291934 222728 291990 222737
rect 291934 222663 291990 222672
rect 295720 222018 295748 318990
rect 295812 317150 295840 319756
rect 295892 318708 295944 318714
rect 295892 318650 295944 318656
rect 295904 317558 295932 318650
rect 295996 318170 296024 319756
rect 296134 319682 296162 320076
rect 297316 320104 297372 320113
rect 296212 320039 296268 320048
rect 296318 319938 296346 320076
rect 296306 319932 296358 319938
rect 296306 319874 296358 319880
rect 296410 319784 296438 320076
rect 296364 319756 296438 319784
rect 296134 319654 296208 319682
rect 296076 319456 296128 319462
rect 296076 319398 296128 319404
rect 295984 318164 296036 318170
rect 295984 318106 296036 318112
rect 296088 318050 296116 319398
rect 295996 318022 296116 318050
rect 295892 317552 295944 317558
rect 295892 317494 295944 317500
rect 295996 317234 296024 318022
rect 296076 317620 296128 317626
rect 296076 317562 296128 317568
rect 295904 317206 296024 317234
rect 295800 317144 295852 317150
rect 295800 317086 295852 317092
rect 295904 312798 295932 317206
rect 295984 317144 296036 317150
rect 295984 317086 296036 317092
rect 295892 312792 295944 312798
rect 295892 312734 295944 312740
rect 295996 232898 296024 317086
rect 295984 232892 296036 232898
rect 295984 232834 296036 232840
rect 295708 222012 295760 222018
rect 295708 221954 295760 221960
rect 292580 209160 292632 209166
rect 292580 209102 292632 209108
rect 292592 208321 292620 209102
rect 292578 208312 292634 208321
rect 292578 208247 292634 208256
rect 292592 200114 292620 208247
rect 292592 200086 292712 200114
rect 292684 16574 292712 200086
rect 293958 166288 294014 166297
rect 293958 166223 294014 166232
rect 293972 16574 294000 166223
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 291844 3664 291896 3670
rect 291844 3606 291896 3612
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 289176 3460 289228 3466
rect 289176 3402 289228 3408
rect 290200 480 290228 3470
rect 291384 3460 291436 3466
rect 291384 3402 291436 3408
rect 291396 480 291424 3402
rect 292580 3392 292632 3398
rect 292580 3334 292632 3340
rect 292592 480 292620 3334
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 295996 3466 296024 232834
rect 296088 221882 296116 317562
rect 296180 317529 296208 319654
rect 296260 317688 296312 317694
rect 296260 317630 296312 317636
rect 296166 317520 296222 317529
rect 296166 317455 296222 317464
rect 296168 313200 296220 313206
rect 296168 313142 296220 313148
rect 296180 225758 296208 313142
rect 296272 235074 296300 317630
rect 296364 317354 296392 319756
rect 296502 319716 296530 320076
rect 296594 319938 296622 320076
rect 296582 319932 296634 319938
rect 296582 319874 296634 319880
rect 296686 319818 296714 320076
rect 296456 319688 296530 319716
rect 296640 319790 296714 319818
rect 296456 319054 296484 319688
rect 296536 319592 296588 319598
rect 296536 319534 296588 319540
rect 296548 319054 296576 319534
rect 296444 319048 296496 319054
rect 296444 318990 296496 318996
rect 296536 319048 296588 319054
rect 296536 318990 296588 318996
rect 296442 318880 296498 318889
rect 296442 318815 296498 318824
rect 296352 317348 296404 317354
rect 296352 317290 296404 317296
rect 296456 312866 296484 318815
rect 296640 318696 296668 319790
rect 296778 319716 296806 320076
rect 296962 319920 296990 320076
rect 296732 319688 296806 319716
rect 296916 319892 296990 319920
rect 296732 318889 296760 319688
rect 296916 319546 296944 319892
rect 297054 319852 297082 320076
rect 296824 319518 296944 319546
rect 297008 319824 297082 319852
rect 296718 318880 296774 318889
rect 296718 318815 296774 318824
rect 296548 318668 296668 318696
rect 296548 313274 296576 318668
rect 296628 318504 296680 318510
rect 296628 318446 296680 318452
rect 296640 317762 296668 318446
rect 296628 317756 296680 317762
rect 296628 317698 296680 317704
rect 296824 317286 296852 319518
rect 296902 318472 296958 318481
rect 296902 318407 296958 318416
rect 296812 317280 296864 317286
rect 296812 317222 296864 317228
rect 296628 316736 296680 316742
rect 296628 316678 296680 316684
rect 296536 313268 296588 313274
rect 296536 313210 296588 313216
rect 296444 312860 296496 312866
rect 296444 312802 296496 312808
rect 296640 238814 296668 316678
rect 296916 304366 296944 318407
rect 297008 307630 297036 319824
rect 297146 319784 297174 320076
rect 297238 319954 297266 320076
rect 299064 320104 299120 320113
rect 297316 320039 297372 320048
rect 297238 319926 297312 319954
rect 297100 319756 297174 319784
rect 297100 318374 297128 319756
rect 297178 318880 297234 318889
rect 297178 318815 297234 318824
rect 297088 318368 297140 318374
rect 297088 318310 297140 318316
rect 297086 317520 297142 317529
rect 297086 317455 297142 317464
rect 296996 307624 297048 307630
rect 296996 307566 297048 307572
rect 296904 304360 296956 304366
rect 296904 304302 296956 304308
rect 296628 238808 296680 238814
rect 296628 238750 296680 238756
rect 296260 235068 296312 235074
rect 296260 235010 296312 235016
rect 296720 231124 296772 231130
rect 296720 231066 296772 231072
rect 296168 225752 296220 225758
rect 296168 225694 296220 225700
rect 296076 221876 296128 221882
rect 296076 221818 296128 221824
rect 296732 16574 296760 231066
rect 297100 229498 297128 317455
rect 297192 239426 297220 318815
rect 297284 317490 297312 319926
rect 297422 319784 297450 320076
rect 297376 319756 297450 319784
rect 297376 318986 297404 319756
rect 297514 319716 297542 320076
rect 297606 319784 297634 320076
rect 297882 319784 297910 320076
rect 297974 319818 298002 320076
rect 298158 319920 298186 320076
rect 298112 319892 298186 319920
rect 297974 319790 298048 319818
rect 297606 319756 297772 319784
rect 297514 319688 297588 319716
rect 297364 318980 297416 318986
rect 297364 318922 297416 318928
rect 297364 317756 297416 317762
rect 297364 317698 297416 317704
rect 297272 317484 297324 317490
rect 297272 317426 297324 317432
rect 297180 239420 297232 239426
rect 297180 239362 297232 239368
rect 297088 229492 297140 229498
rect 297088 229434 297140 229440
rect 297376 221542 297404 317698
rect 297456 312860 297508 312866
rect 297456 312802 297508 312808
rect 297468 235657 297496 312802
rect 297560 304298 297588 319688
rect 297744 313818 297772 319756
rect 297836 319756 297910 319784
rect 297836 314022 297864 319756
rect 298020 319138 298048 319790
rect 297928 319110 298048 319138
rect 297928 318753 297956 319110
rect 298112 319002 298140 319892
rect 298250 319818 298278 320076
rect 298342 319938 298370 320076
rect 298330 319932 298382 319938
rect 298330 319874 298382 319880
rect 298020 318974 298140 319002
rect 298204 319790 298278 319818
rect 297914 318744 297970 318753
rect 297914 318679 297970 318688
rect 298020 317234 298048 318974
rect 298100 318844 298152 318850
rect 298100 318786 298152 318792
rect 298112 318238 298140 318786
rect 298100 318232 298152 318238
rect 298100 318174 298152 318180
rect 298204 318084 298232 319790
rect 298434 319784 298462 320076
rect 298388 319756 298462 319784
rect 298284 319728 298336 319734
rect 298284 319670 298336 319676
rect 298296 318850 298324 319670
rect 298284 318844 298336 318850
rect 298284 318786 298336 318792
rect 298284 318640 298336 318646
rect 298284 318582 298336 318588
rect 298112 318056 298232 318084
rect 298112 317393 298140 318056
rect 298192 317552 298244 317558
rect 298192 317494 298244 317500
rect 298098 317384 298154 317393
rect 298098 317319 298154 317328
rect 298020 317206 298140 317234
rect 297824 314016 297876 314022
rect 297824 313958 297876 313964
rect 297732 313812 297784 313818
rect 297732 313754 297784 313760
rect 298112 312905 298140 317206
rect 298098 312896 298154 312905
rect 298098 312831 298154 312840
rect 297548 304292 297600 304298
rect 297548 304234 297600 304240
rect 298204 296714 298232 317494
rect 298112 296686 298232 296714
rect 298112 237182 298140 296686
rect 298296 241777 298324 318582
rect 298388 317626 298416 319756
rect 298526 319716 298554 320076
rect 298710 319938 298738 320076
rect 298802 319938 298830 320076
rect 298698 319932 298750 319938
rect 298698 319874 298750 319880
rect 298790 319932 298842 319938
rect 298790 319874 298842 319880
rect 298894 319784 298922 320076
rect 298480 319688 298554 319716
rect 298848 319756 298922 319784
rect 298480 317898 298508 319688
rect 298744 319660 298796 319666
rect 298744 319602 298796 319608
rect 298560 319592 298612 319598
rect 298560 319534 298612 319540
rect 298468 317892 298520 317898
rect 298468 317834 298520 317840
rect 298376 317620 298428 317626
rect 298376 317562 298428 317568
rect 298572 312769 298600 319534
rect 298756 317830 298784 319602
rect 298744 317824 298796 317830
rect 298744 317766 298796 317772
rect 298848 317642 298876 319756
rect 298986 319716 299014 320076
rect 299708 320104 299764 320113
rect 299064 320039 299120 320048
rect 299170 319870 299198 320076
rect 299262 319938 299290 320076
rect 299250 319932 299302 319938
rect 299250 319874 299302 319880
rect 299158 319864 299210 319870
rect 299538 319852 299566 320076
rect 299158 319806 299210 319812
rect 299492 319824 299566 319852
rect 298940 319688 299014 319716
rect 298940 318753 298968 319688
rect 299388 319592 299440 319598
rect 299388 319534 299440 319540
rect 299296 319456 299348 319462
rect 299296 319398 299348 319404
rect 299018 318880 299074 318889
rect 299018 318815 299074 318824
rect 298926 318744 298982 318753
rect 298926 318679 298982 318688
rect 298756 317614 298876 317642
rect 298756 314226 298784 317614
rect 298836 317484 298888 317490
rect 298836 317426 298888 317432
rect 298744 314220 298796 314226
rect 298744 314162 298796 314168
rect 298558 312760 298614 312769
rect 298558 312695 298614 312704
rect 298744 311160 298796 311166
rect 298744 311102 298796 311108
rect 298282 241768 298338 241777
rect 298282 241703 298338 241712
rect 298100 237176 298152 237182
rect 298100 237118 298152 237124
rect 298756 235686 298784 311102
rect 298744 235680 298796 235686
rect 297454 235648 297510 235657
rect 298744 235622 298796 235628
rect 297454 235583 297510 235592
rect 298008 231124 298060 231130
rect 298008 231066 298060 231072
rect 298020 230450 298048 231066
rect 298008 230444 298060 230450
rect 298008 230386 298060 230392
rect 297364 221536 297416 221542
rect 297364 221478 297416 221484
rect 298098 188320 298154 188329
rect 298098 188255 298154 188264
rect 296732 16546 297312 16574
rect 296076 3596 296128 3602
rect 296076 3538 296128 3544
rect 295984 3460 296036 3466
rect 295984 3402 296036 3408
rect 296088 480 296116 3538
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 188255
rect 298756 3602 298784 235622
rect 298848 234258 298876 317426
rect 298836 234252 298888 234258
rect 298836 234194 298888 234200
rect 299032 231538 299060 318815
rect 299202 318744 299258 318753
rect 299202 318679 299258 318688
rect 299112 314560 299164 314566
rect 299112 314502 299164 314508
rect 299124 311166 299152 314502
rect 299112 311160 299164 311166
rect 299112 311102 299164 311108
rect 299216 234462 299244 318679
rect 299308 318322 299336 319398
rect 299400 318646 299428 319534
rect 299388 318640 299440 318646
rect 299388 318582 299440 318588
rect 299308 318294 299428 318322
rect 299296 318232 299348 318238
rect 299296 318174 299348 318180
rect 299308 314566 299336 318174
rect 299400 315110 299428 318294
rect 299492 317937 299520 319824
rect 299630 319784 299658 320076
rect 300260 320104 300316 320113
rect 299708 320039 299764 320048
rect 299814 319784 299842 320076
rect 299584 319756 299658 319784
rect 299768 319756 299842 319784
rect 299478 317928 299534 317937
rect 299478 317863 299534 317872
rect 299584 317694 299612 319756
rect 299662 318880 299718 318889
rect 299662 318815 299718 318824
rect 299572 317688 299624 317694
rect 299572 317630 299624 317636
rect 299388 315104 299440 315110
rect 299388 315046 299440 315052
rect 299296 314560 299348 314566
rect 299296 314502 299348 314508
rect 299676 311894 299704 318815
rect 299768 315994 299796 319756
rect 299906 319648 299934 320076
rect 299998 319716 300026 320076
rect 300090 319870 300118 320076
rect 300182 319920 300210 320076
rect 300720 320104 300776 320113
rect 300260 320039 300316 320048
rect 300366 319920 300394 320076
rect 300182 319892 300256 319920
rect 300078 319864 300130 319870
rect 300078 319806 300130 319812
rect 300228 319716 300256 319892
rect 299998 319688 300072 319716
rect 299906 319620 299980 319648
rect 299846 319424 299902 319433
rect 299846 319359 299902 319368
rect 299756 315988 299808 315994
rect 299756 315930 299808 315936
rect 299676 311866 299796 311894
rect 299768 305697 299796 311866
rect 299754 305688 299810 305697
rect 299754 305623 299810 305632
rect 299204 234456 299256 234462
rect 299204 234398 299256 234404
rect 299020 231532 299072 231538
rect 299020 231474 299072 231480
rect 299860 231470 299888 319359
rect 299952 318306 299980 319620
rect 299940 318300 299992 318306
rect 299940 318242 299992 318248
rect 300044 317914 300072 319688
rect 299952 317886 300072 317914
rect 300136 319688 300256 319716
rect 300320 319892 300394 319920
rect 299952 315586 299980 317886
rect 300032 317824 300084 317830
rect 300032 317766 300084 317772
rect 299940 315580 299992 315586
rect 299940 315522 299992 315528
rect 300044 313206 300072 317766
rect 300136 317558 300164 319688
rect 300216 319592 300268 319598
rect 300216 319534 300268 319540
rect 300228 318306 300256 319534
rect 300216 318300 300268 318306
rect 300216 318242 300268 318248
rect 300216 318164 300268 318170
rect 300216 318106 300268 318112
rect 300124 317552 300176 317558
rect 300124 317494 300176 317500
rect 300124 313404 300176 313410
rect 300124 313346 300176 313352
rect 300032 313200 300084 313206
rect 300032 313142 300084 313148
rect 300136 311658 300164 313346
rect 300044 311630 300164 311658
rect 300044 306374 300072 311630
rect 300124 311500 300176 311506
rect 300124 311442 300176 311448
rect 300136 311114 300164 311442
rect 300228 311250 300256 318106
rect 300320 317830 300348 319892
rect 300458 319818 300486 320076
rect 300550 319920 300578 320076
rect 302100 320104 302156 320113
rect 300720 320039 300776 320048
rect 300550 319892 300624 319920
rect 300596 319852 300624 319892
rect 300826 319852 300854 320076
rect 300596 319824 300670 319852
rect 300412 319790 300486 319818
rect 300412 319512 300440 319790
rect 300642 319784 300670 319824
rect 300596 319756 300670 319784
rect 300780 319824 300854 319852
rect 300412 319484 300532 319512
rect 300398 319424 300454 319433
rect 300398 319359 300454 319368
rect 300308 317824 300360 317830
rect 300308 317766 300360 317772
rect 300308 317620 300360 317626
rect 300308 317562 300360 317568
rect 300320 311506 300348 317562
rect 300308 311500 300360 311506
rect 300308 311442 300360 311448
rect 300228 311222 300348 311250
rect 300136 311086 300256 311114
rect 300044 306346 300164 306374
rect 299848 231464 299900 231470
rect 299848 231406 299900 231412
rect 299572 228336 299624 228342
rect 299572 228278 299624 228284
rect 299584 227798 299612 228278
rect 299572 227792 299624 227798
rect 299572 227734 299624 227740
rect 298744 3596 298796 3602
rect 298744 3538 298796 3544
rect 299584 3466 299612 227734
rect 300136 217870 300164 306346
rect 300228 227798 300256 311086
rect 300320 232558 300348 311222
rect 300412 240922 300440 319359
rect 300504 317490 300532 319484
rect 300596 317529 300624 319756
rect 300780 319682 300808 319824
rect 300918 319784 300946 320076
rect 301102 319784 301130 320076
rect 300918 319756 300992 319784
rect 300688 319654 300808 319682
rect 300582 317520 300638 317529
rect 300492 317484 300544 317490
rect 300582 317455 300638 317464
rect 300492 317426 300544 317432
rect 300492 315988 300544 315994
rect 300492 315930 300544 315936
rect 300504 300121 300532 315930
rect 300688 315246 300716 319654
rect 300768 319592 300820 319598
rect 300768 319534 300820 319540
rect 300780 318714 300808 319534
rect 300860 319456 300912 319462
rect 300860 319398 300912 319404
rect 300768 318708 300820 318714
rect 300768 318650 300820 318656
rect 300872 318578 300900 319398
rect 300860 318572 300912 318578
rect 300860 318514 300912 318520
rect 300860 318368 300912 318374
rect 300860 318310 300912 318316
rect 300768 318300 300820 318306
rect 300768 318242 300820 318248
rect 300676 315240 300728 315246
rect 300676 315182 300728 315188
rect 300780 312633 300808 318242
rect 300766 312624 300822 312633
rect 300766 312559 300822 312568
rect 300490 300112 300546 300121
rect 300490 300047 300546 300056
rect 300872 291825 300900 318310
rect 300964 317529 300992 319756
rect 301056 319756 301130 319784
rect 301056 319462 301084 319756
rect 301194 319716 301222 320076
rect 301286 319938 301314 320076
rect 301378 319938 301406 320076
rect 301274 319932 301326 319938
rect 301274 319874 301326 319880
rect 301366 319932 301418 319938
rect 301366 319874 301418 319880
rect 301470 319870 301498 320076
rect 301458 319864 301510 319870
rect 301458 319806 301510 319812
rect 301320 319796 301372 319802
rect 301320 319738 301372 319744
rect 301148 319688 301222 319716
rect 301044 319456 301096 319462
rect 301044 319398 301096 319404
rect 301042 318880 301098 318889
rect 301042 318815 301098 318824
rect 301056 318782 301084 318815
rect 301044 318776 301096 318782
rect 301044 318718 301096 318724
rect 301044 318640 301096 318646
rect 301044 318582 301096 318588
rect 300950 317520 301006 317529
rect 300950 317455 301006 317464
rect 301056 316062 301084 318582
rect 301148 317762 301176 319688
rect 301332 319546 301360 319738
rect 301412 319728 301464 319734
rect 301562 319716 301590 320076
rect 301654 319784 301682 320076
rect 301746 319938 301774 320076
rect 301734 319932 301786 319938
rect 301734 319874 301786 319880
rect 301838 319818 301866 320076
rect 301930 319938 301958 320076
rect 301918 319932 301970 319938
rect 301918 319874 301970 319880
rect 301792 319790 301866 319818
rect 301654 319756 301728 319784
rect 301412 319670 301464 319676
rect 301516 319688 301590 319716
rect 301240 319518 301360 319546
rect 301240 317762 301268 319518
rect 301320 319456 301372 319462
rect 301320 319398 301372 319404
rect 301136 317756 301188 317762
rect 301136 317698 301188 317704
rect 301228 317756 301280 317762
rect 301228 317698 301280 317704
rect 301044 316056 301096 316062
rect 301044 315998 301096 316004
rect 300952 311160 301004 311166
rect 300952 311102 301004 311108
rect 300858 291816 300914 291825
rect 300858 291751 300914 291760
rect 300400 240916 300452 240922
rect 300400 240858 300452 240864
rect 300964 233986 300992 311102
rect 301332 300393 301360 319398
rect 301424 317914 301452 319670
rect 301516 318034 301544 319688
rect 301596 319592 301648 319598
rect 301596 319534 301648 319540
rect 301608 319462 301636 319534
rect 301596 319456 301648 319462
rect 301596 319398 301648 319404
rect 301504 318028 301556 318034
rect 301504 317970 301556 317976
rect 301424 317886 301544 317914
rect 301412 317824 301464 317830
rect 301412 317766 301464 317772
rect 301424 312361 301452 317766
rect 301516 313041 301544 317886
rect 301700 315722 301728 319756
rect 301792 318102 301820 319790
rect 301872 319728 301924 319734
rect 302022 319716 302050 320076
rect 302744 320104 302800 320113
rect 302100 320039 302156 320048
rect 302206 319920 302234 320076
rect 302160 319892 302234 319920
rect 302022 319688 302096 319716
rect 301872 319670 301924 319676
rect 301780 318096 301832 318102
rect 301780 318038 301832 318044
rect 301688 315716 301740 315722
rect 301688 315658 301740 315664
rect 301502 313032 301558 313041
rect 301502 312967 301558 312976
rect 301410 312352 301466 312361
rect 301410 312287 301466 312296
rect 301884 311894 301912 319670
rect 301964 319592 302016 319598
rect 301964 319534 302016 319540
rect 301976 317778 302004 319534
rect 302068 318510 302096 319688
rect 302160 319598 302188 319892
rect 302298 319852 302326 320076
rect 302252 319824 302326 319852
rect 302148 319592 302200 319598
rect 302148 319534 302200 319540
rect 302146 319424 302202 319433
rect 302146 319359 302202 319368
rect 302056 318504 302108 318510
rect 302056 318446 302108 318452
rect 301976 317750 302096 317778
rect 301964 317688 302016 317694
rect 301964 317630 302016 317636
rect 301424 311866 301912 311894
rect 301318 300384 301374 300393
rect 301318 300319 301374 300328
rect 300952 233980 301004 233986
rect 300952 233922 301004 233928
rect 300308 232552 300360 232558
rect 300308 232494 300360 232500
rect 300216 227792 300268 227798
rect 300216 227734 300268 227740
rect 301424 224262 301452 311866
rect 301976 311166 302004 317630
rect 302068 315450 302096 317750
rect 302160 317422 302188 319359
rect 302252 318374 302280 319824
rect 302390 319784 302418 320076
rect 302344 319756 302418 319784
rect 302482 319784 302510 320076
rect 302574 319852 302602 320076
rect 302666 319954 302694 320076
rect 303848 320104 303904 320113
rect 302744 320039 302800 320048
rect 302666 319926 302740 319954
rect 302712 319852 302740 319926
rect 302850 319920 302878 320076
rect 302850 319892 302924 319920
rect 302574 319824 302648 319852
rect 302712 319824 302832 319852
rect 302482 319756 302556 319784
rect 302240 318368 302292 318374
rect 302344 318345 302372 319756
rect 302424 319660 302476 319666
rect 302424 319602 302476 319608
rect 302240 318310 302292 318316
rect 302330 318336 302386 318345
rect 302330 318271 302386 318280
rect 302148 317416 302200 317422
rect 302148 317358 302200 317364
rect 302056 315444 302108 315450
rect 302056 315386 302108 315392
rect 301964 311160 302016 311166
rect 301964 311102 302016 311108
rect 302436 298790 302464 319602
rect 302528 319546 302556 319756
rect 302620 319666 302648 319824
rect 302700 319728 302752 319734
rect 302700 319670 302752 319676
rect 302608 319660 302660 319666
rect 302608 319602 302660 319608
rect 302528 319518 302648 319546
rect 302514 319424 302570 319433
rect 302514 319359 302570 319368
rect 302528 319326 302556 319359
rect 302516 319320 302568 319326
rect 302516 319262 302568 319268
rect 302620 316946 302648 319518
rect 302608 316940 302660 316946
rect 302608 316882 302660 316888
rect 302516 315988 302568 315994
rect 302516 315930 302568 315936
rect 302528 301510 302556 315930
rect 302516 301504 302568 301510
rect 302516 301446 302568 301452
rect 302424 298784 302476 298790
rect 302424 298726 302476 298732
rect 302712 238134 302740 319670
rect 302804 318170 302832 319824
rect 302792 318164 302844 318170
rect 302792 318106 302844 318112
rect 302896 317830 302924 319892
rect 303034 319852 303062 320076
rect 302988 319824 303062 319852
rect 302988 318850 303016 319824
rect 303126 319784 303154 320076
rect 303080 319756 303154 319784
rect 302976 318844 303028 318850
rect 302976 318786 303028 318792
rect 302974 318744 303030 318753
rect 302974 318679 303030 318688
rect 302988 318481 303016 318679
rect 302974 318472 303030 318481
rect 302974 318407 303030 318416
rect 302884 317824 302936 317830
rect 302884 317766 302936 317772
rect 303080 317642 303108 319756
rect 303218 319716 303246 320076
rect 303310 319938 303338 320076
rect 303298 319932 303350 319938
rect 303298 319874 303350 319880
rect 303402 319818 303430 320076
rect 303494 319938 303522 320076
rect 303482 319932 303534 319938
rect 303482 319874 303534 319880
rect 302988 317614 303108 317642
rect 303172 319688 303246 319716
rect 303356 319790 303430 319818
rect 302884 315580 302936 315586
rect 302884 315522 302936 315528
rect 302700 238128 302752 238134
rect 302700 238070 302752 238076
rect 302238 231160 302294 231169
rect 302238 231095 302294 231104
rect 302054 227624 302110 227633
rect 302054 227559 302110 227568
rect 302068 227186 302096 227559
rect 302056 227180 302108 227186
rect 302056 227122 302108 227128
rect 302068 226370 302096 227122
rect 302056 226364 302108 226370
rect 302056 226306 302108 226312
rect 301412 224256 301464 224262
rect 301412 224198 301464 224204
rect 300124 217864 300176 217870
rect 300124 217806 300176 217812
rect 300136 3534 300164 217806
rect 302252 16574 302280 231095
rect 302896 223106 302924 315522
rect 302988 312225 303016 317614
rect 303068 317552 303120 317558
rect 303068 317494 303120 317500
rect 302974 312216 303030 312225
rect 302974 312151 303030 312160
rect 302976 312112 303028 312118
rect 302976 312054 303028 312060
rect 302988 229945 303016 312054
rect 303080 311574 303108 317494
rect 303172 315994 303200 319688
rect 303252 318844 303304 318850
rect 303252 318786 303304 318792
rect 303160 315988 303212 315994
rect 303160 315930 303212 315936
rect 303160 315240 303212 315246
rect 303160 315182 303212 315188
rect 303172 312118 303200 315182
rect 303160 312112 303212 312118
rect 303160 312054 303212 312060
rect 303068 311568 303120 311574
rect 303068 311510 303120 311516
rect 302974 229936 303030 229945
rect 302974 229871 303030 229880
rect 303264 227254 303292 318786
rect 303356 315489 303384 319790
rect 303586 319784 303614 320076
rect 303678 319818 303706 320076
rect 303770 319938 303798 320076
rect 304400 320104 304456 320113
rect 303848 320039 303904 320048
rect 303758 319932 303810 319938
rect 303758 319874 303810 319880
rect 303678 319790 303752 319818
rect 303540 319756 303614 319784
rect 303436 319728 303488 319734
rect 303436 319670 303488 319676
rect 303448 318442 303476 319670
rect 303436 318436 303488 318442
rect 303436 318378 303488 318384
rect 303436 317960 303488 317966
rect 303436 317902 303488 317908
rect 303448 316674 303476 317902
rect 303436 316668 303488 316674
rect 303436 316610 303488 316616
rect 303540 315654 303568 319756
rect 303724 318322 303752 319790
rect 303804 319796 303856 319802
rect 303954 319784 303982 320076
rect 304046 319938 304074 320076
rect 304034 319932 304086 319938
rect 304034 319874 304086 319880
rect 304138 319784 304166 320076
rect 303954 319756 304028 319784
rect 303804 319738 303856 319744
rect 303816 318646 303844 319738
rect 303804 318640 303856 318646
rect 303804 318582 303856 318588
rect 303632 318294 303752 318322
rect 303632 317082 303660 318294
rect 303710 318200 303766 318209
rect 303710 318135 303766 318144
rect 303620 317076 303672 317082
rect 303620 317018 303672 317024
rect 303724 317014 303752 318135
rect 303804 317824 303856 317830
rect 303804 317766 303856 317772
rect 303816 317490 303844 317766
rect 304000 317694 304028 319756
rect 304092 319756 304166 319784
rect 304322 319784 304350 320076
rect 305136 320104 305192 320113
rect 304400 320039 304456 320048
rect 304506 319852 304534 320076
rect 304460 319824 304534 319852
rect 304322 319756 304396 319784
rect 303988 317688 304040 317694
rect 303988 317630 304040 317636
rect 303804 317484 303856 317490
rect 303804 317426 303856 317432
rect 303988 317484 304040 317490
rect 303988 317426 304040 317432
rect 303712 317008 303764 317014
rect 303712 316950 303764 316956
rect 303896 316056 303948 316062
rect 303896 315998 303948 316004
rect 303804 315988 303856 315994
rect 303804 315930 303856 315936
rect 303528 315648 303580 315654
rect 303528 315590 303580 315596
rect 303342 315480 303398 315489
rect 303342 315415 303398 315424
rect 303816 307426 303844 315930
rect 303908 307494 303936 315998
rect 303896 307488 303948 307494
rect 303896 307430 303948 307436
rect 303804 307420 303856 307426
rect 303804 307362 303856 307368
rect 303710 233200 303766 233209
rect 303710 233135 303766 233144
rect 303724 233102 303752 233135
rect 303712 233096 303764 233102
rect 303712 233038 303764 233044
rect 303724 231878 303752 233038
rect 303712 231872 303764 231878
rect 303712 231814 303764 231820
rect 303620 228404 303672 228410
rect 303620 228346 303672 228352
rect 303632 228002 303660 228346
rect 303620 227996 303672 228002
rect 303620 227938 303672 227944
rect 303252 227248 303304 227254
rect 303252 227190 303304 227196
rect 302884 223100 302936 223106
rect 302884 223042 302936 223048
rect 303434 219192 303490 219201
rect 303434 219127 303490 219136
rect 303448 218958 303476 219127
rect 303436 218952 303488 218958
rect 303436 218894 303488 218900
rect 303448 218074 303476 218894
rect 303436 218068 303488 218074
rect 303436 218010 303488 218016
rect 303632 16574 303660 227938
rect 304000 227526 304028 317426
rect 304092 228274 304120 319756
rect 304264 319592 304316 319598
rect 304264 319534 304316 319540
rect 304170 319424 304226 319433
rect 304170 319359 304226 319368
rect 304184 305726 304212 319359
rect 304276 314430 304304 319534
rect 304368 317966 304396 319756
rect 304356 317960 304408 317966
rect 304356 317902 304408 317908
rect 304264 314424 304316 314430
rect 304264 314366 304316 314372
rect 304460 311894 304488 319824
rect 304598 319784 304626 320076
rect 304552 319756 304626 319784
rect 304552 313138 304580 319756
rect 304690 319682 304718 320076
rect 304782 319870 304810 320076
rect 304874 319938 304902 320076
rect 304862 319932 304914 319938
rect 304862 319874 304914 319880
rect 304770 319864 304822 319870
rect 304770 319806 304822 319812
rect 304966 319784 304994 320076
rect 304644 319654 304718 319682
rect 304920 319756 304994 319784
rect 304644 315994 304672 319654
rect 304920 319648 304948 319756
rect 305058 319682 305086 320076
rect 306056 320104 306112 320113
rect 305136 320039 305192 320048
rect 305242 319938 305270 320076
rect 305334 319938 305362 320076
rect 305230 319932 305282 319938
rect 305230 319874 305282 319880
rect 305322 319932 305374 319938
rect 305322 319874 305374 319880
rect 305426 319870 305454 320076
rect 305518 319938 305546 320076
rect 305506 319932 305558 319938
rect 305506 319874 305558 319880
rect 305414 319864 305466 319870
rect 305414 319806 305466 319812
rect 305184 319796 305236 319802
rect 305184 319738 305236 319744
rect 305276 319796 305328 319802
rect 305610 319784 305638 320076
rect 305276 319738 305328 319744
rect 305564 319756 305638 319784
rect 305058 319654 305132 319682
rect 304828 319620 304948 319648
rect 304724 319592 304776 319598
rect 304724 319534 304776 319540
rect 304736 317665 304764 319534
rect 304722 317656 304778 317665
rect 304722 317591 304778 317600
rect 304828 316062 304856 319620
rect 304998 318880 305054 318889
rect 304998 318815 305054 318824
rect 305012 316810 305040 318815
rect 305104 317665 305132 319654
rect 305090 317656 305146 317665
rect 305090 317591 305146 317600
rect 305196 317529 305224 319738
rect 305288 317801 305316 319738
rect 305368 319728 305420 319734
rect 305368 319670 305420 319676
rect 305380 319546 305408 319670
rect 305380 319518 305500 319546
rect 305368 319456 305420 319462
rect 305368 319398 305420 319404
rect 305274 317792 305330 317801
rect 305274 317727 305330 317736
rect 305276 317688 305328 317694
rect 305276 317630 305328 317636
rect 305182 317520 305238 317529
rect 305182 317455 305238 317464
rect 305000 316804 305052 316810
rect 305000 316746 305052 316752
rect 304816 316056 304868 316062
rect 304816 315998 304868 316004
rect 304632 315988 304684 315994
rect 304632 315930 304684 315936
rect 304540 313132 304592 313138
rect 304540 313074 304592 313080
rect 305288 311894 305316 317630
rect 304276 311866 304488 311894
rect 305196 311866 305316 311894
rect 304276 307358 304304 311866
rect 304264 307352 304316 307358
rect 304264 307294 304316 307300
rect 304172 305720 304224 305726
rect 304172 305662 304224 305668
rect 304264 300416 304316 300422
rect 304264 300358 304316 300364
rect 304080 228268 304132 228274
rect 304080 228210 304132 228216
rect 304276 228002 304304 300358
rect 304264 227996 304316 228002
rect 304264 227938 304316 227944
rect 303988 227520 304040 227526
rect 303988 227462 304040 227468
rect 305196 221610 305224 311866
rect 305380 230450 305408 319398
rect 305472 317558 305500 319518
rect 305460 317552 305512 317558
rect 305564 317529 305592 319756
rect 305702 319716 305730 320076
rect 305656 319688 305730 319716
rect 305794 319716 305822 320076
rect 305886 319784 305914 320076
rect 305978 319938 306006 320076
rect 306240 320104 306296 320113
rect 306056 320039 306112 320048
rect 305966 319932 306018 319938
rect 305966 319874 306018 319880
rect 306162 319784 306190 320076
rect 306884 320104 306940 320113
rect 306240 320039 306296 320048
rect 306346 319852 306374 320076
rect 305886 319756 306052 319784
rect 305794 319688 305868 319716
rect 305460 317494 305512 317500
rect 305550 317520 305606 317529
rect 305550 317455 305606 317464
rect 305656 317150 305684 319688
rect 305734 319424 305790 319433
rect 305734 319359 305790 319368
rect 305644 317144 305696 317150
rect 305644 317086 305696 317092
rect 305748 316010 305776 319359
rect 305840 317694 305868 319688
rect 305920 319660 305972 319666
rect 305920 319602 305972 319608
rect 305932 317937 305960 319602
rect 305918 317928 305974 317937
rect 305918 317863 305974 317872
rect 305828 317688 305880 317694
rect 305828 317630 305880 317636
rect 305828 317552 305880 317558
rect 305828 317494 305880 317500
rect 305564 315982 305776 316010
rect 305564 300422 305592 315982
rect 305840 311894 305868 317494
rect 306024 313410 306052 319756
rect 306116 319756 306190 319784
rect 306300 319824 306374 319852
rect 306116 319025 306144 319756
rect 306300 319682 306328 319824
rect 306438 319784 306466 320076
rect 306530 319938 306558 320076
rect 306518 319932 306570 319938
rect 306518 319874 306570 319880
rect 306622 319784 306650 320076
rect 306714 319938 306742 320076
rect 306702 319932 306754 319938
rect 306702 319874 306754 319880
rect 306806 319784 306834 320076
rect 307160 320104 307216 320113
rect 306884 320039 306940 320048
rect 306208 319654 306328 319682
rect 306392 319756 306466 319784
rect 306576 319756 306650 319784
rect 306760 319756 306834 319784
rect 306102 319016 306158 319025
rect 306102 318951 306158 318960
rect 306104 317620 306156 317626
rect 306104 317562 306156 317568
rect 306116 315314 306144 317562
rect 306208 315858 306236 319654
rect 306286 319424 306342 319433
rect 306286 319359 306342 319368
rect 306300 317626 306328 319359
rect 306288 317620 306340 317626
rect 306288 317562 306340 317568
rect 306392 317506 306420 319756
rect 306472 319660 306524 319666
rect 306472 319602 306524 319608
rect 306300 317478 306420 317506
rect 306196 315852 306248 315858
rect 306196 315794 306248 315800
rect 306104 315308 306156 315314
rect 306104 315250 306156 315256
rect 306012 313404 306064 313410
rect 306012 313346 306064 313352
rect 305656 311866 305868 311894
rect 305552 300416 305604 300422
rect 305552 300358 305604 300364
rect 305368 230444 305420 230450
rect 305368 230386 305420 230392
rect 305656 228614 305684 311866
rect 306104 230172 306156 230178
rect 306104 230114 306156 230120
rect 306116 229265 306144 230114
rect 306102 229256 306158 229265
rect 306102 229191 306158 229200
rect 306116 229158 306144 229191
rect 306104 229152 306156 229158
rect 306104 229094 306156 229100
rect 305644 228608 305696 228614
rect 305644 228550 305696 228556
rect 305274 226264 305330 226273
rect 305274 226199 305330 226208
rect 305288 225894 305316 226199
rect 305276 225888 305328 225894
rect 305276 225830 305328 225836
rect 305288 225010 305316 225830
rect 305276 225004 305328 225010
rect 305276 224946 305328 224952
rect 305184 221604 305236 221610
rect 305184 221546 305236 221552
rect 304998 213208 305054 213217
rect 304998 213143 305054 213152
rect 305012 16574 305040 213143
rect 305092 208344 305144 208350
rect 305092 208286 305144 208292
rect 305104 207942 305132 208286
rect 305092 207936 305144 207942
rect 305092 207878 305144 207884
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 300124 3528 300176 3534
rect 300124 3470 300176 3476
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 299572 3460 299624 3466
rect 299572 3402 299624 3408
rect 300768 3460 300820 3466
rect 300768 3402 300820 3408
rect 299664 3392 299716 3398
rect 299664 3334 299716 3340
rect 299676 480 299704 3334
rect 300780 480 300808 3402
rect 301976 480 302004 3470
rect 303172 480 303200 16546
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 305656 3466 305684 228550
rect 306300 207942 306328 317478
rect 306380 315988 306432 315994
rect 306380 315930 306432 315936
rect 306392 315722 306420 315930
rect 306380 315716 306432 315722
rect 306380 315658 306432 315664
rect 306484 228750 306512 319602
rect 306576 316062 306604 319756
rect 306760 319682 306788 319756
rect 306990 319716 307018 320076
rect 307082 319818 307110 320076
rect 307620 320104 307676 320113
rect 307160 320039 307216 320048
rect 307266 319852 307294 320076
rect 307220 319824 307294 319852
rect 307082 319790 307156 319818
rect 306990 319688 307064 319716
rect 306668 319654 306788 319682
rect 306668 318238 306696 319654
rect 306932 319592 306984 319598
rect 306932 319534 306984 319540
rect 306838 319424 306894 319433
rect 306838 319359 306894 319368
rect 306746 319288 306802 319297
rect 306746 319223 306802 319232
rect 306656 318232 306708 318238
rect 306656 318174 306708 318180
rect 306564 316056 306616 316062
rect 306564 315998 306616 316004
rect 306656 315988 306708 315994
rect 306656 315930 306708 315936
rect 306564 315920 306616 315926
rect 306564 315862 306616 315868
rect 306576 231606 306604 315862
rect 306668 239222 306696 315930
rect 306760 240106 306788 319223
rect 306852 316198 306880 319359
rect 306840 316192 306892 316198
rect 306840 316134 306892 316140
rect 306840 316056 306892 316062
rect 306840 315998 306892 316004
rect 306852 260166 306880 315998
rect 306944 311894 306972 319534
rect 307036 317529 307064 319688
rect 307128 317762 307156 319790
rect 307116 317756 307168 317762
rect 307116 317698 307168 317704
rect 307022 317520 307078 317529
rect 307022 317455 307078 317464
rect 307024 316192 307076 316198
rect 307024 316134 307076 316140
rect 307036 315790 307064 316134
rect 307024 315784 307076 315790
rect 307024 315726 307076 315732
rect 306944 311866 307156 311894
rect 307128 311409 307156 311866
rect 307114 311400 307170 311409
rect 307114 311335 307170 311344
rect 306840 260160 306892 260166
rect 306840 260102 306892 260108
rect 306748 240100 306800 240106
rect 306748 240042 306800 240048
rect 306656 239216 306708 239222
rect 306656 239158 306708 239164
rect 306668 234394 306696 239158
rect 306656 234388 306708 234394
rect 306656 234330 306708 234336
rect 306564 231600 306616 231606
rect 306564 231542 306616 231548
rect 306472 228744 306524 228750
rect 306472 228686 306524 228692
rect 306484 227798 306512 228686
rect 306472 227792 306524 227798
rect 306472 227734 306524 227740
rect 307220 211070 307248 319824
rect 307358 319784 307386 320076
rect 307312 319756 307386 319784
rect 307312 315926 307340 319756
rect 307450 319716 307478 320076
rect 307542 319954 307570 320076
rect 308172 320104 308228 320113
rect 307620 320039 307676 320048
rect 307542 319926 307616 319954
rect 307404 319688 307478 319716
rect 307404 315994 307432 319688
rect 307484 319592 307536 319598
rect 307482 319560 307484 319569
rect 307536 319560 307538 319569
rect 307482 319495 307538 319504
rect 307588 317665 307616 319926
rect 307726 319852 307754 320076
rect 307680 319824 307754 319852
rect 307574 317656 307630 317665
rect 307574 317591 307630 317600
rect 307576 317484 307628 317490
rect 307576 317426 307628 317432
rect 307392 315988 307444 315994
rect 307392 315930 307444 315936
rect 307300 315920 307352 315926
rect 307300 315862 307352 315868
rect 307588 237114 307616 317426
rect 307680 316062 307708 319824
rect 307818 319784 307846 320076
rect 307772 319756 307846 319784
rect 307668 316056 307720 316062
rect 307668 315998 307720 316004
rect 307772 316010 307800 319756
rect 307910 319716 307938 320076
rect 308002 319784 308030 320076
rect 308094 319852 308122 320076
rect 309736 320104 309792 320113
rect 308172 320039 308228 320048
rect 308278 319954 308306 320076
rect 308232 319926 308306 319954
rect 308370 319954 308398 320076
rect 308554 319954 308582 320076
rect 308370 319926 308444 319954
rect 308508 319938 308582 319954
rect 308094 319824 308168 319852
rect 308002 319756 308076 319784
rect 307864 319688 307938 319716
rect 307864 318617 307892 319688
rect 307850 318608 307906 318617
rect 307850 318543 307906 318552
rect 308048 317558 308076 319756
rect 308036 317552 308088 317558
rect 308036 317494 308088 317500
rect 307772 315982 308076 316010
rect 307944 315852 307996 315858
rect 307944 315794 307996 315800
rect 307668 315648 307720 315654
rect 307668 315590 307720 315596
rect 307576 237108 307628 237114
rect 307576 237050 307628 237056
rect 307588 236706 307616 237050
rect 307576 236700 307628 236706
rect 307576 236642 307628 236648
rect 307576 231600 307628 231606
rect 307576 231542 307628 231548
rect 307588 231198 307616 231542
rect 307576 231192 307628 231198
rect 307576 231134 307628 231140
rect 307680 213858 307708 315590
rect 307956 228478 307984 315794
rect 308048 311273 308076 315982
rect 308140 315926 308168 319824
rect 308232 317490 308260 319926
rect 308312 319864 308364 319870
rect 308312 319806 308364 319812
rect 308220 317484 308272 317490
rect 308220 317426 308272 317432
rect 308324 316946 308352 319806
rect 308312 316940 308364 316946
rect 308312 316882 308364 316888
rect 308312 316736 308364 316742
rect 308312 316678 308364 316684
rect 308128 315920 308180 315926
rect 308128 315862 308180 315868
rect 308324 311894 308352 316678
rect 308416 315994 308444 319926
rect 308496 319932 308582 319938
rect 308548 319926 308582 319932
rect 308496 319874 308548 319880
rect 308646 319852 308674 320076
rect 308600 319824 308674 319852
rect 308494 319424 308550 319433
rect 308494 319359 308550 319368
rect 308508 317801 308536 319359
rect 308494 317792 308550 317801
rect 308494 317727 308550 317736
rect 308496 317620 308548 317626
rect 308496 317562 308548 317568
rect 308404 315988 308456 315994
rect 308404 315930 308456 315936
rect 308508 315450 308536 317562
rect 308496 315444 308548 315450
rect 308496 315386 308548 315392
rect 308324 311866 308444 311894
rect 308034 311264 308090 311273
rect 308034 311199 308090 311208
rect 308416 238066 308444 311866
rect 308404 238060 308456 238066
rect 308404 238002 308456 238008
rect 307944 228472 307996 228478
rect 307944 228414 307996 228420
rect 307668 213852 307720 213858
rect 307668 213794 307720 213800
rect 307680 213246 307708 213794
rect 307668 213240 307720 213246
rect 307668 213182 307720 213188
rect 307208 211064 307260 211070
rect 307208 211006 307260 211012
rect 307668 211064 307720 211070
rect 307668 211006 307720 211012
rect 307680 210458 307708 211006
rect 307668 210452 307720 210458
rect 307668 210394 307720 210400
rect 306288 207936 306340 207942
rect 306288 207878 306340 207884
rect 307024 207936 307076 207942
rect 307024 207878 307076 207884
rect 306748 3664 306800 3670
rect 306748 3606 306800 3612
rect 305644 3460 305696 3466
rect 305644 3402 305696 3408
rect 306760 480 306788 3606
rect 307036 3534 307064 207878
rect 307024 3528 307076 3534
rect 307024 3470 307076 3476
rect 307956 480 307984 228414
rect 308600 222873 308628 319824
rect 308738 319818 308766 320076
rect 308830 319920 308858 320076
rect 308830 319892 308904 319920
rect 308876 319852 308904 319892
rect 308876 319824 308950 319852
rect 308738 319790 308812 319818
rect 308784 319682 308812 319790
rect 308922 319784 308950 319824
rect 309014 319818 309042 320076
rect 309106 319938 309134 320076
rect 309094 319932 309146 319938
rect 309094 319874 309146 319880
rect 309014 319790 309088 319818
rect 308692 319654 308812 319682
rect 308876 319756 308950 319784
rect 308692 317937 308720 319654
rect 308770 319560 308826 319569
rect 308770 319495 308826 319504
rect 308678 317928 308734 317937
rect 308678 317863 308734 317872
rect 308784 316010 308812 319495
rect 308876 317014 308904 319756
rect 308956 319660 309008 319666
rect 308956 319602 309008 319608
rect 308968 317626 308996 319602
rect 309060 318986 309088 319790
rect 309198 319784 309226 320076
rect 309290 319938 309318 320076
rect 309382 319938 309410 320076
rect 309278 319932 309330 319938
rect 309278 319874 309330 319880
rect 309370 319932 309422 319938
rect 309370 319874 309422 319880
rect 309324 319796 309376 319802
rect 309198 319756 309272 319784
rect 309244 319666 309272 319756
rect 309474 319784 309502 320076
rect 309566 319938 309594 320076
rect 309554 319932 309606 319938
rect 309554 319874 309606 319880
rect 309658 319818 309686 320076
rect 310104 320104 310160 320113
rect 309736 320039 309792 320048
rect 309842 319938 309870 320076
rect 309830 319932 309882 319938
rect 309830 319874 309882 319880
rect 310026 319818 310054 320076
rect 310472 320104 310528 320113
rect 310104 320039 310160 320048
rect 310210 319920 310238 320076
rect 310302 319938 310330 320076
rect 310164 319892 310238 319920
rect 310290 319932 310342 319938
rect 310164 319852 310192 319892
rect 310290 319874 310342 319880
rect 309324 319738 309376 319744
rect 309428 319756 309502 319784
rect 309612 319790 309686 319818
rect 309784 319796 309836 319802
rect 309232 319660 309284 319666
rect 309232 319602 309284 319608
rect 309336 319512 309364 319738
rect 309152 319484 309364 319512
rect 309048 318980 309100 318986
rect 309048 318922 309100 318928
rect 308956 317620 309008 317626
rect 308956 317562 309008 317568
rect 309152 317506 309180 319484
rect 309322 319424 309378 319433
rect 309322 319359 309378 319368
rect 309230 319288 309286 319297
rect 309336 319258 309364 319359
rect 309230 319223 309286 319232
rect 309324 319252 309376 319258
rect 309244 319190 309272 319223
rect 309324 319194 309376 319200
rect 309232 319184 309284 319190
rect 309232 319126 309284 319132
rect 308956 317484 309008 317490
rect 308956 317426 309008 317432
rect 309060 317478 309180 317506
rect 308864 317008 308916 317014
rect 308864 316950 308916 316956
rect 308692 315982 308812 316010
rect 308864 315988 308916 315994
rect 308692 311817 308720 315982
rect 308864 315930 308916 315936
rect 308772 315920 308824 315926
rect 308772 315862 308824 315868
rect 308678 311808 308734 311817
rect 308678 311743 308734 311752
rect 308784 311681 308812 315862
rect 308770 311672 308826 311681
rect 308770 311607 308826 311616
rect 308876 223281 308904 315930
rect 308968 259418 308996 317426
rect 308956 259412 309008 259418
rect 308956 259354 309008 259360
rect 309060 245818 309088 317478
rect 309428 316130 309456 319756
rect 309506 319560 309562 319569
rect 309506 319495 309562 319504
rect 309416 316124 309468 316130
rect 309416 316066 309468 316072
rect 309520 316010 309548 319495
rect 309612 317490 309640 319790
rect 309784 319738 309836 319744
rect 309980 319790 310054 319818
rect 310118 319824 310192 319852
rect 309692 319728 309744 319734
rect 309692 319670 309744 319676
rect 309704 319569 309732 319670
rect 309690 319560 309746 319569
rect 309690 319495 309746 319504
rect 309796 319326 309824 319738
rect 309876 319660 309928 319666
rect 309876 319602 309928 319608
rect 309784 319320 309836 319326
rect 309784 319262 309836 319268
rect 309782 319016 309838 319025
rect 309782 318951 309838 318960
rect 309796 318152 309824 318951
rect 309704 318124 309824 318152
rect 309600 317484 309652 317490
rect 309600 317426 309652 317432
rect 309600 316260 309652 316266
rect 309600 316202 309652 316208
rect 309244 315982 309548 316010
rect 309244 311370 309272 315982
rect 309324 315920 309376 315926
rect 309324 315862 309376 315868
rect 309232 311364 309284 311370
rect 309232 311306 309284 311312
rect 309048 245812 309100 245818
rect 309048 245754 309100 245760
rect 309060 240990 309088 245754
rect 309048 240984 309100 240990
rect 309048 240926 309100 240932
rect 309140 227792 309192 227798
rect 309140 227734 309192 227740
rect 308862 223272 308918 223281
rect 308862 223207 308918 223216
rect 308586 222864 308642 222873
rect 308586 222799 308642 222808
rect 309152 16574 309180 227734
rect 309336 224602 309364 315862
rect 309416 315784 309468 315790
rect 309416 315726 309468 315732
rect 309428 228818 309456 315726
rect 309612 311894 309640 316202
rect 309704 312798 309732 318124
rect 309784 318028 309836 318034
rect 309784 317970 309836 317976
rect 309692 312792 309744 312798
rect 309692 312734 309744 312740
rect 309520 311866 309640 311894
rect 309520 311438 309548 311866
rect 309508 311432 309560 311438
rect 309508 311374 309560 311380
rect 309508 259412 309560 259418
rect 309508 259354 309560 259360
rect 309520 233034 309548 259354
rect 309796 240242 309824 317970
rect 309888 311894 309916 319602
rect 309980 319546 310008 319790
rect 310118 319784 310146 319824
rect 310118 319756 310192 319784
rect 309980 319518 310100 319546
rect 309968 319456 310020 319462
rect 309968 319398 310020 319404
rect 309980 315382 310008 319398
rect 309968 315376 310020 315382
rect 309968 315318 310020 315324
rect 309888 311866 310008 311894
rect 309980 311545 310008 311866
rect 309966 311536 310022 311545
rect 309966 311471 310022 311480
rect 309874 254008 309930 254017
rect 309874 253943 309930 253952
rect 309784 240236 309836 240242
rect 309784 240178 309836 240184
rect 309508 233028 309560 233034
rect 309508 232970 309560 232976
rect 309416 228812 309468 228818
rect 309416 228754 309468 228760
rect 309428 227798 309456 228754
rect 309416 227792 309468 227798
rect 309416 227734 309468 227740
rect 309796 225690 309824 240178
rect 309888 230081 309916 253943
rect 309874 230072 309930 230081
rect 309874 230007 309930 230016
rect 309876 227792 309928 227798
rect 309876 227734 309928 227740
rect 309784 225684 309836 225690
rect 309784 225626 309836 225632
rect 309324 224596 309376 224602
rect 309324 224538 309376 224544
rect 309152 16546 309824 16574
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 309888 3194 309916 227734
rect 310072 223009 310100 319518
rect 310164 319462 310192 319756
rect 310244 319728 310296 319734
rect 310394 319716 310422 320076
rect 310748 320104 310804 320113
rect 310472 320039 310528 320048
rect 310578 319784 310606 320076
rect 310670 319954 310698 320076
rect 312496 320104 312552 320113
rect 310748 320039 310804 320048
rect 310670 319926 310744 319954
rect 310946 319938 310974 320076
rect 310244 319670 310296 319676
rect 310348 319688 310422 319716
rect 310532 319756 310606 319784
rect 310152 319456 310204 319462
rect 310152 319398 310204 319404
rect 310150 319288 310206 319297
rect 310150 319223 310206 319232
rect 310164 233170 310192 319223
rect 310256 316266 310284 319670
rect 310244 316260 310296 316266
rect 310244 316202 310296 316208
rect 310244 316124 310296 316130
rect 310244 316066 310296 316072
rect 310256 311137 310284 316066
rect 310348 315926 310376 319688
rect 310532 315994 310560 319756
rect 310610 319288 310666 319297
rect 310610 319223 310666 319232
rect 310520 315988 310572 315994
rect 310520 315930 310572 315936
rect 310336 315920 310388 315926
rect 310336 315862 310388 315868
rect 310624 311302 310652 319223
rect 310716 319122 310744 319926
rect 310934 319932 310986 319938
rect 310934 319874 310986 319880
rect 310794 319832 310850 319841
rect 311038 319818 311066 320076
rect 311130 319938 311158 320076
rect 311118 319932 311170 319938
rect 311118 319874 311170 319880
rect 311314 319818 311342 320076
rect 311038 319790 311112 319818
rect 310794 319767 310850 319776
rect 310808 319462 310836 319767
rect 310888 319524 310940 319530
rect 310888 319466 310940 319472
rect 310796 319456 310848 319462
rect 310900 319433 310928 319466
rect 310796 319398 310848 319404
rect 310886 319424 310942 319433
rect 310886 319359 310942 319368
rect 310704 319116 310756 319122
rect 310704 319058 310756 319064
rect 310794 319016 310850 319025
rect 310794 318951 310850 318960
rect 310808 316742 310836 318951
rect 310796 316736 310848 316742
rect 310796 316678 310848 316684
rect 310796 316056 310848 316062
rect 310796 315998 310848 316004
rect 310612 311296 310664 311302
rect 310612 311238 310664 311244
rect 310242 311128 310298 311137
rect 310242 311063 310298 311072
rect 310808 245206 310836 315998
rect 310888 315716 310940 315722
rect 310888 315658 310940 315664
rect 310796 245200 310848 245206
rect 310796 245142 310848 245148
rect 310152 233164 310204 233170
rect 310152 233106 310204 233112
rect 310428 233164 310480 233170
rect 310428 233106 310480 233112
rect 310440 232558 310468 233106
rect 310428 232552 310480 232558
rect 310428 232494 310480 232500
rect 310900 229094 310928 315658
rect 311084 315246 311112 319790
rect 311176 319790 311342 319818
rect 311176 316062 311204 319790
rect 311256 319728 311308 319734
rect 311256 319670 311308 319676
rect 311164 316056 311216 316062
rect 311164 315998 311216 316004
rect 311072 315240 311124 315246
rect 311072 315182 311124 315188
rect 311162 312080 311218 312089
rect 311162 312015 311218 312024
rect 311176 235385 311204 312015
rect 311268 311894 311296 319670
rect 311406 319648 311434 320076
rect 311498 319938 311526 320076
rect 311486 319932 311538 319938
rect 311486 319874 311538 319880
rect 311590 319818 311618 320076
rect 311544 319790 311618 319818
rect 311406 319620 311480 319648
rect 311346 319560 311402 319569
rect 311346 319495 311402 319504
rect 311360 319394 311388 319495
rect 311348 319388 311400 319394
rect 311348 319330 311400 319336
rect 311346 319288 311402 319297
rect 311346 319223 311402 319232
rect 311360 312934 311388 319223
rect 311348 312928 311400 312934
rect 311348 312870 311400 312876
rect 311268 311866 311388 311894
rect 311256 245200 311308 245206
rect 311256 245142 311308 245148
rect 311268 244390 311296 245142
rect 311256 244384 311308 244390
rect 311256 244326 311308 244332
rect 311162 235376 311218 235385
rect 311162 235311 311218 235320
rect 311268 231674 311296 244326
rect 311256 231668 311308 231674
rect 311256 231610 311308 231616
rect 311256 230308 311308 230314
rect 311256 230250 311308 230256
rect 311268 229770 311296 230250
rect 311256 229764 311308 229770
rect 311256 229706 311308 229712
rect 310532 229066 310928 229094
rect 310532 228546 310560 229066
rect 310520 228540 310572 228546
rect 310520 228482 310572 228488
rect 310058 223000 310114 223009
rect 310058 222935 310114 222944
rect 310532 16574 310560 228482
rect 311360 223310 311388 311866
rect 311348 223304 311400 223310
rect 311348 223246 311400 223252
rect 311452 221649 311480 319620
rect 311544 316130 311572 319790
rect 311774 319716 311802 320076
rect 311866 319870 311894 320076
rect 311854 319864 311906 319870
rect 311854 319806 311906 319812
rect 312050 319716 312078 320076
rect 312142 319784 312170 320076
rect 312326 319938 312354 320076
rect 315808 320104 315864 320113
rect 312496 320039 312552 320048
rect 312314 319932 312366 319938
rect 312314 319874 312366 319880
rect 312602 319870 312630 320076
rect 312694 319870 312722 320076
rect 312786 319870 312814 320076
rect 312878 319870 312906 320076
rect 313062 319938 313090 320076
rect 313050 319932 313102 319938
rect 313050 319874 313102 319880
rect 312590 319864 312642 319870
rect 312266 319832 312322 319841
rect 312590 319806 312642 319812
rect 312682 319864 312734 319870
rect 312682 319806 312734 319812
rect 312774 319864 312826 319870
rect 312774 319806 312826 319812
rect 312866 319864 312918 319870
rect 313338 319852 313366 320076
rect 313430 319938 313458 320076
rect 313418 319932 313470 319938
rect 313418 319874 313470 319880
rect 312866 319806 312918 319812
rect 313186 319832 313242 319841
rect 312142 319756 312216 319784
rect 312266 319767 312268 319776
rect 311774 319688 311848 319716
rect 312050 319688 312124 319716
rect 311624 319456 311676 319462
rect 311624 319398 311676 319404
rect 311532 316124 311584 316130
rect 311532 316066 311584 316072
rect 311532 315988 311584 315994
rect 311532 315930 311584 315936
rect 311544 311234 311572 315930
rect 311532 311228 311584 311234
rect 311532 311170 311584 311176
rect 311636 230314 311664 319398
rect 311716 319252 311768 319258
rect 311716 319194 311768 319200
rect 311728 317529 311756 319194
rect 311820 318306 311848 319688
rect 311900 319592 311952 319598
rect 311900 319534 311952 319540
rect 311912 319258 311940 319534
rect 311900 319252 311952 319258
rect 311900 319194 311952 319200
rect 311990 318880 312046 318889
rect 311990 318815 312046 318824
rect 311808 318300 311860 318306
rect 311808 318242 311860 318248
rect 311808 317960 311860 317966
rect 311808 317902 311860 317908
rect 311714 317520 311770 317529
rect 311714 317455 311770 317464
rect 311716 316124 311768 316130
rect 311716 316066 311768 316072
rect 311728 314809 311756 316066
rect 311714 314800 311770 314809
rect 311714 314735 311770 314744
rect 311820 234190 311848 317902
rect 312004 315654 312032 318815
rect 312096 318646 312124 319688
rect 312084 318640 312136 318646
rect 312084 318582 312136 318588
rect 312084 315988 312136 315994
rect 312084 315930 312136 315936
rect 311992 315648 312044 315654
rect 311992 315590 312044 315596
rect 312096 263634 312124 315930
rect 312188 294030 312216 319756
rect 312320 319767 312322 319776
rect 313186 319767 313242 319776
rect 313292 319824 313366 319852
rect 312268 319738 312320 319744
rect 312544 319728 312596 319734
rect 312544 319670 312596 319676
rect 312634 319696 312690 319705
rect 312360 319660 312412 319666
rect 312360 319602 312412 319608
rect 312268 319456 312320 319462
rect 312268 319398 312320 319404
rect 312280 317898 312308 319398
rect 312268 317892 312320 317898
rect 312268 317834 312320 317840
rect 312372 315874 312400 319602
rect 312450 319560 312506 319569
rect 312450 319495 312506 319504
rect 312464 315994 312492 319495
rect 312556 318034 312584 319670
rect 312634 319631 312690 319640
rect 312728 319660 312780 319666
rect 312648 319462 312676 319631
rect 312728 319602 312780 319608
rect 313096 319660 313148 319666
rect 313096 319602 313148 319608
rect 312636 319456 312688 319462
rect 312636 319398 312688 319404
rect 312634 319016 312690 319025
rect 312634 318951 312690 318960
rect 312544 318028 312596 318034
rect 312544 317970 312596 317976
rect 312452 315988 312504 315994
rect 312452 315930 312504 315936
rect 312372 315858 312492 315874
rect 312372 315852 312504 315858
rect 312372 315846 312452 315852
rect 312452 315794 312504 315800
rect 312360 315784 312412 315790
rect 312360 315726 312412 315732
rect 312372 310622 312400 315726
rect 312648 314770 312676 318951
rect 312740 315994 312768 319602
rect 312820 319592 312872 319598
rect 312820 319534 312872 319540
rect 313002 319560 313058 319569
rect 312728 315988 312780 315994
rect 312728 315930 312780 315936
rect 312728 315852 312780 315858
rect 312728 315794 312780 315800
rect 312636 314764 312688 314770
rect 312636 314706 312688 314712
rect 312648 311894 312676 314706
rect 312556 311866 312676 311894
rect 312360 310616 312412 310622
rect 312360 310558 312412 310564
rect 312176 294024 312228 294030
rect 312176 293966 312228 293972
rect 312084 263628 312136 263634
rect 312084 263570 312136 263576
rect 311808 234184 311860 234190
rect 311808 234126 311860 234132
rect 311624 230308 311676 230314
rect 311624 230250 311676 230256
rect 312556 225826 312584 311866
rect 312636 310616 312688 310622
rect 312636 310558 312688 310564
rect 312648 233889 312676 310558
rect 312740 309505 312768 315794
rect 312832 313070 312860 319534
rect 313002 319495 313058 319504
rect 312912 319456 312964 319462
rect 312912 319398 312964 319404
rect 312924 315625 312952 319398
rect 313016 318345 313044 319495
rect 313002 318336 313058 318345
rect 313002 318271 313058 318280
rect 313004 315988 313056 315994
rect 313004 315930 313056 315936
rect 312910 315616 312966 315625
rect 312910 315551 312966 315560
rect 312820 313064 312872 313070
rect 312820 313006 312872 313012
rect 312726 309496 312782 309505
rect 312726 309431 312782 309440
rect 312728 294024 312780 294030
rect 312728 293966 312780 293972
rect 312634 233880 312690 233889
rect 312634 233815 312690 233824
rect 312740 227322 312768 293966
rect 313016 258074 313044 315930
rect 312832 258046 313044 258074
rect 312832 248470 312860 258046
rect 312912 250504 312964 250510
rect 312912 250446 312964 250452
rect 312820 248464 312872 248470
rect 312820 248406 312872 248412
rect 312728 227316 312780 227322
rect 312728 227258 312780 227264
rect 312832 226166 312860 248406
rect 312924 227118 312952 250446
rect 313108 228682 313136 319602
rect 313200 315790 313228 319767
rect 313292 319705 313320 319824
rect 313522 319784 313550 320076
rect 313384 319756 313550 319784
rect 313278 319696 313334 319705
rect 313278 319631 313334 319640
rect 313280 319456 313332 319462
rect 313280 319398 313332 319404
rect 313292 317558 313320 319398
rect 313384 318034 313412 319756
rect 313614 319716 313642 320076
rect 313706 319784 313734 320076
rect 313798 319938 313826 320076
rect 313786 319932 313838 319938
rect 313786 319874 313838 319880
rect 313890 319870 313918 320076
rect 313878 319864 313930 319870
rect 313878 319806 313930 319812
rect 313706 319756 313780 319784
rect 313462 319696 313518 319705
rect 313614 319688 313688 319716
rect 313462 319631 313518 319640
rect 313476 319546 313504 319631
rect 313476 319518 313596 319546
rect 313464 319456 313516 319462
rect 313464 319398 313516 319404
rect 313372 318028 313424 318034
rect 313372 317970 313424 317976
rect 313280 317552 313332 317558
rect 313280 317494 313332 317500
rect 313476 315976 313504 319398
rect 313384 315948 313504 315976
rect 313188 315784 313240 315790
rect 313188 315726 313240 315732
rect 313188 315648 313240 315654
rect 313188 315590 313240 315596
rect 313200 300257 313228 315590
rect 313280 313268 313332 313274
rect 313280 313210 313332 313216
rect 313292 311914 313320 313210
rect 313280 311908 313332 311914
rect 313280 311850 313332 311856
rect 313292 307222 313320 311850
rect 313280 307216 313332 307222
rect 313280 307158 313332 307164
rect 313186 300248 313242 300257
rect 313186 300183 313242 300192
rect 313384 259418 313412 315948
rect 313464 315852 313516 315858
rect 313464 315794 313516 315800
rect 313476 269074 313504 315794
rect 313568 294545 313596 319518
rect 313660 315994 313688 319688
rect 313752 316878 313780 319756
rect 313830 319696 313886 319705
rect 313830 319631 313886 319640
rect 313982 319648 314010 320076
rect 314074 319870 314102 320076
rect 314062 319864 314114 319870
rect 314062 319806 314114 319812
rect 314166 319716 314194 320076
rect 314258 319852 314286 320076
rect 314442 319954 314470 320076
rect 314396 319926 314470 319954
rect 314258 319824 314332 319852
rect 314120 319688 314194 319716
rect 313740 316872 313792 316878
rect 313740 316814 313792 316820
rect 313648 315988 313700 315994
rect 313648 315930 313700 315936
rect 313844 313274 313872 319631
rect 313982 319620 314056 319648
rect 313924 319524 313976 319530
rect 313924 319466 313976 319472
rect 313936 314702 313964 319466
rect 314028 317966 314056 319620
rect 314016 317960 314068 317966
rect 314016 317902 314068 317908
rect 314120 315858 314148 319688
rect 314200 319592 314252 319598
rect 314200 319534 314252 319540
rect 314108 315852 314160 315858
rect 314108 315794 314160 315800
rect 314106 315072 314162 315081
rect 314106 315007 314162 315016
rect 313924 314696 313976 314702
rect 313924 314638 313976 314644
rect 313832 313268 313884 313274
rect 313832 313210 313884 313216
rect 313936 311894 313964 314638
rect 314120 313342 314148 315007
rect 314108 313336 314160 313342
rect 314108 313278 314160 313284
rect 313936 311866 314056 311894
rect 313924 308440 313976 308446
rect 313924 308382 313976 308388
rect 313554 294536 313610 294545
rect 313554 294471 313610 294480
rect 313464 269068 313516 269074
rect 313464 269010 313516 269016
rect 313464 263628 313516 263634
rect 313464 263570 313516 263576
rect 313372 259412 313424 259418
rect 313372 259354 313424 259360
rect 313476 239018 313504 263570
rect 313936 241058 313964 308382
rect 313924 241052 313976 241058
rect 313924 240994 313976 241000
rect 313464 239012 313516 239018
rect 313464 238954 313516 238960
rect 313924 233980 313976 233986
rect 313924 233922 313976 233928
rect 313096 228676 313148 228682
rect 313096 228618 313148 228624
rect 313108 228410 313136 228618
rect 313096 228404 313148 228410
rect 313096 228346 313148 228352
rect 312912 227112 312964 227118
rect 312912 227054 312964 227060
rect 312820 226160 312872 226166
rect 312820 226102 312872 226108
rect 312544 225820 312596 225826
rect 312544 225762 312596 225768
rect 313278 223000 313334 223009
rect 313278 222935 313280 222944
rect 313332 222935 313334 222944
rect 313280 222906 313332 222912
rect 313280 221944 313332 221950
rect 313280 221886 313332 221892
rect 311438 221640 311494 221649
rect 311438 221575 311494 221584
rect 313292 221542 313320 221886
rect 313280 221536 313332 221542
rect 313280 221478 313332 221484
rect 311162 192536 311218 192545
rect 311162 192471 311218 192480
rect 310532 16546 311112 16574
rect 311084 3482 311112 16546
rect 311176 3602 311204 192471
rect 313936 3670 313964 233922
rect 314028 226030 314056 311866
rect 314120 311166 314148 313278
rect 314108 311160 314160 311166
rect 314108 311102 314160 311108
rect 314212 310185 314240 319534
rect 314304 319054 314332 319824
rect 314292 319048 314344 319054
rect 314292 318990 314344 318996
rect 314396 317529 314424 319926
rect 314534 319852 314562 320076
rect 314488 319824 314562 319852
rect 314382 317520 314438 317529
rect 314382 317455 314438 317464
rect 314292 315988 314344 315994
rect 314292 315930 314344 315936
rect 314198 310176 314254 310185
rect 314198 310111 314254 310120
rect 314304 310049 314332 315930
rect 314290 310040 314346 310049
rect 314290 309975 314346 309984
rect 314108 304292 314160 304298
rect 314108 304234 314160 304240
rect 314120 232529 314148 304234
rect 314200 269068 314252 269074
rect 314200 269010 314252 269016
rect 314212 267782 314240 269010
rect 314200 267776 314252 267782
rect 314200 267718 314252 267724
rect 314212 239290 314240 267718
rect 314384 259412 314436 259418
rect 314384 259354 314436 259360
rect 314396 258194 314424 259354
rect 314384 258188 314436 258194
rect 314384 258130 314436 258136
rect 314292 249076 314344 249082
rect 314292 249018 314344 249024
rect 314200 239284 314252 239290
rect 314200 239226 314252 239232
rect 314106 232520 314162 232529
rect 314106 232455 314162 232464
rect 314016 226024 314068 226030
rect 314016 225966 314068 225972
rect 314304 225350 314332 249018
rect 314396 239086 314424 258130
rect 314384 239080 314436 239086
rect 314384 239022 314436 239028
rect 314292 225344 314344 225350
rect 314292 225286 314344 225292
rect 314488 221542 314516 319824
rect 314626 319784 314654 320076
rect 314718 319818 314746 320076
rect 314810 319938 314838 320076
rect 314798 319932 314850 319938
rect 314798 319874 314850 319880
rect 314902 319852 314930 320076
rect 314994 319954 315022 320076
rect 315178 319954 315206 320076
rect 314994 319926 315068 319954
rect 314902 319824 314976 319852
rect 314718 319790 314792 319818
rect 314580 319756 314654 319784
rect 314764 319784 314792 319790
rect 314764 319756 314884 319784
rect 314580 317801 314608 319756
rect 314750 319696 314806 319705
rect 314750 319631 314806 319640
rect 314660 319388 314712 319394
rect 314660 319330 314712 319336
rect 314672 319297 314700 319330
rect 314658 319288 314714 319297
rect 314658 319223 314714 319232
rect 314566 317792 314622 317801
rect 314566 317727 314622 317736
rect 314568 317484 314620 317490
rect 314568 317426 314620 317432
rect 314580 253978 314608 317426
rect 314764 310214 314792 319631
rect 314856 315586 314884 319756
rect 314844 315580 314896 315586
rect 314844 315522 314896 315528
rect 314752 310208 314804 310214
rect 314752 310150 314804 310156
rect 314948 308446 314976 319824
rect 315040 312730 315068 319926
rect 315132 319926 315206 319954
rect 315132 317490 315160 319926
rect 315270 319784 315298 320076
rect 315224 319756 315298 319784
rect 315362 319784 315390 320076
rect 315454 319938 315482 320076
rect 315442 319932 315494 319938
rect 315442 319874 315494 319880
rect 315546 319784 315574 320076
rect 315638 319938 315666 320076
rect 315626 319932 315678 319938
rect 315626 319874 315678 319880
rect 315730 319784 315758 320076
rect 315992 320104 316048 320113
rect 315808 320039 315864 320048
rect 315914 319784 315942 320076
rect 316176 320104 316232 320113
rect 315992 320039 316048 320048
rect 316098 319954 316126 320076
rect 317188 320104 317244 320113
rect 316176 320039 316232 320048
rect 316374 319954 316402 320076
rect 316098 319926 316172 319954
rect 315362 319756 315436 319784
rect 315546 319756 315620 319784
rect 315730 319756 315804 319784
rect 315120 317484 315172 317490
rect 315120 317426 315172 317432
rect 315224 315858 315252 319756
rect 315304 319660 315356 319666
rect 315304 319602 315356 319608
rect 315212 315852 315264 315858
rect 315212 315794 315264 315800
rect 315316 313410 315344 319602
rect 315408 315994 315436 319756
rect 315488 316124 315540 316130
rect 315488 316066 315540 316072
rect 315396 315988 315448 315994
rect 315396 315930 315448 315936
rect 315500 315058 315528 316066
rect 315592 315976 315620 319756
rect 315672 319660 315724 319666
rect 315672 319602 315724 319608
rect 315684 317490 315712 319602
rect 315672 317484 315724 317490
rect 315672 317426 315724 317432
rect 315776 316130 315804 319756
rect 315868 319756 315942 319784
rect 315764 316124 315816 316130
rect 315764 316066 315816 316072
rect 315764 315988 315816 315994
rect 315592 315948 315712 315976
rect 315580 315852 315632 315858
rect 315580 315794 315632 315800
rect 315408 315030 315528 315058
rect 315304 313404 315356 313410
rect 315304 313346 315356 313352
rect 315028 312724 315080 312730
rect 315028 312666 315080 312672
rect 314936 308440 314988 308446
rect 314936 308382 314988 308388
rect 314568 253972 314620 253978
rect 314568 253914 314620 253920
rect 314844 253972 314896 253978
rect 314844 253914 314896 253920
rect 314856 225622 314884 253914
rect 314936 240100 314988 240106
rect 314936 240042 314988 240048
rect 314948 229094 314976 240042
rect 315316 232937 315344 313346
rect 315408 313342 315436 315030
rect 315488 313812 315540 313818
rect 315488 313754 315540 313760
rect 315396 313336 315448 313342
rect 315396 313278 315448 313284
rect 315408 237522 315436 313278
rect 315500 237862 315528 313754
rect 315592 310321 315620 315794
rect 315578 310312 315634 310321
rect 315578 310247 315634 310256
rect 315580 309800 315632 309806
rect 315580 309742 315632 309748
rect 315592 238105 315620 309742
rect 315684 307290 315712 315948
rect 315764 315930 315816 315936
rect 315672 307284 315724 307290
rect 315672 307226 315724 307232
rect 315578 238096 315634 238105
rect 315578 238031 315634 238040
rect 315488 237856 315540 237862
rect 315488 237798 315540 237804
rect 315396 237516 315448 237522
rect 315396 237458 315448 237464
rect 315302 232928 315358 232937
rect 315302 232863 315358 232872
rect 315776 231130 315804 315930
rect 315764 231124 315816 231130
rect 315764 231066 315816 231072
rect 314948 229066 315344 229094
rect 314948 228886 314976 229066
rect 314936 228880 314988 228886
rect 314936 228822 314988 228828
rect 314844 225616 314896 225622
rect 314844 225558 314896 225564
rect 314476 221536 314528 221542
rect 314476 221478 314528 221484
rect 315316 4146 315344 229066
rect 315868 220522 315896 319756
rect 316040 319660 316092 319666
rect 316040 319602 316092 319608
rect 315946 319560 316002 319569
rect 315946 319495 316002 319504
rect 315960 314362 315988 319495
rect 316052 319326 316080 319602
rect 316040 319320 316092 319326
rect 316040 319262 316092 319268
rect 315948 314356 316000 314362
rect 315948 314298 316000 314304
rect 316144 310078 316172 319926
rect 316328 319926 316402 319954
rect 316466 319954 316494 320076
rect 316466 319926 316540 319954
rect 316224 319728 316276 319734
rect 316328 319705 316356 319926
rect 316408 319864 316460 319870
rect 316408 319806 316460 319812
rect 316224 319670 316276 319676
rect 316314 319696 316370 319705
rect 316132 310072 316184 310078
rect 316132 310014 316184 310020
rect 316236 247178 316264 319670
rect 316314 319631 316370 319640
rect 316314 319016 316370 319025
rect 316314 318951 316370 318960
rect 316328 262682 316356 318951
rect 316420 287745 316448 319806
rect 316512 319648 316540 319926
rect 316650 319870 316678 320076
rect 316638 319864 316690 319870
rect 316638 319806 316690 319812
rect 316742 319716 316770 320076
rect 316834 319818 316862 320076
rect 316926 319938 316954 320076
rect 317018 319938 317046 320076
rect 317464 320104 317520 320113
rect 317188 320039 317244 320048
rect 316914 319932 316966 319938
rect 316914 319874 316966 319880
rect 317006 319932 317058 319938
rect 317006 319874 317058 319880
rect 317386 319852 317414 320076
rect 318108 320104 318164 320113
rect 317464 320039 317520 320048
rect 317050 319832 317106 319841
rect 316834 319790 316954 319818
rect 316926 319784 316954 319790
rect 316926 319756 317000 319784
rect 317386 319824 317460 319852
rect 317050 319767 317106 319776
rect 317144 319796 317196 319802
rect 316696 319688 316770 319716
rect 316512 319620 316632 319648
rect 316498 319560 316554 319569
rect 316498 319495 316554 319504
rect 316512 319462 316540 319495
rect 316500 319456 316552 319462
rect 316500 319398 316552 319404
rect 316604 318170 316632 319620
rect 316592 318164 316644 318170
rect 316592 318106 316644 318112
rect 316696 316878 316724 319688
rect 316774 319560 316830 319569
rect 316774 319495 316830 319504
rect 316684 316872 316736 316878
rect 316684 316814 316736 316820
rect 316788 315518 316816 319495
rect 316776 315512 316828 315518
rect 316776 315454 316828 315460
rect 316972 313954 317000 319756
rect 316960 313948 317012 313954
rect 316960 313890 317012 313896
rect 316972 313818 317000 313890
rect 316960 313812 317012 313818
rect 316960 313754 317012 313760
rect 316684 297424 316736 297430
rect 316684 297366 316736 297372
rect 316406 287736 316462 287745
rect 316406 287671 316462 287680
rect 316316 262676 316368 262682
rect 316316 262618 316368 262624
rect 316224 247172 316276 247178
rect 316224 247114 316276 247120
rect 316236 240854 316264 247114
rect 316224 240848 316276 240854
rect 316224 240790 316276 240796
rect 316696 235793 316724 297366
rect 316776 262676 316828 262682
rect 316776 262618 316828 262624
rect 316788 262274 316816 262618
rect 316776 262268 316828 262274
rect 316776 262210 316828 262216
rect 316682 235784 316738 235793
rect 316682 235719 316738 235728
rect 316788 224466 316816 262210
rect 316776 224460 316828 224466
rect 316776 224402 316828 224408
rect 317064 222970 317092 319767
rect 317144 319738 317196 319744
rect 317156 225962 317184 319738
rect 317234 319560 317290 319569
rect 317234 319495 317290 319504
rect 317248 310146 317276 319495
rect 317326 318608 317382 318617
rect 317326 318543 317328 318552
rect 317380 318543 317382 318552
rect 317328 318514 317380 318520
rect 317432 318442 317460 319824
rect 317570 319818 317598 320076
rect 317754 319943 317782 320076
rect 317740 319934 317796 319943
rect 317740 319869 317796 319878
rect 317570 319790 317736 319818
rect 317602 319696 317658 319705
rect 317602 319631 317658 319640
rect 317420 318436 317472 318442
rect 317420 318378 317472 318384
rect 317236 310140 317288 310146
rect 317236 310082 317288 310088
rect 317616 290465 317644 319631
rect 317708 317082 317736 319790
rect 317846 319716 317874 320076
rect 317800 319688 317874 319716
rect 317938 319716 317966 320076
rect 318030 319784 318058 320076
rect 318568 320104 318624 320113
rect 318108 320039 318164 320048
rect 318214 319870 318242 320076
rect 318202 319864 318254 319870
rect 318306 319852 318334 320076
rect 318490 319852 318518 320076
rect 319212 320104 319268 320113
rect 318568 320039 318624 320048
rect 318674 319920 318702 320076
rect 318674 319892 318840 319920
rect 318306 319824 318380 319852
rect 318490 319824 318656 319852
rect 318202 319806 318254 319812
rect 318030 319756 318104 319784
rect 317938 319688 318012 319716
rect 318076 319705 318104 319756
rect 317696 317076 317748 317082
rect 317696 317018 317748 317024
rect 317800 315722 317828 319688
rect 317878 319560 317934 319569
rect 317878 319495 317934 319504
rect 317788 315716 317840 315722
rect 317788 315658 317840 315664
rect 317892 311894 317920 319495
rect 317984 318510 318012 319688
rect 318062 319696 318118 319705
rect 318062 319631 318118 319640
rect 318062 319424 318118 319433
rect 318062 319359 318118 319368
rect 317972 318504 318024 318510
rect 317972 318446 318024 318452
rect 317972 317484 318024 317490
rect 317972 317426 318024 317432
rect 317708 311866 317920 311894
rect 317708 308553 317736 311866
rect 317694 308544 317750 308553
rect 317694 308479 317750 308488
rect 317602 290456 317658 290465
rect 317602 290391 317658 290400
rect 317144 225956 317196 225962
rect 317144 225898 317196 225904
rect 317328 225956 317380 225962
rect 317328 225898 317380 225904
rect 317340 225622 317368 225898
rect 317328 225616 317380 225622
rect 317328 225558 317380 225564
rect 317984 225554 318012 317426
rect 318076 313002 318104 319359
rect 318248 318912 318300 318918
rect 318248 318854 318300 318860
rect 318064 312996 318116 313002
rect 318064 312938 318116 312944
rect 318260 310010 318288 318854
rect 318352 317529 318380 319824
rect 318430 319696 318486 319705
rect 318430 319631 318486 319640
rect 318444 318918 318472 319631
rect 318522 319424 318578 319433
rect 318522 319359 318578 319368
rect 318432 318912 318484 318918
rect 318432 318854 318484 318860
rect 318432 318776 318484 318782
rect 318432 318718 318484 318724
rect 318338 317520 318394 317529
rect 318338 317455 318394 317464
rect 318248 310004 318300 310010
rect 318248 309946 318300 309952
rect 318064 294636 318116 294642
rect 318064 294578 318116 294584
rect 317972 225548 318024 225554
rect 317972 225490 318024 225496
rect 318076 224641 318104 294578
rect 318248 291916 318300 291922
rect 318248 291858 318300 291864
rect 318062 224632 318118 224641
rect 318062 224567 318118 224576
rect 318260 224369 318288 291858
rect 318246 224360 318302 224369
rect 318246 224295 318302 224304
rect 317052 222964 317104 222970
rect 317052 222906 317104 222912
rect 315856 220516 315908 220522
rect 315856 220458 315908 220464
rect 315868 216034 315896 220458
rect 315856 216028 315908 216034
rect 315856 215970 315908 215976
rect 318444 212430 318472 318718
rect 318536 227390 318564 319359
rect 318628 318345 318656 319824
rect 318706 319696 318762 319705
rect 318706 319631 318762 319640
rect 318614 318336 318670 318345
rect 318614 318271 318670 318280
rect 318720 317422 318748 319631
rect 318812 318782 318840 319892
rect 318892 319864 318944 319870
rect 319042 319818 319070 320076
rect 319134 319852 319162 320076
rect 319396 320104 319452 320113
rect 319212 320039 319268 320048
rect 319318 319954 319346 320076
rect 319856 320104 319912 320113
rect 319396 320039 319452 320048
rect 319318 319926 319392 319954
rect 319260 319864 319312 319870
rect 319134 319824 319208 319852
rect 318892 319806 318944 319812
rect 318800 318776 318852 318782
rect 318800 318718 318852 318724
rect 318904 318374 318932 319806
rect 318996 319790 319070 319818
rect 318996 319648 319024 319790
rect 318996 319620 319116 319648
rect 318982 319560 319038 319569
rect 318982 319495 319038 319504
rect 318892 318368 318944 318374
rect 318892 318310 318944 318316
rect 318708 317416 318760 317422
rect 318708 317358 318760 317364
rect 318800 316056 318852 316062
rect 318800 315998 318852 316004
rect 318614 304056 318670 304065
rect 318614 303991 318670 304000
rect 318628 302938 318656 303991
rect 318616 302932 318668 302938
rect 318616 302874 318668 302880
rect 318524 227384 318576 227390
rect 318524 227326 318576 227332
rect 318536 227050 318564 227326
rect 318524 227044 318576 227050
rect 318524 226986 318576 226992
rect 318708 225548 318760 225554
rect 318708 225490 318760 225496
rect 318720 220182 318748 225490
rect 318708 220176 318760 220182
rect 318708 220118 318760 220124
rect 318432 212424 318484 212430
rect 318432 212366 318484 212372
rect 318708 212424 318760 212430
rect 318708 212366 318760 212372
rect 318720 211886 318748 212366
rect 318708 211880 318760 211886
rect 318708 211822 318760 211828
rect 318812 211002 318840 315998
rect 318996 311894 319024 319495
rect 319088 319444 319116 319620
rect 319180 319569 319208 319824
rect 319260 319806 319312 319812
rect 319166 319560 319222 319569
rect 319166 319495 319222 319504
rect 319088 319416 319208 319444
rect 319074 319016 319130 319025
rect 319074 318951 319130 318960
rect 318904 311866 319024 311894
rect 318904 309942 318932 311866
rect 318892 309936 318944 309942
rect 318892 309878 318944 309884
rect 319088 265878 319116 318951
rect 319180 318209 319208 319416
rect 319272 318481 319300 319806
rect 319258 318472 319314 318481
rect 319258 318407 319314 318416
rect 319166 318200 319222 318209
rect 319166 318135 319222 318144
rect 319168 315988 319220 315994
rect 319168 315930 319220 315936
rect 319180 306374 319208 315930
rect 319272 314294 319300 318407
rect 319364 318238 319392 319926
rect 319502 319784 319530 320076
rect 319594 319938 319622 320076
rect 319582 319932 319634 319938
rect 319582 319874 319634 319880
rect 319686 319841 319714 320076
rect 319778 319852 319806 320076
rect 320040 320104 320096 320113
rect 319856 320039 319912 320048
rect 319962 319920 319990 320076
rect 320408 320104 320464 320113
rect 320040 320039 320096 320048
rect 319962 319892 320128 319920
rect 319456 319756 319530 319784
rect 319672 319832 319728 319841
rect 319778 319824 319944 319852
rect 319672 319767 319728 319776
rect 319352 318232 319404 318238
rect 319352 318174 319404 318180
rect 319456 316062 319484 319756
rect 319534 319696 319590 319705
rect 319810 319696 319866 319705
rect 319534 319631 319590 319640
rect 319732 319654 319810 319682
rect 319444 316056 319496 316062
rect 319444 315998 319496 316004
rect 319260 314288 319312 314294
rect 319260 314230 319312 314236
rect 319548 311894 319576 319631
rect 319626 319424 319682 319433
rect 319626 319359 319682 319368
rect 319640 314090 319668 319359
rect 319732 315994 319760 319654
rect 319810 319631 319866 319640
rect 319810 319560 319866 319569
rect 319810 319495 319866 319504
rect 319824 316010 319852 319495
rect 319916 318782 319944 319824
rect 319994 319832 320050 319841
rect 319994 319767 320050 319776
rect 319904 318776 319956 318782
rect 319904 318718 319956 318724
rect 320008 318714 320036 319767
rect 319996 318708 320048 318714
rect 319996 318650 320048 318656
rect 319720 315988 319772 315994
rect 319824 315982 320036 316010
rect 319720 315930 319772 315936
rect 319628 314084 319680 314090
rect 319628 314026 319680 314032
rect 319548 311866 319944 311894
rect 319916 308417 319944 311866
rect 319902 308408 319958 308417
rect 319902 308343 319958 308352
rect 319180 306346 319484 306374
rect 319456 292602 319484 306346
rect 319444 292596 319496 292602
rect 319444 292538 319496 292544
rect 319076 265872 319128 265878
rect 319076 265814 319128 265820
rect 319456 237046 319484 292538
rect 319628 265872 319680 265878
rect 319628 265814 319680 265820
rect 319640 264994 319668 265814
rect 319628 264988 319680 264994
rect 319628 264930 319680 264936
rect 319536 255332 319588 255338
rect 319536 255274 319588 255280
rect 319444 237040 319496 237046
rect 319444 236982 319496 236988
rect 319444 226364 319496 226370
rect 319444 226306 319496 226312
rect 318800 210996 318852 211002
rect 318800 210938 318852 210944
rect 318064 210452 318116 210458
rect 318064 210394 318116 210400
rect 316130 152416 316186 152425
rect 316130 152351 316186 152360
rect 316144 16574 316172 152351
rect 316144 16546 316264 16574
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 313924 3664 313976 3670
rect 313924 3606 313976 3612
rect 311164 3596 311216 3602
rect 311164 3538 311216 3544
rect 312636 3596 312688 3602
rect 312636 3538 312688 3544
rect 311084 3454 311480 3482
rect 309876 3188 309928 3194
rect 309876 3130 309928 3136
rect 311452 480 311480 3454
rect 312648 480 312676 3538
rect 313832 3528 313884 3534
rect 313832 3470 313884 3476
rect 313844 480 313872 3470
rect 315028 3188 315080 3194
rect 315028 3130 315080 3136
rect 315040 480 315068 3130
rect 316236 480 316264 16546
rect 317328 3664 317380 3670
rect 317328 3606 317380 3612
rect 317340 480 317368 3606
rect 318076 3534 318104 210394
rect 318524 4140 318576 4146
rect 318524 4082 318576 4088
rect 318064 3528 318116 3534
rect 318064 3470 318116 3476
rect 318536 480 318564 4082
rect 319456 4010 319484 226306
rect 319548 224670 319576 255274
rect 319640 244089 319668 264930
rect 319626 244080 319682 244089
rect 319626 244015 319682 244024
rect 319536 224664 319588 224670
rect 319536 224606 319588 224612
rect 320008 219162 320036 315982
rect 320100 255338 320128 319892
rect 320238 319818 320266 320076
rect 320330 319870 320358 320076
rect 321144 320104 321200 320113
rect 320408 320039 320464 320048
rect 320192 319790 320266 319818
rect 320318 319864 320370 319870
rect 320318 319806 320370 319812
rect 320192 316062 320220 319790
rect 320514 319784 320542 320076
rect 320606 319870 320634 320076
rect 320698 319938 320726 320076
rect 320686 319932 320738 319938
rect 320686 319874 320738 319880
rect 320594 319864 320646 319870
rect 320594 319806 320646 319812
rect 320790 319784 320818 320076
rect 320882 320074 320910 320076
rect 320870 320068 320922 320074
rect 320870 320010 320922 320016
rect 320974 319954 321002 320076
rect 320468 319756 320542 319784
rect 320744 319756 320818 319784
rect 320928 319926 321002 319954
rect 320272 319728 320324 319734
rect 320272 319670 320324 319676
rect 320364 319728 320416 319734
rect 320364 319670 320416 319676
rect 320284 318918 320312 319670
rect 320272 318912 320324 318918
rect 320272 318854 320324 318860
rect 320180 316056 320232 316062
rect 320180 315998 320232 316004
rect 320088 255332 320140 255338
rect 320088 255274 320140 255280
rect 320376 245750 320404 319670
rect 320468 316674 320496 319756
rect 320638 319696 320694 319705
rect 320638 319631 320640 319640
rect 320692 319631 320694 319640
rect 320640 319602 320692 319608
rect 320638 319560 320694 319569
rect 320638 319495 320694 319504
rect 320652 316849 320680 319495
rect 320744 317694 320772 319756
rect 320732 317688 320784 317694
rect 320732 317630 320784 317636
rect 320732 317552 320784 317558
rect 320732 317494 320784 317500
rect 320638 316840 320694 316849
rect 320638 316775 320694 316784
rect 320456 316668 320508 316674
rect 320456 316610 320508 316616
rect 320640 316056 320692 316062
rect 320640 315998 320692 316004
rect 320456 315988 320508 315994
rect 320456 315930 320508 315936
rect 320468 259418 320496 315930
rect 320548 315852 320600 315858
rect 320548 315794 320600 315800
rect 320560 271862 320588 315794
rect 320652 290873 320680 315998
rect 320638 290864 320694 290873
rect 320638 290799 320694 290808
rect 320548 271856 320600 271862
rect 320548 271798 320600 271804
rect 320548 260160 320600 260166
rect 320548 260102 320600 260108
rect 320456 259412 320508 259418
rect 320456 259354 320508 259360
rect 320364 245744 320416 245750
rect 320364 245686 320416 245692
rect 320180 231192 320232 231198
rect 320180 231134 320232 231140
rect 319996 219156 320048 219162
rect 319996 219098 320048 219104
rect 320088 210996 320140 211002
rect 320088 210938 320140 210944
rect 320100 210458 320128 210938
rect 320088 210452 320140 210458
rect 320088 210394 320140 210400
rect 320192 16574 320220 231134
rect 320560 228954 320588 260102
rect 320548 228948 320600 228954
rect 320548 228890 320600 228896
rect 320560 227798 320588 228890
rect 320548 227792 320600 227798
rect 320548 227734 320600 227740
rect 320744 213926 320772 317494
rect 320928 314430 320956 319926
rect 321066 319852 321094 320076
rect 321512 320104 321568 320113
rect 321144 320039 321200 320048
rect 321020 319824 321094 319852
rect 321020 315994 321048 319824
rect 321250 319784 321278 320076
rect 321204 319756 321278 319784
rect 321342 319784 321370 320076
rect 321698 320078 321750 320084
rect 322156 320104 322212 320113
rect 321710 320076 321738 320078
rect 321512 320039 321568 320048
rect 321618 319784 321646 320076
rect 321342 319756 321508 319784
rect 321618 319756 321692 319784
rect 321098 319560 321154 319569
rect 321098 319495 321154 319504
rect 321008 315988 321060 315994
rect 321008 315930 321060 315936
rect 320916 314424 320968 314430
rect 320916 314366 320968 314372
rect 321112 312866 321140 319495
rect 321204 315858 321232 319756
rect 321282 319696 321338 319705
rect 321282 319631 321338 319640
rect 321296 319258 321324 319631
rect 321284 319252 321336 319258
rect 321284 319194 321336 319200
rect 321376 317688 321428 317694
rect 321376 317630 321428 317636
rect 321192 315852 321244 315858
rect 321192 315794 321244 315800
rect 321100 312860 321152 312866
rect 321100 312802 321152 312808
rect 321112 312730 321140 312802
rect 321100 312724 321152 312730
rect 321100 312666 321152 312672
rect 320916 312588 320968 312594
rect 320916 312530 320968 312536
rect 320824 311976 320876 311982
rect 320824 311918 320876 311924
rect 320836 232801 320864 311918
rect 320928 236745 320956 312530
rect 321100 271856 321152 271862
rect 321100 271798 321152 271804
rect 321112 270570 321140 271798
rect 321100 270564 321152 270570
rect 321100 270506 321152 270512
rect 321008 259412 321060 259418
rect 321008 259354 321060 259360
rect 321020 258126 321048 259354
rect 321008 258120 321060 258126
rect 321008 258062 321060 258068
rect 320914 236736 320970 236745
rect 320914 236671 320970 236680
rect 320822 232792 320878 232801
rect 320822 232727 320878 232736
rect 320824 227792 320876 227798
rect 320824 227734 320876 227740
rect 320732 213920 320784 213926
rect 320732 213862 320784 213868
rect 320744 213314 320772 213862
rect 320732 213308 320784 213314
rect 320732 213250 320784 213256
rect 320192 16546 320496 16574
rect 319444 4004 319496 4010
rect 319444 3946 319496 3952
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 319732 480 319760 3470
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 320836 3534 320864 227734
rect 321020 224738 321048 258062
rect 321112 239494 321140 270506
rect 321284 245744 321336 245750
rect 321284 245686 321336 245692
rect 321192 245676 321244 245682
rect 321192 245618 321244 245624
rect 321100 239488 321152 239494
rect 321100 239430 321152 239436
rect 321204 226098 321232 245618
rect 321296 237250 321324 245686
rect 321388 242962 321416 317630
rect 321480 245682 321508 319756
rect 321664 316062 321692 319756
rect 321802 319716 321830 320076
rect 321894 319784 321922 320076
rect 321986 319920 322014 320076
rect 322616 320104 322672 320113
rect 322156 320039 322212 320048
rect 322262 319943 322290 320076
rect 322248 319934 322304 319943
rect 321986 319892 322106 319920
rect 322078 319818 322106 319892
rect 322248 319869 322304 319878
rect 322078 319790 322244 319818
rect 321894 319756 321968 319784
rect 321802 319688 321876 319716
rect 321652 316056 321704 316062
rect 321652 315998 321704 316004
rect 321560 315988 321612 315994
rect 321560 315930 321612 315936
rect 321572 307154 321600 315930
rect 321744 315920 321796 315926
rect 321744 315862 321796 315868
rect 321560 307148 321612 307154
rect 321560 307090 321612 307096
rect 321756 247926 321784 315862
rect 321848 252550 321876 319688
rect 321940 315926 321968 319756
rect 322110 319696 322166 319705
rect 322110 319631 322166 319640
rect 322018 319560 322074 319569
rect 322124 319530 322152 319631
rect 322018 319495 322074 319504
rect 322112 319524 322164 319530
rect 321928 315920 321980 315926
rect 321928 315862 321980 315868
rect 322032 311894 322060 319495
rect 322112 319466 322164 319472
rect 322216 318850 322244 319790
rect 322354 319716 322382 320076
rect 322308 319688 322382 319716
rect 322446 319716 322474 320076
rect 322538 319818 322566 320076
rect 323628 320104 323684 320113
rect 322616 320039 322672 320048
rect 322722 319920 322750 320076
rect 322722 319892 322796 319920
rect 322662 319832 322718 319841
rect 322538 319790 322612 319818
rect 322446 319688 322520 319716
rect 322204 318844 322256 318850
rect 322204 318786 322256 318792
rect 322204 316260 322256 316266
rect 322204 316202 322256 316208
rect 321940 311866 322060 311894
rect 321940 252618 321968 311866
rect 321928 252612 321980 252618
rect 321928 252554 321980 252560
rect 321836 252544 321888 252550
rect 321836 252486 321888 252492
rect 321744 247920 321796 247926
rect 321744 247862 321796 247868
rect 321468 245676 321520 245682
rect 321468 245618 321520 245624
rect 321376 242956 321428 242962
rect 321376 242898 321428 242904
rect 321388 242049 321416 242898
rect 321374 242040 321430 242049
rect 321374 241975 321430 241984
rect 322216 239329 322244 316202
rect 322308 312662 322336 319688
rect 322386 319560 322442 319569
rect 322386 319495 322442 319504
rect 322400 319394 322428 319495
rect 322388 319388 322440 319394
rect 322388 319330 322440 319336
rect 322388 317960 322440 317966
rect 322492 317937 322520 319688
rect 322584 318986 322612 319790
rect 322662 319767 322718 319776
rect 322572 318980 322624 318986
rect 322572 318922 322624 318928
rect 322388 317902 322440 317908
rect 322478 317928 322534 317937
rect 322296 312656 322348 312662
rect 322296 312598 322348 312604
rect 322308 311982 322336 312598
rect 322296 311976 322348 311982
rect 322296 311918 322348 311924
rect 322296 252612 322348 252618
rect 322296 252554 322348 252560
rect 322202 239320 322258 239329
rect 322202 239255 322258 239264
rect 321560 239216 321612 239222
rect 321560 239158 321612 239164
rect 321284 237244 321336 237250
rect 321284 237186 321336 237192
rect 321192 226092 321244 226098
rect 321192 226034 321244 226040
rect 321008 224732 321060 224738
rect 321008 224674 321060 224680
rect 321572 16574 321600 239158
rect 322308 227497 322336 252554
rect 322400 249082 322428 317902
rect 322478 317863 322534 317872
rect 322480 316056 322532 316062
rect 322480 315998 322532 316004
rect 322388 249076 322440 249082
rect 322388 249018 322440 249024
rect 322388 247920 322440 247926
rect 322388 247862 322440 247868
rect 322400 247110 322428 247862
rect 322388 247104 322440 247110
rect 322388 247046 322440 247052
rect 322294 227488 322350 227497
rect 322294 227423 322350 227432
rect 322400 226137 322428 247046
rect 322492 244322 322520 315998
rect 322572 252544 322624 252550
rect 322572 252486 322624 252492
rect 322584 251258 322612 252486
rect 322572 251252 322624 251258
rect 322572 251194 322624 251200
rect 322480 244316 322532 244322
rect 322480 244258 322532 244264
rect 322386 226128 322442 226137
rect 322386 226063 322442 226072
rect 322492 224806 322520 244258
rect 322584 239154 322612 251194
rect 322572 239148 322624 239154
rect 322572 239090 322624 239096
rect 322676 230217 322704 319767
rect 322768 315994 322796 319892
rect 322906 319818 322934 320076
rect 322860 319790 322934 319818
rect 322998 319818 323026 320076
rect 323274 319954 323302 320076
rect 323274 319926 323348 319954
rect 322998 319790 323164 319818
rect 322860 319682 322888 319790
rect 322860 319654 322980 319682
rect 322846 319560 322902 319569
rect 322846 319495 322902 319504
rect 322860 316062 322888 319495
rect 322952 317354 322980 319654
rect 323032 319524 323084 319530
rect 323032 319466 323084 319472
rect 322940 317348 322992 317354
rect 322940 317290 322992 317296
rect 322848 316056 322900 316062
rect 322848 315998 322900 316004
rect 322756 315988 322808 315994
rect 322756 315930 322808 315936
rect 323044 312594 323072 319466
rect 323032 312588 323084 312594
rect 323032 312530 323084 312536
rect 323136 243681 323164 319790
rect 323216 319796 323268 319802
rect 323216 319738 323268 319744
rect 323228 244905 323256 319738
rect 323320 315926 323348 319926
rect 323458 319784 323486 320076
rect 323550 319938 323578 320076
rect 324088 320104 324144 320113
rect 323628 320039 323684 320048
rect 323538 319932 323590 319938
rect 323538 319874 323590 319880
rect 323734 319784 323762 320076
rect 323458 319756 323532 319784
rect 323398 319560 323454 319569
rect 323504 319530 323532 319756
rect 323596 319756 323762 319784
rect 323826 319784 323854 320076
rect 324010 319852 324038 320076
rect 326388 320104 326444 320113
rect 324088 320039 324144 320048
rect 324194 319920 324222 320076
rect 324378 319954 324406 320076
rect 324332 319926 324406 319954
rect 324194 319892 324268 319920
rect 324010 319824 324176 319852
rect 323826 319756 323900 319784
rect 323398 319495 323454 319504
rect 323492 319524 323544 319530
rect 323412 317626 323440 319495
rect 323492 319466 323544 319472
rect 323492 318640 323544 318646
rect 323492 318582 323544 318588
rect 323400 317620 323452 317626
rect 323400 317562 323452 317568
rect 323400 317416 323452 317422
rect 323400 317358 323452 317364
rect 323308 315920 323360 315926
rect 323308 315862 323360 315868
rect 323214 244896 323270 244905
rect 323214 244831 323270 244840
rect 323122 243672 323178 243681
rect 323122 243607 323178 243616
rect 322662 230208 322718 230217
rect 322662 230143 322718 230152
rect 322480 224800 322532 224806
rect 322480 224742 322532 224748
rect 322940 223440 322992 223446
rect 322940 223382 322992 223388
rect 322952 223038 322980 223382
rect 322940 223032 322992 223038
rect 322940 222974 322992 222980
rect 323412 219366 323440 317358
rect 323504 238754 323532 318582
rect 323596 316742 323624 319756
rect 323674 319696 323730 319705
rect 323674 319631 323730 319640
rect 323584 316736 323636 316742
rect 323584 316678 323636 316684
rect 323596 316266 323624 316678
rect 323584 316260 323636 316266
rect 323584 316202 323636 316208
rect 323688 316169 323716 319631
rect 323872 316198 323900 319756
rect 323950 319424 324006 319433
rect 323950 319359 324006 319368
rect 323860 316192 323912 316198
rect 323674 316160 323730 316169
rect 323584 316124 323636 316130
rect 323860 316134 323912 316140
rect 323674 316095 323730 316104
rect 323584 316066 323636 316072
rect 323596 241233 323624 316066
rect 323688 244934 323716 316095
rect 323964 316010 323992 319359
rect 324148 318794 324176 319824
rect 324240 319297 324268 319892
rect 324226 319288 324282 319297
rect 324226 319223 324282 319232
rect 324056 318766 324176 318794
rect 324056 316266 324084 318766
rect 324044 316260 324096 316266
rect 324044 316202 324096 316208
rect 324056 316130 324084 316202
rect 324136 316192 324188 316198
rect 324136 316134 324188 316140
rect 324044 316124 324096 316130
rect 324044 316066 324096 316072
rect 323780 315982 323992 316010
rect 323676 244928 323728 244934
rect 323676 244870 323728 244876
rect 323582 241224 323638 241233
rect 323582 241159 323638 241168
rect 323504 238726 323624 238754
rect 323596 223038 323624 238726
rect 323584 223032 323636 223038
rect 323584 222974 323636 222980
rect 323780 221474 323808 315982
rect 323952 315920 324004 315926
rect 323952 315862 324004 315868
rect 323964 241913 323992 315862
rect 324148 246362 324176 316134
rect 324136 246356 324188 246362
rect 324136 246298 324188 246304
rect 324332 243953 324360 319926
rect 324562 319920 324590 320076
rect 324470 319892 324590 319920
rect 324470 319852 324498 319892
rect 324654 319852 324682 320076
rect 324424 319824 324498 319852
rect 324608 319824 324682 319852
rect 324424 317558 324452 319824
rect 324502 319696 324558 319705
rect 324502 319631 324558 319640
rect 324412 317552 324464 317558
rect 324412 317494 324464 317500
rect 324412 310548 324464 310554
rect 324412 310490 324464 310496
rect 324424 308514 324452 310490
rect 324412 308508 324464 308514
rect 324412 308450 324464 308456
rect 324318 243944 324374 243953
rect 324318 243879 324374 243888
rect 323950 241904 324006 241913
rect 323950 241839 324006 241848
rect 323768 221468 323820 221474
rect 323768 221410 323820 221416
rect 324516 219434 324544 319631
rect 324608 246265 324636 319824
rect 324746 319784 324774 320076
rect 324700 319756 324774 319784
rect 324700 319025 324728 319756
rect 324838 319682 324866 320076
rect 324930 319784 324958 320076
rect 324930 319756 325004 319784
rect 324792 319654 324866 319682
rect 324686 319016 324742 319025
rect 324686 318951 324742 318960
rect 324688 315988 324740 315994
rect 324688 315930 324740 315936
rect 324700 258777 324728 315930
rect 324792 310554 324820 319654
rect 324976 318730 325004 319756
rect 325114 319716 325142 320076
rect 325206 319943 325234 320076
rect 325192 319934 325248 319943
rect 325192 319869 325248 319878
rect 325298 319784 325326 320076
rect 325252 319756 325326 319784
rect 325114 319688 325188 319716
rect 324884 318702 325004 318730
rect 324884 315994 324912 318702
rect 324964 318640 325016 318646
rect 324964 318582 325016 318588
rect 324976 316334 325004 318582
rect 324964 316328 325016 316334
rect 324964 316270 325016 316276
rect 324872 315988 324924 315994
rect 324872 315930 324924 315936
rect 324780 310548 324832 310554
rect 324780 310490 324832 310496
rect 324686 258768 324742 258777
rect 324686 258703 324742 258712
rect 324594 246256 324650 246265
rect 324594 246191 324650 246200
rect 324976 237969 325004 316270
rect 325056 316192 325108 316198
rect 325056 316134 325108 316140
rect 325068 239193 325096 316134
rect 325160 316130 325188 319688
rect 325252 319433 325280 319756
rect 325390 319716 325418 320076
rect 325482 319920 325510 320076
rect 325666 319954 325694 320076
rect 325620 319926 325694 319954
rect 325482 319892 325556 319920
rect 325344 319688 325418 319716
rect 325238 319424 325294 319433
rect 325238 319359 325294 319368
rect 325344 319138 325372 319688
rect 325252 319110 325372 319138
rect 325252 316470 325280 319110
rect 325528 319054 325556 319892
rect 325332 319048 325384 319054
rect 325332 318990 325384 318996
rect 325516 319048 325568 319054
rect 325516 318990 325568 318996
rect 325240 316464 325292 316470
rect 325240 316406 325292 316412
rect 325252 316198 325280 316406
rect 325240 316192 325292 316198
rect 325240 316134 325292 316140
rect 325148 316124 325200 316130
rect 325148 316066 325200 316072
rect 325160 241097 325188 316066
rect 325146 241088 325202 241097
rect 325146 241023 325202 241032
rect 325054 239184 325110 239193
rect 325054 239119 325110 239128
rect 324962 237960 325018 237969
rect 324962 237895 325018 237904
rect 324596 231872 324648 231878
rect 324596 231814 324648 231820
rect 324332 219406 324544 219434
rect 323400 219360 323452 219366
rect 323400 219302 323452 219308
rect 323412 218822 323440 219302
rect 323400 218816 323452 218822
rect 323400 218758 323452 218764
rect 322940 217320 322992 217326
rect 322940 217262 322992 217268
rect 321572 16546 322152 16574
rect 320824 3528 320876 3534
rect 320824 3470 320876 3476
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 217262
rect 324332 215150 324360 219406
rect 324320 215144 324372 215150
rect 324320 215086 324372 215092
rect 324332 214606 324360 215086
rect 324320 214600 324372 214606
rect 324320 214542 324372 214548
rect 324608 6914 324636 231814
rect 325344 205562 325372 318990
rect 325620 318646 325648 319926
rect 325758 319784 325786 320076
rect 325712 319756 325786 319784
rect 325608 318640 325660 318646
rect 325608 318582 325660 318588
rect 325608 318504 325660 318510
rect 325608 318446 325660 318452
rect 325422 318336 325478 318345
rect 325422 318271 325478 318280
rect 325436 318073 325464 318271
rect 325422 318064 325478 318073
rect 325620 318034 325648 318446
rect 325422 317999 325478 318008
rect 325608 318028 325660 318034
rect 325608 317970 325660 317976
rect 325712 243574 325740 319756
rect 325850 319716 325878 320076
rect 325942 319784 325970 320076
rect 326034 319920 326062 320076
rect 326218 319920 326246 320076
rect 326034 319892 326108 319920
rect 325942 319756 326016 319784
rect 325804 319688 325878 319716
rect 325804 318510 325832 319688
rect 325884 319456 325936 319462
rect 325884 319398 325936 319404
rect 325792 318504 325844 318510
rect 325792 318446 325844 318452
rect 325792 315988 325844 315994
rect 325792 315930 325844 315936
rect 325804 243817 325832 315930
rect 325896 245041 325924 319398
rect 325988 317801 326016 319756
rect 326080 319462 326108 319892
rect 326172 319892 326246 319920
rect 326068 319456 326120 319462
rect 326068 319398 326120 319404
rect 326068 319048 326120 319054
rect 326068 318990 326120 318996
rect 325974 317792 326030 317801
rect 325974 317727 326030 317736
rect 326080 311894 326108 318990
rect 326172 317490 326200 319892
rect 326310 319784 326338 320076
rect 326940 320104 326996 320113
rect 326388 320039 326444 320048
rect 326264 319756 326338 319784
rect 326494 319784 326522 320076
rect 326586 319920 326614 320076
rect 326586 319892 326660 319920
rect 326494 319756 326568 319784
rect 326160 317484 326212 317490
rect 326160 317426 326212 317432
rect 326264 315994 326292 319756
rect 326344 318640 326396 318646
rect 326540 318617 326568 319756
rect 326632 319054 326660 319892
rect 326770 319648 326798 320076
rect 326862 319784 326890 320076
rect 326940 320039 326996 320048
rect 327046 319954 327074 320076
rect 327000 319926 327074 319954
rect 327000 319841 327028 319926
rect 326986 319832 327042 319841
rect 326862 319756 326936 319784
rect 327138 319818 327166 320076
rect 326986 319767 327042 319776
rect 327092 319790 327166 319818
rect 326770 319620 326844 319648
rect 326710 319560 326766 319569
rect 326710 319495 326766 319504
rect 326620 319048 326672 319054
rect 326620 318990 326672 318996
rect 326344 318582 326396 318588
rect 326526 318608 326582 318617
rect 326356 318306 326384 318582
rect 326526 318543 326582 318552
rect 326618 318472 326674 318481
rect 326528 318436 326580 318442
rect 326618 318407 326674 318416
rect 326528 318378 326580 318384
rect 326344 318300 326396 318306
rect 326344 318242 326396 318248
rect 326436 318232 326488 318238
rect 326436 318174 326488 318180
rect 326448 317966 326476 318174
rect 326540 318170 326568 318378
rect 326528 318164 326580 318170
rect 326528 318106 326580 318112
rect 326436 317960 326488 317966
rect 326436 317902 326488 317908
rect 326528 317892 326580 317898
rect 326528 317834 326580 317840
rect 326252 315988 326304 315994
rect 326252 315930 326304 315936
rect 326540 311894 326568 317834
rect 326632 317665 326660 318407
rect 326618 317656 326674 317665
rect 326618 317591 326674 317600
rect 326724 317642 326752 319495
rect 326816 318794 326844 319620
rect 326908 319444 326936 319756
rect 326908 319416 327028 319444
rect 326816 318766 326936 318794
rect 326802 317656 326858 317665
rect 326724 317614 326802 317642
rect 326724 311894 326752 317614
rect 326802 317591 326858 317600
rect 326908 317257 326936 318766
rect 326894 317248 326950 317257
rect 326894 317183 326950 317192
rect 326908 316713 326936 317183
rect 326894 316704 326950 316713
rect 326894 316639 326950 316648
rect 325988 311866 326108 311894
rect 326448 311866 326568 311894
rect 326632 311866 326752 311894
rect 325988 250481 326016 311866
rect 326448 250510 326476 311866
rect 326632 271153 326660 311866
rect 327000 272513 327028 319416
rect 327092 315994 327120 319790
rect 327230 319716 327258 320076
rect 327322 319784 327350 320076
rect 327428 320062 328040 320090
rect 327322 319756 327396 319784
rect 327184 319688 327258 319716
rect 327080 315988 327132 315994
rect 327080 315930 327132 315936
rect 326986 272504 327042 272513
rect 326986 272439 327042 272448
rect 326618 271144 326674 271153
rect 326618 271079 326674 271088
rect 326436 250504 326488 250510
rect 325974 250472 326030 250481
rect 326436 250446 326488 250452
rect 325974 250407 326030 250416
rect 325882 245032 325938 245041
rect 325882 244967 325938 244976
rect 325790 243808 325846 243817
rect 325790 243743 325846 243752
rect 325700 243568 325752 243574
rect 325700 243510 325752 243516
rect 327078 224224 327134 224233
rect 327078 224159 327134 224168
rect 324872 205556 324924 205562
rect 324872 205498 324924 205504
rect 325332 205556 325384 205562
rect 325332 205498 325384 205504
rect 324884 204950 324912 205498
rect 324872 204944 324924 204950
rect 324872 204886 324924 204892
rect 324962 199336 325018 199345
rect 324962 199271 325018 199280
rect 324424 6886 324636 6914
rect 324424 480 324452 6886
rect 324976 3398 325004 199271
rect 327092 16574 327120 224159
rect 327184 216578 327212 319688
rect 327262 318608 327318 318617
rect 327262 318543 327318 318552
rect 327276 316146 327304 318543
rect 327368 317529 327396 319756
rect 327722 317792 327778 317801
rect 327722 317727 327778 317736
rect 327632 317552 327684 317558
rect 327354 317520 327410 317529
rect 327632 317494 327684 317500
rect 327354 317455 327410 317464
rect 327540 317484 327592 317490
rect 327540 317426 327592 317432
rect 327276 316118 327396 316146
rect 327264 315988 327316 315994
rect 327264 315930 327316 315936
rect 327276 258913 327304 315930
rect 327368 309806 327396 316118
rect 327448 316056 327500 316062
rect 327448 315998 327500 316004
rect 327356 309800 327408 309806
rect 327356 309742 327408 309748
rect 327262 258904 327318 258913
rect 327262 258839 327318 258848
rect 327460 234161 327488 315998
rect 327552 304298 327580 317426
rect 327644 305658 327672 317494
rect 327736 309194 327764 317727
rect 327816 317620 327868 317626
rect 327816 317562 327868 317568
rect 327724 309188 327776 309194
rect 327724 309130 327776 309136
rect 327632 305652 327684 305658
rect 327632 305594 327684 305600
rect 327540 304292 327592 304298
rect 327540 304234 327592 304240
rect 327736 240961 327764 309130
rect 327828 307834 327856 317562
rect 327908 316328 327960 316334
rect 327908 316270 327960 316276
rect 327920 316062 327948 316270
rect 327908 316056 327960 316062
rect 327908 315998 327960 316004
rect 327816 307828 327868 307834
rect 327816 307770 327868 307776
rect 327828 306374 327856 307770
rect 327828 306346 327948 306374
rect 327722 240952 327778 240961
rect 327722 240887 327778 240896
rect 327920 240825 327948 306346
rect 328012 247625 328040 320062
rect 328196 311894 328224 320622
rect 328460 319660 328512 319666
rect 328460 319602 328512 319608
rect 328104 311866 328224 311894
rect 327998 247616 328054 247625
rect 327998 247551 328054 247560
rect 327906 240816 327962 240825
rect 327906 240751 327962 240760
rect 327446 234152 327502 234161
rect 327446 234087 327502 234096
rect 327722 234152 327778 234161
rect 327722 234087 327778 234096
rect 327172 216572 327224 216578
rect 327172 216514 327224 216520
rect 327092 16546 327672 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 327644 3482 327672 16546
rect 327736 3602 327764 234087
rect 328104 215218 328132 311866
rect 328366 231840 328422 231849
rect 328366 231775 328422 231784
rect 328380 231169 328408 231775
rect 328366 231160 328422 231169
rect 328366 231095 328422 231104
rect 328368 216572 328420 216578
rect 328368 216514 328420 216520
rect 328380 215966 328408 216514
rect 328368 215960 328420 215966
rect 328368 215902 328420 215908
rect 328092 215212 328144 215218
rect 328092 215154 328144 215160
rect 328368 215212 328420 215218
rect 328368 215154 328420 215160
rect 328380 214742 328408 215154
rect 328368 214736 328420 214742
rect 328368 214678 328420 214684
rect 328472 205630 328500 319602
rect 328564 212498 328592 320719
rect 328642 319968 328698 319977
rect 328642 319903 328698 319912
rect 328656 226953 328684 319903
rect 328736 317348 328788 317354
rect 328736 317290 328788 317296
rect 328748 231849 328776 317290
rect 328828 317008 328880 317014
rect 328828 316950 328880 316956
rect 328734 231840 328790 231849
rect 328734 231775 328790 231784
rect 328748 231441 328776 231775
rect 328840 231742 328868 316950
rect 328920 314424 328972 314430
rect 328920 314366 328972 314372
rect 328828 231736 328880 231742
rect 328932 231713 328960 314366
rect 329024 291854 329052 369378
rect 329116 325650 329144 370330
rect 331862 370288 331918 370297
rect 331862 370223 331918 370232
rect 329196 370116 329248 370122
rect 329196 370058 329248 370064
rect 329208 353258 329236 370058
rect 330484 369980 330536 369986
rect 330484 369922 330536 369928
rect 329196 353252 329248 353258
rect 329196 353194 329248 353200
rect 329104 325644 329156 325650
rect 329104 325586 329156 325592
rect 330206 320512 330262 320521
rect 330206 320447 330262 320456
rect 330024 318844 330076 318850
rect 330024 318786 330076 318792
rect 329840 318776 329892 318782
rect 329840 318718 329892 318724
rect 329104 318572 329156 318578
rect 329104 318514 329156 318520
rect 329116 300898 329144 318514
rect 329194 318064 329250 318073
rect 329194 317999 329250 318008
rect 329104 300892 329156 300898
rect 329104 300834 329156 300840
rect 329012 291848 329064 291854
rect 329012 291790 329064 291796
rect 329116 240786 329144 300834
rect 329208 294642 329236 317999
rect 329656 302932 329708 302938
rect 329656 302874 329708 302880
rect 329668 300150 329696 302874
rect 329656 300144 329708 300150
rect 329656 300086 329708 300092
rect 329196 294636 329248 294642
rect 329196 294578 329248 294584
rect 329104 240780 329156 240786
rect 329104 240722 329156 240728
rect 329286 231840 329342 231849
rect 329286 231775 329342 231784
rect 329196 231736 329248 231742
rect 328828 231678 328880 231684
rect 328918 231704 328974 231713
rect 329196 231678 329248 231684
rect 328918 231639 328974 231648
rect 328734 231432 328790 231441
rect 328734 231367 328790 231376
rect 328932 229094 328960 231639
rect 328932 229066 329144 229094
rect 328642 226944 328698 226953
rect 328642 226879 328698 226888
rect 328552 212492 328604 212498
rect 328552 212434 328604 212440
rect 328460 205624 328512 205630
rect 328460 205566 328512 205572
rect 329116 3602 329144 229066
rect 329208 4078 329236 231678
rect 329196 4072 329248 4078
rect 329196 4014 329248 4020
rect 327724 3596 327776 3602
rect 327724 3538 327776 3544
rect 329104 3596 329156 3602
rect 329104 3538 329156 3544
rect 324964 3392 325016 3398
rect 324964 3334 325016 3340
rect 325620 480 325648 3470
rect 327644 3454 328040 3482
rect 329300 3466 329328 231775
rect 329852 222086 329880 318718
rect 329932 316940 329984 316946
rect 329932 316882 329984 316888
rect 329944 227662 329972 316882
rect 330036 232665 330064 318786
rect 330116 318708 330168 318714
rect 330116 318650 330168 318656
rect 330128 234297 330156 318650
rect 330220 237318 330248 320447
rect 330392 318912 330444 318918
rect 330392 318854 330444 318860
rect 330300 314084 330352 314090
rect 330300 314026 330352 314032
rect 330312 238754 330340 314026
rect 330404 240106 330432 318854
rect 330496 273222 330524 369922
rect 331404 320136 331456 320142
rect 331404 320078 331456 320084
rect 331220 319116 331272 319122
rect 331220 319058 331272 319064
rect 330576 318028 330628 318034
rect 330576 317970 330628 317976
rect 330588 297430 330616 317970
rect 330576 297424 330628 297430
rect 330576 297366 330628 297372
rect 330484 273216 330536 273222
rect 330484 273158 330536 273164
rect 330392 240100 330444 240106
rect 330392 240042 330444 240048
rect 331128 240100 331180 240106
rect 331128 240042 331180 240048
rect 331140 238950 331168 240042
rect 331128 238944 331180 238950
rect 331128 238886 331180 238892
rect 330312 238726 330524 238754
rect 330208 237312 330260 237318
rect 330208 237254 330260 237260
rect 330220 236774 330248 237254
rect 330208 236768 330260 236774
rect 330208 236710 330260 236716
rect 330496 234433 330524 238726
rect 331140 236910 331168 238886
rect 331128 236904 331180 236910
rect 331128 236846 331180 236852
rect 330482 234424 330538 234433
rect 330482 234359 330538 234368
rect 330114 234288 330170 234297
rect 330114 234223 330170 234232
rect 330022 232656 330078 232665
rect 330022 232591 330078 232600
rect 329932 227656 329984 227662
rect 329932 227598 329984 227604
rect 329944 226370 329972 227598
rect 329932 226364 329984 226370
rect 329932 226306 329984 226312
rect 329840 222080 329892 222086
rect 329840 222022 329892 222028
rect 330300 222080 330352 222086
rect 330300 222022 330352 222028
rect 330312 221474 330340 222022
rect 330300 221468 330352 221474
rect 330300 221410 330352 221416
rect 329748 212492 329800 212498
rect 329748 212434 329800 212440
rect 329760 211818 329788 212434
rect 329748 211812 329800 211818
rect 329748 211754 329800 211760
rect 329748 205624 329800 205630
rect 329748 205566 329800 205572
rect 329760 205018 329788 205566
rect 329748 205012 329800 205018
rect 329748 204954 329800 204960
rect 329838 186960 329894 186969
rect 329838 186895 329894 186904
rect 329852 16574 329880 186895
rect 329852 16546 330432 16574
rect 326804 3392 326856 3398
rect 326804 3334 326856 3340
rect 326816 480 326844 3334
rect 328012 480 328040 3454
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 329288 3460 329340 3466
rect 329288 3402 329340 3408
rect 329208 480 329236 3402
rect 330404 480 330432 16546
rect 330496 3670 330524 234359
rect 330576 226364 330628 226370
rect 330576 226306 330628 226312
rect 330588 4146 330616 226306
rect 331232 223514 331260 319058
rect 331312 315444 331364 315450
rect 331312 315386 331364 315392
rect 331324 227594 331352 315386
rect 331416 234025 331444 320078
rect 331494 319424 331550 319433
rect 331494 319359 331550 319368
rect 331508 235890 331536 319359
rect 331588 319252 331640 319258
rect 331588 319194 331640 319200
rect 331600 240174 331628 319194
rect 331678 318200 331734 318209
rect 331678 318135 331734 318144
rect 331692 291922 331720 318135
rect 331680 291916 331732 291922
rect 331680 291858 331732 291864
rect 331588 240168 331640 240174
rect 331588 240110 331640 240116
rect 331496 235884 331548 235890
rect 331496 235826 331548 235832
rect 331508 235278 331536 235826
rect 331600 235346 331628 240110
rect 331588 235340 331640 235346
rect 331588 235282 331640 235288
rect 331496 235272 331548 235278
rect 331496 235214 331548 235220
rect 331496 234660 331548 234666
rect 331496 234602 331548 234608
rect 331402 234016 331458 234025
rect 331402 233951 331458 233960
rect 331508 231577 331536 234602
rect 331494 231568 331550 231577
rect 331494 231503 331550 231512
rect 331312 227588 331364 227594
rect 331312 227530 331364 227536
rect 331324 226370 331352 227530
rect 331312 226364 331364 226370
rect 331312 226306 331364 226312
rect 331220 223508 331272 223514
rect 331220 223450 331272 223456
rect 331876 73166 331904 370223
rect 334622 369880 334678 369889
rect 334622 369815 334678 369824
rect 332782 321056 332838 321065
rect 332782 320991 332838 321000
rect 331956 318980 332008 318986
rect 331956 318922 332008 318928
rect 331968 234666 331996 318922
rect 332690 318880 332746 318889
rect 332690 318815 332746 318824
rect 332046 317520 332102 317529
rect 332046 317455 332102 317464
rect 332060 298790 332088 317455
rect 332048 298784 332100 298790
rect 332048 298726 332100 298732
rect 332600 236700 332652 236706
rect 332600 236642 332652 236648
rect 331956 234660 332008 234666
rect 331956 234602 332008 234608
rect 331956 226364 332008 226370
rect 331956 226306 332008 226312
rect 331864 73160 331916 73166
rect 331864 73102 331916 73108
rect 330576 4140 330628 4146
rect 330576 4082 330628 4088
rect 331968 4078 331996 226306
rect 332048 223508 332100 223514
rect 332048 223450 332100 223456
rect 331956 4072 332008 4078
rect 331956 4014 332008 4020
rect 331588 4004 331640 4010
rect 331588 3946 331640 3952
rect 330484 3664 330536 3670
rect 330484 3606 330536 3612
rect 331600 480 331628 3946
rect 332060 3398 332088 223450
rect 332612 16574 332640 236642
rect 332704 219434 332732 318815
rect 332796 226114 332824 320991
rect 334438 320648 334494 320657
rect 334438 320583 334494 320592
rect 334346 320240 334402 320249
rect 334346 320175 334402 320184
rect 332968 320068 333020 320074
rect 332968 320010 333020 320016
rect 332876 319184 332928 319190
rect 332876 319126 332928 319132
rect 332888 226386 332916 319126
rect 332980 238882 333008 320010
rect 333060 320000 333112 320006
rect 333060 319942 333112 319948
rect 332968 238876 333020 238882
rect 332968 238818 333020 238824
rect 332980 236842 333008 238818
rect 332968 236836 333020 236842
rect 332968 236778 333020 236784
rect 333072 231169 333100 319942
rect 334254 319288 334310 319297
rect 334254 319223 334310 319232
rect 334162 319016 334218 319025
rect 334162 318951 334218 318960
rect 334072 317076 334124 317082
rect 334072 317018 334124 317024
rect 333980 237380 334032 237386
rect 333980 237322 334032 237328
rect 333992 236706 334020 237322
rect 333980 236700 334032 236706
rect 333980 236642 334032 236648
rect 333058 231160 333114 231169
rect 333058 231095 333114 231104
rect 333980 229152 334032 229158
rect 333980 229094 334032 229100
rect 332888 226358 333100 226386
rect 332796 226086 332916 226114
rect 332784 224936 332836 224942
rect 332784 224878 332836 224884
rect 332796 224330 332824 224878
rect 332888 224874 332916 226086
rect 333072 224942 333100 226358
rect 333060 224936 333112 224942
rect 333060 224878 333112 224884
rect 332876 224868 332928 224874
rect 332876 224810 332928 224816
rect 332784 224324 332836 224330
rect 332784 224266 332836 224272
rect 332888 224262 332916 224810
rect 332876 224256 332928 224262
rect 332876 224198 332928 224204
rect 332692 219428 332744 219434
rect 332692 219370 332744 219376
rect 332704 218754 332732 219370
rect 332692 218748 332744 218754
rect 332692 218690 332744 218696
rect 333992 16574 334020 229094
rect 334084 215286 334112 317018
rect 334176 229094 334204 318951
rect 334268 230353 334296 319223
rect 334360 232393 334388 320175
rect 334452 237386 334480 320583
rect 334532 318640 334584 318646
rect 334532 318582 334584 318588
rect 334440 237380 334492 237386
rect 334440 237322 334492 237328
rect 334346 232384 334402 232393
rect 334346 232319 334402 232328
rect 334254 230344 334310 230353
rect 334254 230279 334310 230288
rect 334176 229066 334296 229094
rect 334164 227724 334216 227730
rect 334164 227666 334216 227672
rect 334176 227118 334204 227666
rect 334164 227112 334216 227118
rect 334164 227054 334216 227060
rect 334268 223378 334296 229066
rect 334544 227730 334572 318582
rect 334532 227724 334584 227730
rect 334532 227666 334584 227672
rect 334256 223372 334308 223378
rect 334256 223314 334308 223320
rect 334072 215280 334124 215286
rect 334072 215222 334124 215228
rect 334084 214674 334112 215222
rect 334072 214668 334124 214674
rect 334072 214610 334124 214616
rect 334636 153202 334664 369815
rect 335358 321600 335414 321609
rect 335358 321535 335414 321544
rect 334714 318472 334770 318481
rect 334714 318407 334770 318416
rect 334728 293282 334756 318407
rect 334716 293276 334768 293282
rect 334716 293218 334768 293224
rect 334806 230344 334862 230353
rect 334806 230279 334862 230288
rect 334820 229809 334848 230279
rect 334806 229800 334862 229809
rect 334806 229735 334862 229744
rect 334808 223372 334860 223378
rect 334808 223314 334860 223320
rect 334820 222902 334848 223314
rect 334808 222896 334860 222902
rect 334808 222838 334860 222844
rect 335372 204270 335400 321535
rect 335450 321192 335506 321201
rect 335450 321127 335506 321136
rect 335464 225593 335492 321127
rect 335820 320272 335872 320278
rect 335820 320214 335872 320220
rect 335634 319152 335690 319161
rect 335634 319087 335690 319096
rect 335544 318368 335596 318374
rect 335544 318310 335596 318316
rect 335556 226234 335584 318310
rect 335648 228993 335676 319087
rect 335728 318504 335780 318510
rect 335728 318446 335780 318452
rect 335634 228984 335690 228993
rect 335634 228919 335690 228928
rect 335740 228313 335768 318446
rect 335832 231810 335860 320214
rect 335912 320204 335964 320210
rect 335912 320146 335964 320152
rect 335924 234569 335952 320146
rect 336016 319462 336044 371486
rect 345664 369912 345716 369918
rect 345664 369854 345716 369860
rect 338580 320612 338632 320618
rect 338580 320554 338632 320560
rect 336740 320476 336792 320482
rect 336740 320418 336792 320424
rect 336004 319456 336056 319462
rect 336004 319398 336056 319404
rect 336004 315376 336056 315382
rect 336004 315318 336056 315324
rect 336016 237454 336044 315318
rect 336004 237448 336056 237454
rect 336004 237390 336056 237396
rect 335910 234560 335966 234569
rect 335910 234495 335966 234504
rect 335820 231804 335872 231810
rect 335820 231746 335872 231752
rect 335726 228304 335782 228313
rect 335726 228239 335782 228248
rect 335544 226228 335596 226234
rect 335544 226170 335596 226176
rect 335450 225584 335506 225593
rect 335450 225519 335506 225528
rect 335360 204264 335412 204270
rect 335360 204206 335412 204212
rect 334624 153196 334676 153202
rect 334624 153138 334676 153144
rect 332612 16546 332732 16574
rect 333992 16546 334664 16574
rect 332048 3392 332100 3398
rect 332048 3334 332100 3340
rect 332704 480 332732 16546
rect 333886 6080 333942 6089
rect 333886 6015 333942 6024
rect 333900 480 333928 6015
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336016 4078 336044 237390
rect 336646 234560 336702 234569
rect 336646 234495 336702 234504
rect 336660 233889 336688 234495
rect 336646 233880 336702 233889
rect 336646 233815 336702 233824
rect 336648 231804 336700 231810
rect 336648 231746 336700 231752
rect 336660 231198 336688 231746
rect 336648 231192 336700 231198
rect 336648 231134 336700 231140
rect 336096 226228 336148 226234
rect 336096 226170 336148 226176
rect 336108 6526 336136 226170
rect 336752 211138 336780 320418
rect 338304 320408 338356 320414
rect 338304 320350 338356 320356
rect 336832 320340 336884 320346
rect 336832 320282 336884 320288
rect 336844 220794 336872 320282
rect 338212 319796 338264 319802
rect 338212 319738 338264 319744
rect 337016 319388 337068 319394
rect 337016 319330 337068 319336
rect 336924 316872 336976 316878
rect 336924 316814 336976 316820
rect 336936 229945 336964 316814
rect 337028 235958 337056 319330
rect 337016 235952 337068 235958
rect 337016 235894 337068 235900
rect 338028 235952 338080 235958
rect 338028 235894 338080 235900
rect 338040 235414 338068 235894
rect 338028 235408 338080 235414
rect 338028 235350 338080 235356
rect 336922 229936 336978 229945
rect 336922 229871 336978 229880
rect 338120 225004 338172 225010
rect 338120 224946 338172 224952
rect 336832 220788 336884 220794
rect 336832 220730 336884 220736
rect 338028 220788 338080 220794
rect 338028 220730 338080 220736
rect 338040 220250 338068 220730
rect 338028 220244 338080 220250
rect 338028 220186 338080 220192
rect 336740 211132 336792 211138
rect 336740 211074 336792 211080
rect 338028 211132 338080 211138
rect 338028 211074 338080 211080
rect 338040 210526 338068 211074
rect 338028 210520 338080 210526
rect 338028 210462 338080 210468
rect 336648 204264 336700 204270
rect 336648 204206 336700 204212
rect 336660 203590 336688 204206
rect 336648 203584 336700 203590
rect 336648 203526 336700 203532
rect 336738 197976 336794 197985
rect 336738 197911 336794 197920
rect 336752 16574 336780 197911
rect 338132 16574 338160 224946
rect 338224 216646 338252 319738
rect 338316 218006 338344 320350
rect 338394 320104 338450 320113
rect 338394 320039 338450 320048
rect 338304 218000 338356 218006
rect 338304 217942 338356 217948
rect 338316 217394 338344 217942
rect 338408 217938 338436 320039
rect 338488 319320 338540 319326
rect 338488 319262 338540 319268
rect 338500 222154 338528 319262
rect 338592 229022 338620 320554
rect 338670 320376 338726 320385
rect 338670 320311 338726 320320
rect 338580 229016 338632 229022
rect 338580 228958 338632 228964
rect 338488 222148 338540 222154
rect 338488 222090 338540 222096
rect 338684 220658 338712 320311
rect 340880 319728 340932 319734
rect 340880 319670 340932 319676
rect 339408 222148 339460 222154
rect 339408 222090 339460 222096
rect 339420 221610 339448 222090
rect 339408 221604 339460 221610
rect 339408 221546 339460 221552
rect 340892 220726 340920 319670
rect 340972 318232 341024 318238
rect 340972 318174 341024 318180
rect 340984 223582 341012 318174
rect 342260 312792 342312 312798
rect 342260 312734 342312 312740
rect 342272 228206 342300 312734
rect 345676 233238 345704 369854
rect 349252 318164 349304 318170
rect 349252 318106 349304 318112
rect 349160 259480 349212 259486
rect 349160 259422 349212 259428
rect 346400 245812 346452 245818
rect 346400 245754 346452 245760
rect 345664 233232 345716 233238
rect 345664 233174 345716 233180
rect 345020 229016 345072 229022
rect 345020 228958 345072 228964
rect 342260 228200 342312 228206
rect 342260 228142 342312 228148
rect 342272 227798 342300 228142
rect 342260 227792 342312 227798
rect 342260 227734 342312 227740
rect 342904 227792 342956 227798
rect 342904 227734 342956 227740
rect 340972 223576 341024 223582
rect 340972 223518 341024 223524
rect 341524 223576 341576 223582
rect 341524 223518 341576 223524
rect 340880 220720 340932 220726
rect 340880 220662 340932 220668
rect 338672 220652 338724 220658
rect 338672 220594 338724 220600
rect 339408 220652 339460 220658
rect 339408 220594 339460 220600
rect 339420 220114 339448 220594
rect 340892 220522 340920 220662
rect 340880 220516 340932 220522
rect 340880 220458 340932 220464
rect 339408 220108 339460 220114
rect 339408 220050 339460 220056
rect 338396 217932 338448 217938
rect 338396 217874 338448 217880
rect 338304 217388 338356 217394
rect 338304 217330 338356 217336
rect 338408 217326 338436 217874
rect 338396 217320 338448 217326
rect 338396 217262 338448 217268
rect 338212 216640 338264 216646
rect 338212 216582 338264 216588
rect 339408 216640 339460 216646
rect 339408 216582 339460 216588
rect 339420 216102 339448 216582
rect 339408 216096 339460 216102
rect 339408 216038 339460 216044
rect 341536 207670 341564 223518
rect 341616 220516 341668 220522
rect 341616 220458 341668 220464
rect 341628 209166 341656 220458
rect 341616 209160 341668 209166
rect 341616 209102 341668 209108
rect 341524 207664 341576 207670
rect 341524 207606 341576 207612
rect 340972 196648 341024 196654
rect 340972 196590 341024 196596
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 336096 6520 336148 6526
rect 336096 6462 336148 6468
rect 336280 4140 336332 4146
rect 336280 4082 336332 4088
rect 335912 4072 335964 4078
rect 335912 4014 335964 4020
rect 336004 4072 336056 4078
rect 336004 4014 336056 4020
rect 335924 3330 335952 4014
rect 335912 3324 335964 3330
rect 335912 3266 335964 3272
rect 336292 480 336320 4082
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339868 4004 339920 4010
rect 339868 3946 339920 3952
rect 339880 480 339908 3946
rect 340984 480 341012 196590
rect 342916 4078 342944 227734
rect 345032 16574 345060 228958
rect 346412 16574 346440 245754
rect 347778 167648 347834 167657
rect 347778 167583 347834 167592
rect 347792 16574 347820 167583
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 344560 7608 344612 7614
rect 344560 7550 344612 7556
rect 342904 4072 342956 4078
rect 342904 4014 342956 4020
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 343364 3324 343416 3330
rect 343364 3266 343416 3272
rect 343376 480 343404 3266
rect 344572 480 344600 7550
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3398 349200 259422
rect 349264 226302 349292 318106
rect 354680 318096 354732 318102
rect 354680 318038 354732 318044
rect 354692 236745 354720 318038
rect 358082 314936 358138 314945
rect 358082 314871 358138 314880
rect 354678 236736 354734 236745
rect 354678 236671 354734 236680
rect 355322 236736 355378 236745
rect 355322 236671 355378 236680
rect 351184 231192 351236 231198
rect 351184 231134 351236 231140
rect 349252 226296 349304 226302
rect 349252 226238 349304 226244
rect 349264 225010 349292 226238
rect 349252 225004 349304 225010
rect 349252 224946 349304 224952
rect 349804 225004 349856 225010
rect 349804 224946 349856 224952
rect 349252 216096 349304 216102
rect 349252 216038 349304 216044
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 349264 480 349292 216038
rect 349816 4826 349844 224946
rect 350538 178664 350594 178673
rect 350538 178599 350594 178608
rect 350552 6914 350580 178599
rect 351196 16574 351224 231134
rect 353944 220244 353996 220250
rect 353944 220186 353996 220192
rect 351196 16546 351316 16574
rect 350552 6886 351224 6914
rect 349804 4820 349856 4826
rect 349804 4762 349856 4768
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 6886
rect 351288 3058 351316 16546
rect 353956 4146 353984 220186
rect 354678 202192 354734 202201
rect 354678 202127 354734 202136
rect 354692 16574 354720 202127
rect 354692 16546 355272 16574
rect 353944 4140 353996 4146
rect 353944 4082 353996 4088
rect 354036 4072 354088 4078
rect 354036 4014 354088 4020
rect 351276 3052 351328 3058
rect 351276 2994 351328 3000
rect 352840 3052 352892 3058
rect 352840 2994 352892 3000
rect 352852 480 352880 2994
rect 354048 480 354076 4014
rect 355244 480 355272 16546
rect 355336 7614 355364 236671
rect 356060 232552 356112 232558
rect 356060 232494 356112 232500
rect 356072 16574 356100 232494
rect 357532 195288 357584 195294
rect 357532 195230 357584 195236
rect 356072 16546 356376 16574
rect 355324 7608 355376 7614
rect 355324 7550 355376 7556
rect 356348 480 356376 16546
rect 357440 4004 357492 4010
rect 357440 3946 357492 3952
rect 357452 1986 357480 3946
rect 357544 3398 357572 195230
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 358096 2922 358124 314871
rect 363616 259418 363644 372098
rect 577504 372088 577556 372094
rect 577504 372030 577556 372036
rect 475382 317520 475438 317529
rect 475382 317455 475438 317464
rect 364340 316804 364392 316810
rect 364340 316746 364392 316752
rect 363604 259412 363656 259418
rect 363604 259354 363656 259360
rect 358820 224392 358872 224398
rect 358820 224334 358872 224340
rect 358832 16574 358860 224334
rect 362960 221604 363012 221610
rect 362960 221546 363012 221552
rect 361580 164892 361632 164898
rect 361580 164834 361632 164840
rect 361592 16574 361620 164834
rect 362972 16574 363000 221546
rect 364352 16574 364380 316746
rect 400864 316736 400916 316742
rect 400864 316678 400916 316684
rect 367100 315308 367152 315314
rect 367100 315250 367152 315256
rect 365810 138680 365866 138689
rect 365810 138615 365866 138624
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 364352 16546 364656 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358084 2916 358136 2922
rect 358084 2858 358136 2864
rect 357452 1958 357572 1986
rect 357544 480 357572 1958
rect 358740 480 358768 3334
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 2916 361172 2922
rect 361120 2858 361172 2864
rect 361132 480 361160 2858
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364628 480 364656 16546
rect 365824 480 365852 138615
rect 367112 16574 367140 315250
rect 373998 314800 374054 314809
rect 373998 314735 374054 314744
rect 396080 314764 396132 314770
rect 371240 244384 371292 244390
rect 371240 244326 371292 244332
rect 369860 235408 369912 235414
rect 369860 235350 369912 235356
rect 369872 16574 369900 235350
rect 367112 16546 367784 16574
rect 369872 16546 370176 16574
rect 367008 4072 367060 4078
rect 367008 4014 367060 4020
rect 367020 480 367048 4014
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369400 8968 369452 8974
rect 369400 8910 369452 8916
rect 369412 480 369440 8910
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 244326
rect 372896 3936 372948 3942
rect 372896 3878 372948 3884
rect 372908 480 372936 3878
rect 374012 3398 374040 314735
rect 396080 314706 396132 314712
rect 378138 312080 378194 312089
rect 378138 312015 378194 312024
rect 374092 229764 374144 229770
rect 374092 229706 374144 229712
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 229706
rect 376024 227112 376076 227118
rect 376024 227054 376076 227060
rect 376036 3398 376064 227054
rect 378152 16574 378180 312015
rect 391940 310616 391992 310622
rect 391940 310558 391992 310564
rect 382280 294024 382332 294030
rect 382280 293966 382332 293972
rect 380900 223032 380952 223038
rect 380900 222974 380952 222980
rect 378784 214736 378836 214742
rect 378784 214678 378836 214684
rect 378152 16546 378456 16574
rect 376484 3868 376536 3874
rect 376484 3810 376536 3816
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 376024 3392 376076 3398
rect 376024 3334 376076 3340
rect 375300 480 375328 3334
rect 376496 480 376524 3810
rect 377680 3392 377732 3398
rect 377680 3334 377732 3340
rect 377692 480 377720 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378796 4146 378824 214678
rect 380912 16574 380940 222974
rect 382292 16574 382320 293966
rect 386420 263628 386472 263634
rect 386420 263570 386472 263576
rect 385040 250504 385092 250510
rect 385040 250446 385092 250452
rect 385052 16574 385080 250446
rect 385684 225684 385736 225690
rect 385684 225626 385736 225632
rect 380912 16546 381216 16574
rect 382292 16546 382412 16574
rect 385052 16546 385632 16574
rect 378784 4140 378836 4146
rect 378784 4082 378836 4088
rect 379978 3632 380034 3641
rect 379978 3567 380034 3576
rect 379992 480 380020 3567
rect 381188 480 381216 16546
rect 382384 480 382412 16546
rect 384764 4140 384816 4146
rect 384764 4082 384816 4088
rect 383566 3496 383622 3505
rect 383566 3431 383622 3440
rect 383580 480 383608 3431
rect 384776 480 384804 4082
rect 385604 3482 385632 16546
rect 385696 3738 385724 225626
rect 386432 16574 386460 263570
rect 389180 248464 389232 248470
rect 389180 248406 389232 248412
rect 389192 16574 389220 248406
rect 390652 228404 390704 228410
rect 390652 228346 390704 228352
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 385684 3732 385736 3738
rect 385684 3674 385736 3680
rect 385604 3454 386000 3482
rect 385972 480 386000 3454
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 388260 3732 388312 3738
rect 388260 3674 388312 3680
rect 388272 480 388300 3674
rect 389468 480 389496 16546
rect 390560 3868 390612 3874
rect 390560 3810 390612 3816
rect 390572 1850 390600 3810
rect 390664 3398 390692 228346
rect 391952 16574 391980 310558
rect 394700 218068 394752 218074
rect 394700 218010 394752 218016
rect 394712 16574 394740 218010
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 1822 390692 1850
rect 390664 480 390692 1822
rect 391860 480 391888 3334
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394240 6452 394292 6458
rect 394240 6394 394292 6400
rect 394252 480 394280 6394
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 314706
rect 398840 249076 398892 249082
rect 398840 249018 398892 249024
rect 397736 6384 397788 6390
rect 397736 6326 397788 6332
rect 397748 480 397776 6326
rect 398852 2650 398880 249018
rect 398932 213308 398984 213314
rect 398932 213250 398984 213256
rect 398840 2644 398892 2650
rect 398840 2586 398892 2592
rect 398944 480 398972 213250
rect 400876 3738 400904 316678
rect 407120 314696 407172 314702
rect 407120 314638 407172 314644
rect 402980 258188 403032 258194
rect 402980 258130 403032 258136
rect 402992 16574 403020 258130
rect 405740 233912 405792 233918
rect 405740 233854 405792 233860
rect 405752 16574 405780 233854
rect 406384 224324 406436 224330
rect 406384 224266 406436 224272
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 401322 6896 401378 6905
rect 401322 6831 401378 6840
rect 400864 3732 400916 3738
rect 400864 3674 400916 3680
rect 400128 2644 400180 2650
rect 400128 2586 400180 2592
rect 400140 480 400168 2586
rect 401336 480 401364 6831
rect 402520 3936 402572 3942
rect 402520 3878 402572 3884
rect 402532 480 402560 3878
rect 403636 480 403664 16546
rect 404818 6760 404874 6769
rect 404818 6695 404874 6704
rect 404832 480 404860 6695
rect 406028 480 406056 16546
rect 406396 3126 406424 224266
rect 407132 3210 407160 314638
rect 431960 314016 432012 314022
rect 431960 313958 432012 313964
rect 422944 313404 422996 313410
rect 422944 313346 422996 313352
rect 409880 311908 409932 311914
rect 409880 311850 409932 311856
rect 407212 267776 407264 267782
rect 407212 267718 407264 267724
rect 407224 3398 407252 267718
rect 409892 16574 409920 311850
rect 414020 311160 414072 311166
rect 414020 311102 414072 311108
rect 411904 221536 411956 221542
rect 411904 221478 411956 221484
rect 411260 171828 411312 171834
rect 411260 171770 411312 171776
rect 409892 16546 410840 16574
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 406384 3120 406436 3126
rect 406384 3062 406436 3068
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 409604 3120 409656 3126
rect 409604 3062 409656 3068
rect 409616 480 409644 3062
rect 410812 480 410840 16546
rect 411272 6914 411300 171770
rect 411916 16574 411944 221478
rect 414032 16574 414060 311102
rect 416780 308440 416832 308446
rect 416780 308382 416832 308388
rect 415400 217388 415452 217394
rect 415400 217330 415452 217336
rect 411916 16546 412036 16574
rect 414032 16546 414336 16574
rect 411272 6886 411944 6914
rect 411916 480 411944 6886
rect 412008 4146 412036 16546
rect 411996 4140 412048 4146
rect 411996 4082 412048 4088
rect 413100 4140 413152 4146
rect 413100 4082 413152 4088
rect 413112 480 413140 4082
rect 414308 480 414336 16546
rect 415412 3398 415440 217330
rect 415492 189780 415544 189786
rect 415492 189722 415544 189728
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 189722
rect 416792 6914 416820 308382
rect 418802 283520 418858 283529
rect 418802 283455 418858 283464
rect 417424 210520 417476 210526
rect 417424 210462 417476 210468
rect 417436 16574 417464 210462
rect 418158 156632 418214 156641
rect 418158 156567 418214 156576
rect 418172 16574 418200 156567
rect 418816 20670 418844 283455
rect 420920 253972 420972 253978
rect 420920 253914 420972 253920
rect 418804 20664 418856 20670
rect 418804 20606 418856 20612
rect 417436 16546 417556 16574
rect 418172 16546 418568 16574
rect 416792 6886 417464 6914
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 6886
rect 417528 3330 417556 16546
rect 417516 3324 417568 3330
rect 417516 3266 417568 3272
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420184 3324 420236 3330
rect 420184 3266 420236 3272
rect 420196 480 420224 3266
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 253914
rect 421564 231124 421616 231130
rect 421564 231066 421616 231072
rect 421576 3330 421604 231066
rect 422576 14476 422628 14482
rect 422576 14418 422628 14424
rect 421564 3324 421616 3330
rect 421564 3266 421616 3272
rect 422588 480 422616 14418
rect 422956 3398 422984 313346
rect 427820 313336 427872 313342
rect 427820 313278 427872 313284
rect 426440 220176 426492 220182
rect 426440 220118 426492 220124
rect 425704 209160 425756 209166
rect 425704 209102 425756 209108
rect 425716 4146 425744 209102
rect 426452 16574 426480 220118
rect 427832 16574 427860 313278
rect 430580 216028 430632 216034
rect 430580 215970 430632 215976
rect 430592 16574 430620 215970
rect 431972 16574 432000 313958
rect 441620 313948 441672 313954
rect 441620 313890 441672 313896
rect 438860 262268 438912 262274
rect 438860 262210 438912 262216
rect 434718 254008 434774 254017
rect 434718 253943 434774 253952
rect 434732 16574 434760 253943
rect 436744 207664 436796 207670
rect 436744 207606 436796 207612
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 431972 16546 432092 16574
rect 434732 16546 435128 16574
rect 426162 6624 426218 6633
rect 426162 6559 426218 6568
rect 425704 4140 425756 4146
rect 425704 4082 425756 4088
rect 422944 3392 422996 3398
rect 422944 3334 422996 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423772 3324 423824 3330
rect 423772 3266 423824 3272
rect 423784 480 423812 3266
rect 424980 480 425008 3334
rect 426176 480 426204 6559
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 6316 429712 6322
rect 429660 6258 429712 6264
rect 429672 480 429700 6258
rect 430868 480 430896 16546
rect 432064 480 432092 16546
rect 433248 6248 433300 6254
rect 433248 6190 433300 6196
rect 433260 480 433288 6190
rect 434444 4140 434496 4146
rect 434444 4082 434496 4088
rect 434456 480 434484 4082
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 436650 6488 436706 6497
rect 436650 6423 436706 6432
rect 436664 3210 436692 6423
rect 436756 3398 436784 207606
rect 438872 16574 438900 262210
rect 440238 229936 440294 229945
rect 440238 229871 440294 229880
rect 438872 16546 439176 16574
rect 436744 3392 436796 3398
rect 436744 3334 436796 3340
rect 437940 3392 437992 3398
rect 437940 3334 437992 3340
rect 436664 3182 436784 3210
rect 436756 480 436784 3182
rect 437952 480 437980 3334
rect 439148 480 439176 16546
rect 440252 3398 440280 229871
rect 441632 16574 441660 313890
rect 445760 300892 445812 300898
rect 445760 300834 445812 300840
rect 443000 247172 443052 247178
rect 443000 247114 443052 247120
rect 443012 16574 443040 247114
rect 443644 225616 443696 225622
rect 443644 225558 443696 225564
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 440330 6352 440386 6361
rect 440330 6287 440386 6296
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 6287
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 443656 3398 443684 225558
rect 443644 3392 443696 3398
rect 443644 3334 443696 3340
rect 445024 3392 445076 3398
rect 445024 3334 445076 3340
rect 445036 480 445064 3334
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 300834
rect 452660 300144 452712 300150
rect 452660 300086 452712 300092
rect 447784 222964 447836 222970
rect 447784 222906 447836 222912
rect 447138 169008 447194 169017
rect 447138 168943 447194 168952
rect 447152 16574 447180 168943
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 447796 3058 447824 222906
rect 451280 214668 451332 214674
rect 451280 214610 451332 214616
rect 449898 151056 449954 151065
rect 449898 150991 449954 151000
rect 449912 16574 449940 150991
rect 451292 16574 451320 214610
rect 452672 16574 452700 300086
rect 456800 297424 456852 297430
rect 456800 297366 456852 297372
rect 454684 213240 454736 213246
rect 454684 213182 454736 213188
rect 454040 149728 454092 149734
rect 454040 149670 454092 149676
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 449808 4820 449860 4826
rect 449808 4762 449860 4768
rect 447784 3052 447836 3058
rect 447784 2994 447836 3000
rect 448612 3052 448664 3058
rect 448612 2994 448664 3000
rect 448624 480 448652 2994
rect 449820 480 449848 4762
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 149670
rect 454696 3330 454724 213182
rect 454684 3324 454736 3330
rect 454684 3266 454736 3272
rect 455696 3324 455748 3330
rect 455696 3266 455748 3272
rect 455708 480 455736 3266
rect 456812 3210 456840 297366
rect 463700 294636 463752 294642
rect 463700 294578 463752 294584
rect 458180 227044 458232 227050
rect 458180 226986 458232 226992
rect 458192 16574 458220 226986
rect 462320 218816 462372 218822
rect 462320 218758 462372 218764
rect 461584 205012 461636 205018
rect 461584 204954 461636 204960
rect 461596 16574 461624 204954
rect 458192 16546 459232 16574
rect 461596 16546 461716 16574
rect 456890 15872 456946 15881
rect 456890 15807 456946 15816
rect 456904 3398 456932 15807
rect 456892 3392 456944 3398
rect 456892 3334 456944 3340
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 456812 3182 456932 3210
rect 456904 480 456932 3182
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 460388 6520 460440 6526
rect 460388 6462 460440 6468
rect 460400 480 460428 6462
rect 461584 6180 461636 6186
rect 461584 6122 461636 6128
rect 461596 480 461624 6122
rect 461688 3398 461716 16546
rect 461676 3392 461728 3398
rect 461676 3334 461728 3340
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 354 462360 218758
rect 463712 16574 463740 294578
rect 466460 293276 466512 293282
rect 466460 293218 466512 293224
rect 465080 211880 465132 211886
rect 465080 211822 465132 211828
rect 465092 16574 465120 211822
rect 466472 16574 466500 293218
rect 470600 291848 470652 291854
rect 470600 291790 470652 291796
rect 467840 264988 467892 264994
rect 467840 264930 467892 264936
rect 467852 16574 467880 264930
rect 463712 16546 464016 16574
rect 465092 16546 465856 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 463988 480 464016 16546
rect 465170 6216 465226 6225
rect 465170 6151 465226 6160
rect 465184 480 465212 6151
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469864 3392 469916 3398
rect 469864 3334 469916 3340
rect 469876 480 469904 3334
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 291790
rect 472624 203584 472676 203590
rect 472624 203526 472676 203532
rect 471978 146976 472034 146985
rect 471978 146911 472034 146920
rect 471992 16574 472020 146911
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3058 472664 203526
rect 474738 25528 474794 25537
rect 474738 25463 474794 25472
rect 474752 16574 474780 25463
rect 474752 16546 475332 16574
rect 474556 7608 474608 7614
rect 474556 7550 474608 7556
rect 472624 3052 472676 3058
rect 472624 2994 472676 3000
rect 473452 3052 473504 3058
rect 473452 2994 473504 3000
rect 473464 480 473492 2994
rect 474568 480 474596 7550
rect 475304 3482 475332 16546
rect 475396 5574 475424 317455
rect 488538 316840 488594 316849
rect 488538 316775 488594 316784
rect 481640 292596 481692 292602
rect 481640 292538 481692 292544
rect 478144 221468 478196 221474
rect 478144 221410 478196 221416
rect 476120 210452 476172 210458
rect 476120 210394 476172 210400
rect 476132 16574 476160 210394
rect 476132 16546 476528 16574
rect 475384 5568 475436 5574
rect 475384 5510 475436 5516
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478052 5568 478104 5574
rect 478052 5510 478104 5516
rect 478064 3482 478092 5510
rect 478156 4146 478184 221410
rect 478880 145580 478932 145586
rect 478880 145522 478932 145528
rect 478144 4140 478196 4146
rect 478144 4082 478196 4088
rect 478064 3454 478184 3482
rect 478156 480 478184 3454
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 145522
rect 481652 6914 481680 292538
rect 481732 255332 481784 255338
rect 481732 255274 481784 255280
rect 481744 16574 481772 255274
rect 487160 236904 487212 236910
rect 487160 236846 487212 236852
rect 483018 234152 483074 234161
rect 483018 234087 483074 234096
rect 483032 16574 483060 234087
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 481652 6886 481772 6914
rect 480536 4140 480588 4146
rect 480536 4082 480588 4088
rect 480548 480 480576 4082
rect 481744 480 481772 6886
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 485228 3664 485280 3670
rect 485228 3606 485280 3612
rect 485240 480 485268 3606
rect 486422 3360 486478 3369
rect 486422 3295 486478 3304
rect 486436 480 486464 3295
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 236846
rect 488552 16574 488580 316775
rect 569958 316704 570014 316713
rect 569958 316639 570014 316648
rect 493324 316260 493376 316266
rect 493324 316202 493376 316208
rect 491300 245744 491352 245750
rect 491300 245686 491352 245692
rect 489920 238808 489972 238814
rect 489920 238750 489972 238756
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 480 489960 238750
rect 490010 231160 490066 231169
rect 490010 231095 490066 231104
rect 490024 16574 490052 231095
rect 491312 16574 491340 245686
rect 492680 242956 492732 242962
rect 492680 242898 492732 242904
rect 492692 16574 492720 242898
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 493336 3670 493364 316202
rect 534080 316192 534132 316198
rect 534080 316134 534132 316140
rect 538218 316160 538274 316169
rect 500224 312724 500276 312730
rect 500224 312666 500276 312672
rect 498200 270564 498252 270570
rect 498200 270506 498252 270512
rect 496820 258120 496872 258126
rect 496820 258062 496872 258068
rect 494060 236836 494112 236842
rect 494060 236778 494112 236784
rect 494072 16574 494100 236778
rect 496832 16574 496860 258062
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 493324 3664 493376 3670
rect 493324 3606 493376 3612
rect 494716 480 494744 16546
rect 495900 3596 495952 3602
rect 495900 3538 495952 3544
rect 495912 480 495940 3538
rect 497108 480 497136 16546
rect 498212 3602 498240 270506
rect 499580 245676 499632 245682
rect 499580 245618 499632 245624
rect 498292 235340 498344 235346
rect 498292 235282 498344 235288
rect 498200 3596 498252 3602
rect 498200 3538 498252 3544
rect 498304 3482 498332 235282
rect 499592 16574 499620 245618
rect 499592 16546 500172 16574
rect 499028 3596 499080 3602
rect 499028 3538 499080 3544
rect 498212 3454 498332 3482
rect 498212 480 498240 3454
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3538
rect 500144 3482 500172 16546
rect 500236 3602 500264 312666
rect 511264 312656 511316 312662
rect 511264 312598 511316 312604
rect 508502 311944 508558 311953
rect 508502 311879 508558 311888
rect 506480 251252 506532 251258
rect 506480 251194 506532 251200
rect 503720 244316 503772 244322
rect 503720 244258 503772 244264
rect 502982 234016 503038 234025
rect 502982 233951 503038 233960
rect 500960 218748 501012 218754
rect 500960 218690 501012 218696
rect 500972 16574 501000 218690
rect 500972 16546 501368 16574
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 500144 3454 500632 3482
rect 500604 480 500632 3454
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 3602 503024 233951
rect 502892 3596 502944 3602
rect 502892 3538 502944 3544
rect 502984 3596 503036 3602
rect 502984 3538 503036 3544
rect 502904 3482 502932 3538
rect 502904 3454 503024 3482
rect 502996 480 503024 3454
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 244258
rect 505376 3596 505428 3602
rect 505376 3538 505428 3544
rect 505388 480 505416 3538
rect 506492 480 506520 251194
rect 506572 247104 506624 247110
rect 506572 247046 506624 247052
rect 506584 16574 506612 247046
rect 507858 232656 507914 232665
rect 507858 232591 507914 232600
rect 507872 16574 507900 232591
rect 506584 16546 507256 16574
rect 507872 16546 508452 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508424 3482 508452 16546
rect 508516 4146 508544 311879
rect 510620 252612 510672 252618
rect 510620 252554 510672 252560
rect 510632 6914 510660 252554
rect 511276 16574 511304 312598
rect 526444 312588 526496 312594
rect 526444 312530 526496 312536
rect 523040 307828 523092 307834
rect 523040 307770 523092 307776
rect 512644 234660 512696 234666
rect 512644 234602 512696 234608
rect 512000 144220 512052 144226
rect 512000 144162 512052 144168
rect 511276 16546 511396 16574
rect 510632 6886 511304 6914
rect 508504 4140 508556 4146
rect 508504 4082 508556 4088
rect 510068 4140 510120 4146
rect 510068 4082 510120 4088
rect 508424 3454 508912 3482
rect 508884 480 508912 3454
rect 510080 480 510108 4082
rect 511276 480 511304 6886
rect 511368 2922 511396 16546
rect 511356 2916 511408 2922
rect 511356 2858 511408 2864
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 144162
rect 512656 3194 512684 234602
rect 518900 211812 518952 211818
rect 518900 211754 518952 211760
rect 514850 191040 514906 191049
rect 514850 190975 514906 190984
rect 514864 6914 514892 190975
rect 517518 189680 517574 189689
rect 517518 189615 517574 189624
rect 517532 16574 517560 189615
rect 517532 16546 517928 16574
rect 514772 6886 514892 6914
rect 512644 3188 512696 3194
rect 512644 3130 512696 3136
rect 513564 2916 513616 2922
rect 513564 2858 513616 2864
rect 513576 480 513604 2858
rect 514772 480 514800 6886
rect 517152 3528 517204 3534
rect 517152 3470 517204 3476
rect 515956 3188 516008 3194
rect 515956 3130 516008 3136
rect 515968 480 515996 3130
rect 517164 480 517192 3470
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 518912 6914 518940 211754
rect 521660 186992 521712 186998
rect 521660 186934 521712 186940
rect 519544 141432 519596 141438
rect 519544 141374 519596 141380
rect 519556 16574 519584 141374
rect 519556 16546 519676 16574
rect 518912 6886 519584 6914
rect 519556 480 519584 6886
rect 519648 3262 519676 16546
rect 520740 3460 520792 3466
rect 520740 3402 520792 3408
rect 519636 3256 519688 3262
rect 519636 3198 519688 3204
rect 520752 480 520780 3402
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521672 354 521700 186934
rect 523052 3534 523080 307770
rect 523130 228440 523186 228449
rect 523130 228375 523186 228384
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 228375
rect 525798 225584 525854 225593
rect 525798 225519 525854 225528
rect 525812 16574 525840 225519
rect 525812 16546 526208 16574
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525432 3256 525484 3262
rect 525432 3198 525484 3204
rect 525444 480 525472 3198
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 526456 3534 526484 312530
rect 529204 236768 529256 236774
rect 529204 236710 529256 236716
rect 527824 29640 527876 29646
rect 527824 29582 527876 29588
rect 527836 4146 527864 29582
rect 528558 10296 528614 10305
rect 528558 10231 528614 10240
rect 527824 4140 527876 4146
rect 527824 4082 527876 4088
rect 526444 3528 526496 3534
rect 526444 3470 526496 3476
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 527836 480 527864 3470
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 10231
rect 529216 3466 529244 236710
rect 532698 233880 532754 233889
rect 532698 233815 532754 233824
rect 530584 209092 530636 209098
rect 530584 209034 530636 209040
rect 530124 4140 530176 4146
rect 530124 4082 530176 4088
rect 529204 3460 529256 3466
rect 529204 3402 529256 3408
rect 530136 480 530164 4082
rect 530596 3058 530624 209034
rect 532712 16574 532740 233815
rect 534092 16574 534120 316134
rect 538218 316095 538274 316104
rect 547972 316124 548024 316130
rect 536102 229800 536158 229809
rect 536102 229735 536158 229744
rect 535460 185632 535512 185638
rect 535460 185574 535512 185580
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 531320 3732 531372 3738
rect 531320 3674 531372 3680
rect 530584 3052 530636 3058
rect 530584 2994 530636 3000
rect 531332 480 531360 3674
rect 532516 3052 532568 3058
rect 532516 2994 532568 3000
rect 532528 480 532556 2994
rect 533724 480 533752 16546
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 535472 6914 535500 185574
rect 536116 16574 536144 229735
rect 537484 224256 537536 224262
rect 537484 224198 537536 224204
rect 536116 16546 536236 16574
rect 535472 6886 536144 6914
rect 536116 480 536144 6886
rect 536208 3534 536236 16546
rect 537496 3942 537524 224198
rect 537484 3936 537536 3942
rect 537484 3878 537536 3884
rect 536196 3528 536248 3534
rect 536196 3470 536248 3476
rect 537208 3528 537260 3534
rect 537208 3470 537260 3476
rect 537220 480 537248 3470
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 316095
rect 547972 316066 548024 316072
rect 543004 310548 543056 310554
rect 543004 310490 543056 310496
rect 540980 305652 541032 305658
rect 540980 305594 541032 305600
rect 540244 236700 540296 236706
rect 540244 236642 540296 236648
rect 539692 184204 539744 184210
rect 539692 184146 539744 184152
rect 539704 6914 539732 184146
rect 539612 6886 539732 6914
rect 539612 480 539640 6886
rect 540256 3534 540284 236642
rect 540992 16574 541020 305594
rect 542360 181484 542412 181490
rect 542360 181426 542412 181432
rect 542372 16574 542400 181426
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 540796 3936 540848 3942
rect 540796 3878 540848 3884
rect 540244 3528 540296 3534
rect 540244 3470 540296 3476
rect 540808 480 540836 3878
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3126 543044 310490
rect 543740 222896 543792 222902
rect 543740 222838 543792 222844
rect 543752 16574 543780 222838
rect 547144 214600 547196 214606
rect 547144 214542 547196 214548
rect 546498 182880 546554 182889
rect 546498 182815 546554 182824
rect 543752 16546 544424 16574
rect 543004 3120 543056 3126
rect 543004 3062 543056 3068
rect 544396 480 544424 16546
rect 545488 3120 545540 3126
rect 545488 3062 545540 3068
rect 545500 480 545528 3062
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 182815
rect 547156 4010 547184 214542
rect 547984 16574 548012 316066
rect 554044 316056 554096 316062
rect 554044 315998 554096 316004
rect 550640 235272 550692 235278
rect 550640 235214 550692 235220
rect 550652 16574 550680 235214
rect 553400 204944 553452 204950
rect 553400 204886 553452 204892
rect 553412 16574 553440 204886
rect 547984 16546 548656 16574
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 547144 4004 547196 4010
rect 547144 3946 547196 3952
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547892 480 547920 3470
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550272 4004 550324 4010
rect 550272 3946 550324 3952
rect 550284 480 550312 3946
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 3664 552716 3670
rect 552664 3606 552716 3612
rect 552676 480 552704 3606
rect 553780 480 553808 16546
rect 554056 3602 554084 315998
rect 565820 309800 565872 309806
rect 565820 309742 565872 309748
rect 558920 309188 558972 309194
rect 558920 309130 558972 309136
rect 555422 232520 555478 232529
rect 555422 232455 555478 232464
rect 554044 3596 554096 3602
rect 554044 3538 554096 3544
rect 555436 3466 555464 232455
rect 557538 228304 557594 228313
rect 557538 228239 557594 228248
rect 555516 137284 555568 137290
rect 555516 137226 555568 137232
rect 555528 3534 555556 137226
rect 557552 16574 557580 228239
rect 558932 16574 558960 309130
rect 563060 304292 563112 304298
rect 563060 304234 563112 304240
rect 562322 226944 562378 226953
rect 562322 226879 562378 226888
rect 559564 180124 559616 180130
rect 559564 180066 559616 180072
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 556160 3596 556212 3602
rect 556160 3538 556212 3544
rect 555516 3528 555568 3534
rect 555516 3470 555568 3476
rect 554964 3460 555016 3466
rect 554964 3402 555016 3408
rect 555424 3460 555476 3466
rect 555424 3402 555476 3408
rect 554976 480 555004 3402
rect 556172 480 556200 3538
rect 557356 3528 557408 3534
rect 557356 3470 557408 3476
rect 557368 480 557396 3470
rect 558564 480 558592 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559576 3534 559604 180066
rect 559564 3528 559616 3534
rect 559564 3470 559616 3476
rect 560852 3528 560904 3534
rect 560852 3470 560904 3476
rect 560864 480 560892 3470
rect 562048 3460 562100 3466
rect 562048 3402 562100 3408
rect 562060 480 562088 3402
rect 562336 3330 562364 226879
rect 562324 3324 562376 3330
rect 562324 3266 562376 3272
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 304234
rect 565084 217320 565136 217326
rect 565084 217262 565136 217268
rect 564532 177336 564584 177342
rect 564532 177278 564584 177284
rect 563704 175976 563756 175982
rect 563704 175918 563756 175924
rect 563716 4010 563744 175918
rect 564544 6914 564572 177278
rect 564452 6886 564572 6914
rect 563704 4004 563756 4010
rect 563704 3946 563756 3952
rect 564452 480 564480 6886
rect 565096 3466 565124 217262
rect 565832 16574 565860 309742
rect 568580 220108 568632 220114
rect 568580 220050 568632 220056
rect 568592 16574 568620 220050
rect 569972 16574 570000 316639
rect 574742 302288 574798 302297
rect 574742 302223 574798 302232
rect 572812 298784 572864 298790
rect 572812 298726 572864 298732
rect 571340 174548 571392 174554
rect 571340 174490 571392 174496
rect 565832 16546 566872 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 565084 3460 565136 3466
rect 565084 3402 565136 3408
rect 565636 3324 565688 3330
rect 565636 3266 565688 3272
rect 565648 480 565676 3266
rect 566844 480 566872 16546
rect 568028 4004 568080 4010
rect 568028 3946 568080 3952
rect 568040 480 568068 3946
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 174490
rect 572824 16574 572852 298726
rect 574100 170400 574152 170406
rect 574100 170342 574152 170348
rect 574112 16574 574140 170342
rect 572824 16546 573496 16574
rect 574112 16546 574692 16574
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 572732 480 572760 3402
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 574664 3482 574692 16546
rect 574756 3874 574784 302223
rect 575480 215960 575532 215966
rect 575480 215902 575532 215908
rect 575492 16574 575520 215902
rect 577516 179382 577544 372030
rect 577608 193186 577636 372982
rect 580262 371784 580318 371793
rect 580262 371719 580318 371728
rect 580172 370524 580224 370530
rect 580172 370466 580224 370472
rect 580184 365129 580212 370466
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 579620 353252 579672 353258
rect 579620 353194 579672 353200
rect 579632 351937 579660 353194
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 577596 193180 577648 193186
rect 577596 193122 577648 193128
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 577504 179376 577556 179382
rect 577504 179318 577556 179324
rect 579712 179376 579764 179382
rect 579712 179318 579764 179324
rect 579724 179217 579752 179318
rect 579710 179208 579766 179217
rect 579710 179143 579766 179152
rect 578240 173188 578292 173194
rect 578240 173130 578292 173136
rect 578252 16574 578280 173130
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580276 112849 580304 371719
rect 580356 370660 580408 370666
rect 580356 370602 580408 370608
rect 580368 139369 580396 370602
rect 580540 370592 580592 370598
rect 580540 370534 580592 370540
rect 580448 319456 580500 319462
rect 580448 319398 580500 319404
rect 580460 312089 580488 319398
rect 580446 312080 580502 312089
rect 580446 312015 580502 312024
rect 580448 306400 580500 306406
rect 580448 306342 580500 306348
rect 580460 298761 580488 306342
rect 580446 298752 580502 298761
rect 580446 298687 580502 298696
rect 580446 289096 580502 289105
rect 580446 289031 580502 289040
rect 580354 139360 580410 139369
rect 580354 139295 580410 139304
rect 580356 126268 580408 126274
rect 580356 126210 580408 126216
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 579620 100700 579672 100706
rect 579620 100642 579672 100648
rect 579632 99521 579660 100642
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 580264 87644 580316 87650
rect 580264 87586 580316 87592
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 574744 3868 574796 3874
rect 574744 3810 574796 3816
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 577424 480 577452 3810
rect 578620 480 578648 16546
rect 580276 6633 580304 87586
rect 580368 46345 580396 126210
rect 580460 86193 580488 289031
rect 580552 219065 580580 370534
rect 580724 290488 580776 290494
rect 580724 290430 580776 290436
rect 580630 286376 580686 286385
rect 580630 286311 580686 286320
rect 580538 219056 580594 219065
rect 580538 218991 580594 219000
rect 580644 165889 580672 286311
rect 580736 245585 580764 290430
rect 580722 245576 580778 245585
rect 580722 245511 580778 245520
rect 580630 165880 580686 165889
rect 580630 165815 580686 165824
rect 580446 86184 580502 86193
rect 580446 86119 580502 86128
rect 580354 46336 580410 46345
rect 580354 46271 580410 46280
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3422 579944 3478 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2778 527856 2834 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 7562 381520 7618 381576
rect 4802 380160 4858 380216
rect 46202 389816 46258 389872
rect 90362 403552 90418 403608
rect 40038 378664 40094 378720
rect 169758 377304 169814 377360
rect 104898 374584 104954 374640
rect 3422 371320 3478 371376
rect 227718 367648 227774 367704
rect 226982 367512 227038 367568
rect 224222 363568 224278 363624
rect 3422 358400 3478 358456
rect 3330 345344 3386 345400
rect 220726 322088 220782 322144
rect 217966 321952 218022 322008
rect 213734 321816 213790 321872
rect 213642 321544 213698 321600
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 43442 291216 43498 291272
rect 7562 289040 7618 289096
rect 3514 267144 3570 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3238 162832 3294 162888
rect 4158 237496 4214 237552
rect 3514 201864 3570 201920
rect 3514 188808 3570 188864
rect 3422 149776 3478 149832
rect 2870 136720 2926 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 34518 236544 34574 236600
rect 3422 6432 3478 6488
rect 25502 226888 25558 226944
rect 44178 233824 44234 233880
rect 51078 231104 51134 231160
rect 57978 225528 58034 225584
rect 62118 200640 62174 200696
rect 71042 229744 71098 229800
rect 66258 196560 66314 196616
rect 69018 213152 69074 213208
rect 71778 228248 71834 228304
rect 82818 222808 82874 222864
rect 93858 224168 93914 224224
rect 97998 233960 98054 234016
rect 102138 199280 102194 199336
rect 104898 203496 104954 203552
rect 110418 229880 110474 229936
rect 114558 220224 114614 220280
rect 186962 289176 187018 289232
rect 118790 182824 118846 182880
rect 131118 221448 131174 221504
rect 138018 232464 138074 232520
rect 152462 235184 152518 235240
rect 142158 207576 142214 207632
rect 143630 193840 143686 193896
rect 144918 188264 144974 188320
rect 155222 231376 155278 231432
rect 158718 224304 158774 224360
rect 173898 236816 173954 236872
rect 169758 236680 169814 236736
rect 176658 236952 176714 237008
rect 184938 237224 184994 237280
rect 188342 237904 188398 237960
rect 206282 291352 206338 291408
rect 201498 237088 201554 237144
rect 209686 238448 209742 238504
rect 209042 237768 209098 237824
rect 208398 231240 208454 231296
rect 209870 224440 209926 224496
rect 210698 235864 210754 235920
rect 210698 233824 210754 233880
rect 212170 318416 212226 318472
rect 212078 318144 212134 318200
rect 211986 307128 212042 307184
rect 211066 235864 211122 235920
rect 212354 318280 212410 318336
rect 212170 237768 212226 237824
rect 212446 318008 212502 318064
rect 211986 236408 212042 236464
rect 213274 241032 213330 241088
rect 213550 314336 213606 314392
rect 213090 225528 213146 225584
rect 212538 221584 212594 221640
rect 213642 240488 213698 240544
rect 215114 316648 215170 316704
rect 213734 235728 213790 235784
rect 213642 228248 213698 228304
rect 213734 226888 213790 226944
rect 214470 306992 214526 307048
rect 214838 309712 214894 309768
rect 213826 223488 213882 223544
rect 213826 222808 213882 222864
rect 217782 316512 217838 316568
rect 217598 315288 217654 315344
rect 216218 314200 216274 314256
rect 215206 309848 215262 309904
rect 214838 236544 214894 236600
rect 214838 229880 214894 229936
rect 215666 240216 215722 240272
rect 214746 224848 214802 224904
rect 215206 224848 215262 224904
rect 214746 224168 214802 224224
rect 215758 239944 215814 240000
rect 215758 238992 215814 239048
rect 215942 241032 215998 241088
rect 215942 240216 215998 240272
rect 215666 231104 215722 231160
rect 216494 314064 216550 314120
rect 216126 238992 216182 239048
rect 216310 239944 216366 240000
rect 216218 236952 216274 237008
rect 216586 313928 216642 313984
rect 217138 240624 217194 240680
rect 216586 238040 216642 238096
rect 216494 237224 216550 237280
rect 217506 240896 217562 240952
rect 217506 240624 217562 240680
rect 217598 240352 217654 240408
rect 217414 240216 217470 240272
rect 217322 238720 217378 238776
rect 217138 232464 217194 232520
rect 217322 235592 217378 235648
rect 217230 229744 217286 229800
rect 216678 226888 216734 226944
rect 217874 314472 217930 314528
rect 220634 321680 220690 321736
rect 217598 231376 217654 231432
rect 218702 240624 218758 240680
rect 219254 316920 219310 316976
rect 220450 312432 220506 312488
rect 219162 238992 219218 239048
rect 219438 238176 219494 238232
rect 219254 237768 219310 237824
rect 218886 236952 218942 237008
rect 220082 241168 220138 241224
rect 220082 240488 220138 240544
rect 220358 240488 220414 240544
rect 220358 240216 220414 240272
rect 219990 237904 220046 237960
rect 220450 238176 220506 238232
rect 221922 318688 221978 318744
rect 220726 239536 220782 239592
rect 220910 240216 220966 240272
rect 221186 238584 221242 238640
rect 225602 362208 225658 362264
rect 225234 329024 225290 329080
rect 224590 289992 224646 290048
rect 226430 320728 226486 320784
rect 226430 291080 226486 291136
rect 227626 291080 227682 291136
rect 227626 289856 227682 289912
rect 228730 291488 228786 291544
rect 231122 371592 231178 371648
rect 224958 289584 225014 289640
rect 233054 289720 233110 289776
rect 235630 289720 235686 289776
rect 237378 369960 237434 370016
rect 238666 306312 238722 306368
rect 238850 315424 238906 315480
rect 238666 296792 238722 296848
rect 238666 296656 238722 296712
rect 239034 293120 239090 293176
rect 238666 290264 238722 290320
rect 240414 370368 240470 370424
rect 240230 370096 240286 370152
rect 241610 320592 241666 320648
rect 241610 293256 241666 293312
rect 242714 294752 242770 294808
rect 242990 321000 243046 321056
rect 244370 319368 244426 319424
rect 247130 321272 247186 321328
rect 247222 314608 247278 314664
rect 248418 321136 248474 321192
rect 251178 374040 251234 374096
rect 249890 368600 249946 368656
rect 249614 289992 249670 290048
rect 250718 289992 250774 290048
rect 235906 289584 235962 289640
rect 251270 368872 251326 368928
rect 251362 367784 251418 367840
rect 251086 289720 251142 289776
rect 250994 289584 251050 289640
rect 252650 320864 252706 320920
rect 252650 292032 252706 292088
rect 253938 369008 253994 369064
rect 254122 368736 254178 368792
rect 254030 320456 254086 320512
rect 254214 319504 254270 319560
rect 256514 289992 256570 290048
rect 256238 289720 256294 289776
rect 256514 289756 256516 289776
rect 256516 289756 256568 289776
rect 256568 289756 256570 289776
rect 256514 289720 256570 289756
rect 256790 345616 256846 345672
rect 256974 319640 257030 319696
rect 260930 319776 260986 319832
rect 263598 372816 263654 372872
rect 264334 291352 264390 291408
rect 264978 372680 265034 372736
rect 252558 289584 252614 289640
rect 256606 289584 256662 289640
rect 265898 291216 265954 291272
rect 263874 289584 263930 289640
rect 264978 289584 265034 289640
rect 265162 289312 265218 289368
rect 267554 272448 267610 272504
rect 267646 250416 267702 250472
rect 267554 244160 267610 244216
rect 267554 244024 267610 244080
rect 267554 241576 267610 241632
rect 222290 241304 222346 241360
rect 267922 246200 267978 246256
rect 267830 243480 267886 243536
rect 267462 241168 267518 241224
rect 267646 241068 267648 241088
rect 267648 241068 267700 241088
rect 267700 241068 267702 241088
rect 267646 241032 267702 241068
rect 222290 240252 222292 240272
rect 222292 240252 222344 240272
rect 222344 240252 222346 240272
rect 222290 240216 222346 240252
rect 222290 240080 222346 240136
rect 222198 239128 222254 239184
rect 222382 236272 222438 236328
rect 222750 239708 222752 239728
rect 222752 239708 222804 239728
rect 222804 239708 222806 239728
rect 222750 239672 222806 239708
rect 223072 239842 223128 239898
rect 223118 239692 223174 239728
rect 223118 239672 223120 239692
rect 223120 239672 223172 239692
rect 223172 239672 223174 239692
rect 222612 239400 222668 239456
rect 222934 239400 222990 239456
rect 222842 239264 222898 239320
rect 222842 238856 222898 238912
rect 222842 237768 222898 237824
rect 223394 239692 223450 239728
rect 223394 239672 223396 239692
rect 223396 239672 223448 239692
rect 223448 239672 223450 239692
rect 223302 239400 223358 239456
rect 223210 239128 223266 239184
rect 223578 239536 223634 239592
rect 223486 238448 223542 238504
rect 223670 237768 223726 237824
rect 223854 239692 223910 239728
rect 223854 239672 223856 239692
rect 223856 239672 223908 239692
rect 223908 239672 223910 239692
rect 224176 239842 224232 239898
rect 224314 239708 224316 239728
rect 224316 239708 224368 239728
rect 224368 239708 224370 239728
rect 224314 239672 224370 239708
rect 223946 239536 224002 239592
rect 223762 236272 223818 236328
rect 224590 239536 224646 239592
rect 224590 238584 224646 238640
rect 224498 238312 224554 238368
rect 224038 235728 224094 235784
rect 223762 220768 223818 220824
rect 224038 219272 224094 219328
rect 224590 236136 224646 236192
rect 224866 237632 224922 237688
rect 224498 220768 224554 220824
rect 224498 220496 224554 220552
rect 225188 239808 225244 239864
rect 225326 239572 225328 239592
rect 225328 239572 225380 239592
rect 225380 239572 225382 239592
rect 225326 239536 225382 239572
rect 225510 238992 225566 239048
rect 225050 236408 225106 236464
rect 224958 236136 225014 236192
rect 225234 220632 225290 220688
rect 226016 239808 226072 239864
rect 226062 239672 226118 239728
rect 226384 239808 226440 239864
rect 226982 239808 227038 239864
rect 227120 239808 227176 239864
rect 227304 239842 227360 239898
rect 227672 239842 227728 239898
rect 226154 238448 226210 238504
rect 225878 235864 225934 235920
rect 226706 239672 226762 239728
rect 226890 239708 226892 239728
rect 226892 239708 226944 239728
rect 226944 239708 226946 239728
rect 226890 239672 226946 239708
rect 226522 238448 226578 238504
rect 226614 238040 226670 238096
rect 226798 238720 226854 238776
rect 226798 238176 226854 238232
rect 227948 239808 228004 239864
rect 227258 239556 227314 239592
rect 227258 239536 227260 239556
rect 227260 239536 227312 239556
rect 227312 239536 227314 239556
rect 227258 237904 227314 237960
rect 227626 239672 227682 239728
rect 226982 199416 227038 199472
rect 226338 156576 226394 156632
rect 227718 239572 227720 239592
rect 227720 239572 227772 239592
rect 227772 239572 227774 239592
rect 227718 239536 227774 239572
rect 228500 239808 228556 239864
rect 228776 239808 228832 239864
rect 229052 239844 229054 239864
rect 229054 239844 229106 239864
rect 229106 239844 229108 239864
rect 229052 239808 229108 239844
rect 227902 238856 227958 238912
rect 227718 238720 227774 238776
rect 227994 238040 228050 238096
rect 227994 236000 228050 236056
rect 228178 239400 228234 239456
rect 228362 239400 228418 239456
rect 228914 239672 228970 239728
rect 229328 239808 229384 239864
rect 229006 238856 229062 238912
rect 229006 238604 229062 238640
rect 229006 238584 229008 238604
rect 229008 238584 229060 238604
rect 229060 238584 229062 238604
rect 228914 238176 228970 238232
rect 228822 237904 228878 237960
rect 228730 236544 228786 236600
rect 228270 220768 228326 220824
rect 227994 219136 228050 219192
rect 229466 239400 229522 239456
rect 229466 239128 229522 239184
rect 229466 238584 229522 238640
rect 229742 239148 229798 239184
rect 229742 239128 229744 239148
rect 229744 239128 229796 239148
rect 229796 239128 229798 239148
rect 229650 237360 229706 237416
rect 230202 239672 230258 239728
rect 230386 239708 230388 239728
rect 230388 239708 230440 239728
rect 230440 239708 230442 239728
rect 230110 238720 230166 238776
rect 230110 238176 230166 238232
rect 228730 220768 228786 220824
rect 228730 219816 228786 219872
rect 230386 239672 230442 239708
rect 230386 239572 230388 239592
rect 230388 239572 230440 239592
rect 230440 239572 230442 239592
rect 230386 239536 230442 239572
rect 230386 239128 230442 239184
rect 230754 239672 230810 239728
rect 231168 239808 231224 239864
rect 230662 237496 230718 237552
rect 231214 239672 231270 239728
rect 231306 239572 231308 239592
rect 231308 239572 231360 239592
rect 231360 239572 231362 239592
rect 231306 239536 231362 239572
rect 231490 238720 231546 238776
rect 231996 239808 232052 239864
rect 232640 239842 232696 239898
rect 232916 239842 232972 239898
rect 231674 238040 231730 238096
rect 231950 237904 232006 237960
rect 232594 239536 232650 239592
rect 232870 239536 232926 239592
rect 232042 222128 232098 222184
rect 232870 222128 232926 222184
rect 233652 239808 233708 239864
rect 233928 239842 233984 239898
rect 233146 239692 233202 239728
rect 233146 239672 233148 239692
rect 233148 239672 233200 239692
rect 233200 239672 233202 239692
rect 233330 238584 233386 238640
rect 233514 235320 233570 235376
rect 233698 239536 233754 239592
rect 234296 239808 234352 239864
rect 234250 238584 234306 238640
rect 234664 239808 234720 239864
rect 234618 239572 234620 239592
rect 234620 239572 234672 239592
rect 234672 239572 234674 239592
rect 234618 239536 234674 239572
rect 234434 236952 234490 237008
rect 234618 238584 234674 238640
rect 233606 224848 233662 224904
rect 234894 234776 234950 234832
rect 234802 234504 234858 234560
rect 235952 239808 236008 239864
rect 235722 239672 235778 239728
rect 235630 236680 235686 236736
rect 235998 239672 236054 239728
rect 236596 239808 236652 239864
rect 236964 239842 237020 239898
rect 236182 239128 236238 239184
rect 235262 218048 235318 218104
rect 236458 239536 236514 239592
rect 236642 238040 236698 238096
rect 236550 237224 236606 237280
rect 237286 239672 237342 239728
rect 238160 239808 238216 239864
rect 237930 239264 237986 239320
rect 237378 222128 237434 222184
rect 238206 237088 238262 237144
rect 237930 231240 237986 231296
rect 238390 239672 238446 239728
rect 238712 239808 238768 239864
rect 239264 239808 239320 239864
rect 238574 239400 238630 239456
rect 238850 239264 238906 239320
rect 238482 222128 238538 222184
rect 239218 239708 239220 239728
rect 239220 239708 239272 239728
rect 239272 239708 239274 239728
rect 239218 239672 239274 239708
rect 239218 239264 239274 239320
rect 239494 237904 239550 237960
rect 238850 221720 238906 221776
rect 240046 239536 240102 239592
rect 240644 239842 240700 239898
rect 241334 239556 241390 239592
rect 241334 239536 241336 239556
rect 241336 239536 241388 239556
rect 241388 239536 241390 239556
rect 241748 239808 241804 239864
rect 241610 235864 241666 235920
rect 242346 239808 242402 239864
rect 242484 239808 242540 239864
rect 241978 239128 242034 239184
rect 242760 239808 242816 239864
rect 242530 239692 242586 239728
rect 242530 239672 242532 239692
rect 242532 239672 242584 239692
rect 242584 239672 242586 239692
rect 242438 238584 242494 238640
rect 242346 236680 242402 236736
rect 243036 239808 243092 239864
rect 242898 239536 242954 239592
rect 243174 239536 243230 239592
rect 243358 239400 243414 239456
rect 244278 238584 244334 238640
rect 244830 238584 244886 238640
rect 245198 239692 245254 239728
rect 245198 239672 245200 239692
rect 245200 239672 245252 239692
rect 245252 239672 245254 239692
rect 245198 239556 245254 239592
rect 245198 239536 245200 239556
rect 245200 239536 245252 239556
rect 245252 239536 245254 239556
rect 245474 238584 245530 238640
rect 246210 239828 246266 239864
rect 246210 239808 246212 239828
rect 246212 239808 246264 239828
rect 246264 239808 246266 239828
rect 245566 223080 245622 223136
rect 244922 220768 244978 220824
rect 246026 239536 246082 239592
rect 246762 239672 246818 239728
rect 246762 234504 246818 234560
rect 246946 238584 247002 238640
rect 247820 239808 247876 239864
rect 247866 239708 247868 239728
rect 247868 239708 247920 239728
rect 247920 239708 247922 239728
rect 247866 239672 247922 239708
rect 248050 239672 248106 239728
rect 248050 239400 248106 239456
rect 248418 238584 248474 238640
rect 248602 238584 248658 238640
rect 248878 239572 248880 239592
rect 248880 239572 248932 239592
rect 248932 239572 248934 239592
rect 248878 239536 248934 239572
rect 249246 239672 249302 239728
rect 249752 239808 249808 239864
rect 249338 239400 249394 239456
rect 249522 239536 249578 239592
rect 249614 236136 249670 236192
rect 250074 239400 250130 239456
rect 250350 239692 250406 239728
rect 250350 239672 250352 239692
rect 250352 239672 250404 239692
rect 250404 239672 250406 239692
rect 250856 239808 250912 239864
rect 250534 237904 250590 237960
rect 251408 239808 251464 239864
rect 251960 239808 252016 239864
rect 250626 237224 250682 237280
rect 250810 236136 250866 236192
rect 251086 238584 251142 238640
rect 250994 226208 251050 226264
rect 251638 239536 251694 239592
rect 251822 235320 251878 235376
rect 252098 233688 252154 233744
rect 252466 239536 252522 239592
rect 252282 221584 252338 221640
rect 252650 239692 252706 239728
rect 252650 239672 252652 239692
rect 252652 239672 252704 239692
rect 252704 239672 252706 239692
rect 252650 239128 252706 239184
rect 252926 239536 252982 239592
rect 253110 239708 253112 239728
rect 253112 239708 253164 239728
rect 253164 239708 253166 239728
rect 253110 239672 253166 239708
rect 253340 239808 253396 239864
rect 253386 239536 253442 239592
rect 253478 239128 253534 239184
rect 253110 238584 253166 238640
rect 253202 227160 253258 227216
rect 253754 239692 253810 239728
rect 253754 239672 253756 239692
rect 253756 239672 253808 239692
rect 253808 239672 253810 239692
rect 253754 239536 253810 239592
rect 253662 228656 253718 228712
rect 254168 239808 254224 239864
rect 254536 239808 254592 239864
rect 253846 233144 253902 233200
rect 254582 239536 254638 239592
rect 254674 235864 254730 235920
rect 255180 239808 255236 239864
rect 255042 239572 255044 239592
rect 255044 239572 255096 239592
rect 255096 239572 255098 239592
rect 255042 239536 255098 239572
rect 255042 239400 255098 239456
rect 254950 236000 255006 236056
rect 255226 239672 255282 239728
rect 255594 239572 255596 239592
rect 255596 239572 255648 239592
rect 255648 239572 255650 239592
rect 255226 237904 255282 237960
rect 255134 223760 255190 223816
rect 255594 239536 255650 239572
rect 255502 237904 255558 237960
rect 255410 237632 255466 237688
rect 255318 236952 255374 237008
rect 256652 239808 256708 239864
rect 256146 239400 256202 239456
rect 256330 239572 256332 239592
rect 256332 239572 256384 239592
rect 256384 239572 256386 239592
rect 256330 239536 256386 239572
rect 256514 239672 256570 239728
rect 255686 236544 255742 236600
rect 256974 239672 257030 239728
rect 256790 233824 256846 233880
rect 257480 239842 257536 239898
rect 257158 235184 257214 235240
rect 257940 239842 257996 239898
rect 258216 239842 258272 239898
rect 258078 239672 258134 239728
rect 258262 239672 258318 239728
rect 258584 239808 258640 239864
rect 257894 239536 257950 239592
rect 257526 228520 257582 228576
rect 257986 236680 258042 236736
rect 258078 235728 258134 235784
rect 258446 239672 258502 239728
rect 258354 235184 258410 235240
rect 257986 229608 258042 229664
rect 258078 204856 258134 204912
rect 258814 239264 258870 239320
rect 258722 238040 258778 238096
rect 259136 239808 259192 239864
rect 259090 239572 259092 239592
rect 259092 239572 259144 239592
rect 259144 239572 259146 239592
rect 259090 239536 259146 239572
rect 259182 239400 259238 239456
rect 258998 239128 259054 239184
rect 259090 230016 259146 230072
rect 258998 229880 259054 229936
rect 259596 239808 259652 239864
rect 259458 236816 259514 236872
rect 259366 218048 259422 218104
rect 259642 239672 259698 239728
rect 260424 239808 260480 239864
rect 259642 237088 259698 237144
rect 260102 239556 260158 239592
rect 260102 239536 260104 239556
rect 260104 239536 260156 239556
rect 260156 239536 260158 239556
rect 260470 239264 260526 239320
rect 260378 237496 260434 237552
rect 260102 234368 260158 234424
rect 260010 234232 260066 234288
rect 260102 200640 260158 200696
rect 260930 239536 260986 239592
rect 260654 231784 260710 231840
rect 261022 231648 261078 231704
rect 260746 228928 260802 228984
rect 261896 239842 261952 239898
rect 262080 239842 262136 239898
rect 261666 239264 261722 239320
rect 261850 236680 261906 236736
rect 262586 239828 262642 239864
rect 262586 239808 262588 239828
rect 262588 239808 262640 239828
rect 262640 239808 262642 239828
rect 261942 233008 261998 233064
rect 262126 227432 262182 227488
rect 261850 226072 261906 226128
rect 262494 239672 262550 239728
rect 263000 239896 263056 239898
rect 263000 239844 263002 239896
rect 263002 239844 263054 239896
rect 263054 239844 263056 239896
rect 263000 239842 263056 239844
rect 262586 235184 262642 235240
rect 262678 234096 262734 234152
rect 262494 233960 262550 234016
rect 262402 232736 262458 232792
rect 262954 239672 263010 239728
rect 263506 239692 263562 239728
rect 262770 231376 262826 231432
rect 263046 228928 263102 228984
rect 263506 239672 263508 239692
rect 263508 239672 263560 239692
rect 263560 239672 263562 239692
rect 263828 239808 263884 239864
rect 263230 225664 263286 225720
rect 263598 239128 263654 239184
rect 263782 239264 263838 239320
rect 263874 239128 263930 239184
rect 263874 237632 263930 237688
rect 263874 237360 263930 237416
rect 263414 230152 263470 230208
rect 263874 235456 263930 235512
rect 264058 237904 264114 237960
rect 264472 239808 264528 239864
rect 264334 239672 264390 239728
rect 264242 239536 264298 239592
rect 263966 234504 264022 234560
rect 263782 230288 263838 230344
rect 264334 236544 264390 236600
rect 264610 239672 264666 239728
rect 264518 238448 264574 238504
rect 264932 239842 264988 239898
rect 264610 221176 264666 221232
rect 264978 239708 264980 239728
rect 264980 239708 265032 239728
rect 265032 239708 265034 239728
rect 264978 239672 265034 239708
rect 264886 238448 264942 238504
rect 264978 236680 265034 236736
rect 264886 231512 264942 231568
rect 262218 141344 262274 141400
rect 265346 239692 265402 239728
rect 265346 239672 265348 239692
rect 265348 239672 265400 239692
rect 265400 239672 265402 239692
rect 265714 237904 265770 237960
rect 265944 239808 266000 239864
rect 266588 239808 266644 239864
rect 266082 239672 266138 239728
rect 265714 230968 265770 231024
rect 265622 228792 265678 228848
rect 266542 239672 266598 239728
rect 266634 238040 266690 238096
rect 266266 232328 266322 232384
rect 266542 226888 266598 226944
rect 266818 239708 266820 239728
rect 266820 239708 266872 239728
rect 266872 239708 266874 239728
rect 266818 239672 266874 239708
rect 266818 232464 266874 232520
rect 267094 239808 267150 239864
rect 267554 239980 267556 240000
rect 267556 239980 267608 240000
rect 267608 239980 267610 240000
rect 267554 239944 267610 239980
rect 267646 239808 267702 239864
rect 267554 238312 267610 238368
rect 268014 241032 268070 241088
rect 268474 314608 268530 314664
rect 269302 247560 269358 247616
rect 268842 243616 268898 243672
rect 268750 240760 268806 240816
rect 268842 240216 268898 240272
rect 268658 240080 268714 240136
rect 269118 242256 269174 242312
rect 269118 241168 269174 241224
rect 268934 238584 268990 238640
rect 268658 237224 268714 237280
rect 268566 236952 268622 237008
rect 269486 243752 269542 243808
rect 269118 239536 269174 239592
rect 269118 235592 269174 235648
rect 268474 233688 268530 233744
rect 269486 238176 269542 238232
rect 271142 317192 271198 317248
rect 269118 228248 269174 228304
rect 270130 286456 270186 286512
rect 271142 239672 271198 239728
rect 270958 237496 271014 237552
rect 270038 237088 270094 237144
rect 271602 315832 271658 315888
rect 271786 237632 271842 237688
rect 271510 229744 271566 229800
rect 273902 316784 273958 316840
rect 273902 239400 273958 239456
rect 272522 224032 272578 224088
rect 275466 315016 275522 315072
rect 277582 318588 277584 318608
rect 277584 318588 277636 318608
rect 277636 318588 277638 318608
rect 277582 318552 277638 318588
rect 277766 318144 277822 318200
rect 277766 317736 277822 317792
rect 275374 221312 275430 221368
rect 278410 318588 278412 318608
rect 278412 318588 278464 318608
rect 278464 318588 278466 318608
rect 278410 318552 278466 318588
rect 278410 318416 278466 318472
rect 278410 318008 278466 318064
rect 278318 317328 278374 317384
rect 278042 235456 278098 235512
rect 277306 233144 277362 233200
rect 276662 220088 276718 220144
rect 278134 233144 278190 233200
rect 279974 369824 280030 369880
rect 280710 360204 280712 360224
rect 280712 360204 280764 360224
rect 280764 360204 280766 360224
rect 280710 360168 280766 360204
rect 280710 358828 280766 358864
rect 280710 358808 280712 358828
rect 280712 358808 280764 358828
rect 280764 358808 280766 358828
rect 278410 228656 278466 228712
rect 279514 218728 279570 218784
rect 280158 320320 280214 320376
rect 280158 214512 280214 214568
rect 289082 373224 289138 373280
rect 286782 371728 286838 371784
rect 281262 371456 281318 371512
rect 282090 371320 282146 371376
rect 286046 371320 286102 371376
rect 281262 358808 281318 358864
rect 286046 370232 286102 370288
rect 281998 321952 282054 322008
rect 281906 320184 281962 320240
rect 281906 318144 281962 318200
rect 281998 315152 282054 315208
rect 286184 369824 286240 369880
rect 288254 371592 288310 371648
rect 287058 371456 287114 371512
rect 288024 369824 288080 369880
rect 285218 369552 285274 369608
rect 283654 369416 283710 369472
rect 284482 369416 284538 369472
rect 284942 369416 284998 369472
rect 287426 369416 287482 369472
rect 295614 370368 295670 370424
rect 295614 370096 295670 370152
rect 299570 386280 299626 386336
rect 296718 370096 296774 370152
rect 297960 370096 298016 370152
rect 299110 374176 299166 374232
rect 298926 371320 298982 371376
rect 299662 370368 299718 370424
rect 299662 370096 299718 370152
rect 300168 370096 300224 370152
rect 301502 375672 301558 375728
rect 301042 370504 301098 370560
rect 302606 375536 302662 375592
rect 302330 371592 302386 371648
rect 302974 375536 303030 375592
rect 302882 369688 302938 369744
rect 299294 369416 299350 369472
rect 301778 369416 301834 369472
rect 302882 369416 302938 369472
rect 303480 369688 303536 369744
rect 303986 369416 304042 369472
rect 305642 385600 305698 385656
rect 307942 372544 307998 372600
rect 309598 372544 309654 372600
rect 308402 369688 308458 369744
rect 309368 369688 309424 369744
rect 305458 369416 305514 369472
rect 307298 369416 307354 369472
rect 309874 369416 309930 369472
rect 310104 369416 310160 369472
rect 311898 375400 311954 375456
rect 310978 374040 311034 374096
rect 310702 372544 310758 372600
rect 311714 373224 311770 373280
rect 311346 372544 311402 372600
rect 311346 371864 311402 371920
rect 311714 369688 311770 369744
rect 312450 375400 312506 375456
rect 319534 372816 319590 372872
rect 324962 372680 325018 372736
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580262 458088 580318 458144
rect 579894 431568 579950 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 312818 369552 312874 369608
rect 313278 369552 313334 369608
rect 314520 369552 314576 369608
rect 310978 369416 311034 369472
rect 312082 369416 312138 369472
rect 313922 369416 313978 369472
rect 315026 369416 315082 369472
rect 320914 369416 320970 369472
rect 324226 369416 324282 369472
rect 286552 369280 286608 369336
rect 309000 369280 309056 369336
rect 310104 369280 310160 369336
rect 312312 369280 312368 369336
rect 313416 369280 313472 369336
rect 316728 369280 316784 369336
rect 282366 363568 282422 363624
rect 282274 345616 282330 345672
rect 282182 329024 282238 329080
rect 282274 322088 282330 322144
rect 327722 321272 327778 321328
rect 327538 320864 327594 320920
rect 288024 320728 288080 320784
rect 290140 320728 290196 320784
rect 293452 320728 293508 320784
rect 294096 320728 294152 320784
rect 295384 320728 295440 320784
rect 299432 320728 299488 320784
rect 311208 320728 311264 320784
rect 323352 320728 323408 320784
rect 324456 320728 324512 320784
rect 311944 320592 312000 320648
rect 313140 320592 313196 320648
rect 322800 320592 322856 320648
rect 325008 320592 325064 320648
rect 315072 320456 315128 320512
rect 317648 320456 317704 320512
rect 318844 320456 318900 320512
rect 323904 320456 323960 320512
rect 325560 320456 325616 320512
rect 282964 320320 283020 320376
rect 283240 320320 283296 320376
rect 283792 320320 283848 320376
rect 289680 320320 289736 320376
rect 291060 320320 291116 320376
rect 297684 320320 297740 320376
rect 298052 320320 298108 320376
rect 298604 320320 298660 320376
rect 300628 320320 300684 320376
rect 308908 320320 308964 320376
rect 312220 320320 312276 320376
rect 313232 320320 313288 320376
rect 317096 320320 317152 320376
rect 318752 320320 318808 320376
rect 318936 320320 318992 320376
rect 323168 320320 323224 320376
rect 326664 320320 326720 320376
rect 285172 320184 285228 320240
rect 286460 320184 286516 320240
rect 286644 320184 286700 320240
rect 287380 320184 287436 320240
rect 288116 320184 288172 320240
rect 289036 320184 289092 320240
rect 290324 320184 290380 320240
rect 290968 320184 291024 320240
rect 291336 320184 291392 320240
rect 293544 320184 293600 320240
rect 294188 320184 294244 320240
rect 296856 320184 296912 320240
rect 297776 320184 297832 320240
rect 299340 320184 299396 320240
rect 300996 320184 301052 320240
rect 304216 320184 304272 320240
rect 308448 320184 308504 320240
rect 309920 320184 309976 320240
rect 310840 320184 310896 320240
rect 311668 320184 311724 320240
rect 312404 320184 312460 320240
rect 312956 320184 313012 320240
rect 314336 320184 314392 320240
rect 316268 320184 316324 320240
rect 316544 320184 316600 320240
rect 317280 320184 317336 320240
rect 318384 320184 318440 320240
rect 320132 320184 320188 320240
rect 321420 320184 321476 320240
rect 322064 320184 322120 320240
rect 323076 320184 323132 320240
rect 324272 320184 324328 320240
rect 326112 320184 326168 320240
rect 328550 320728 328606 320784
rect 282274 320048 282330 320104
rect 281446 287000 281502 287056
rect 281446 286320 281502 286376
rect 280986 228520 281042 228576
rect 281170 214512 281226 214568
rect 281170 213832 281226 213888
rect 282366 319232 282422 319288
rect 282872 320048 282928 320104
rect 283056 320048 283112 320104
rect 282458 318688 282514 318744
rect 282550 318552 282606 318608
rect 282550 318144 282606 318200
rect 282366 317872 282422 317928
rect 282274 310392 282330 310448
rect 282274 309848 282330 309904
rect 282274 225936 282330 225992
rect 283286 307400 283342 307456
rect 283102 297608 283158 297664
rect 283470 319232 283526 319288
rect 284160 320048 284216 320104
rect 282918 220244 282974 220280
rect 282918 220224 282920 220244
rect 282920 220224 282972 220244
rect 282972 220224 282974 220244
rect 284022 319232 284078 319288
rect 284712 320048 284768 320104
rect 284022 318280 284078 318336
rect 283654 309576 283710 309632
rect 284206 319096 284262 319152
rect 284206 318144 284262 318200
rect 284206 316512 284262 316568
rect 283930 297744 283986 297800
rect 283838 294616 283894 294672
rect 284574 319232 284630 319288
rect 285034 319232 285090 319288
rect 284758 316920 284814 316976
rect 284942 317872 284998 317928
rect 284850 241304 284906 241360
rect 284758 238992 284814 239048
rect 285218 317600 285274 317656
rect 285540 320048 285596 320104
rect 285494 319232 285550 319288
rect 286092 320048 286148 320104
rect 285770 317736 285826 317792
rect 285678 309848 285734 309904
rect 286138 317464 286194 317520
rect 286230 296112 286286 296168
rect 286690 318688 286746 318744
rect 286598 317056 286654 317112
rect 285034 218592 285090 218648
rect 286598 307128 286654 307184
rect 286966 317600 287022 317656
rect 287656 320048 287712 320104
rect 287150 318144 287206 318200
rect 287150 318008 287206 318064
rect 287058 317464 287114 317520
rect 287150 309304 287206 309360
rect 287794 318688 287850 318744
rect 287794 317736 287850 317792
rect 287702 317464 287758 317520
rect 287426 298696 287482 298752
rect 287334 295976 287390 296032
rect 287242 291896 287298 291952
rect 286690 225800 286746 225856
rect 287426 223488 287482 223544
rect 288070 319232 288126 319288
rect 287978 318688 288034 318744
rect 288392 320048 288448 320104
rect 288346 318688 288402 318744
rect 288852 320048 288908 320104
rect 288622 318144 288678 318200
rect 288530 317464 288586 317520
rect 288438 312044 288494 312080
rect 288438 312024 288440 312044
rect 288440 312024 288492 312044
rect 288492 312024 288494 312044
rect 288070 302776 288126 302832
rect 287978 290672 288034 290728
rect 287794 218864 287850 218920
rect 288898 318688 288954 318744
rect 288530 247696 288586 247752
rect 289404 320048 289460 320104
rect 289082 317600 289138 317656
rect 288990 238856 289046 238912
rect 289864 320048 289920 320104
rect 290416 320048 290472 320104
rect 289542 318416 289598 318472
rect 289542 317872 289598 317928
rect 289358 308624 289414 308680
rect 289910 319232 289966 319288
rect 289818 316648 289874 316704
rect 290094 318688 290150 318744
rect 290370 319232 290426 319288
rect 290186 317736 290242 317792
rect 290094 307264 290150 307320
rect 289542 304136 289598 304192
rect 289450 238448 289506 238504
rect 289174 227024 289230 227080
rect 290876 320048 290932 320104
rect 290830 319232 290886 319288
rect 290370 307536 290426 307592
rect 290922 318688 290978 318744
rect 291520 320048 291576 320104
rect 291704 320048 291760 320104
rect 291198 319232 291254 319288
rect 291014 315696 291070 315752
rect 291290 317464 291346 317520
rect 291566 317464 291622 317520
rect 292348 320048 292404 320104
rect 291934 318824 291990 318880
rect 291382 238720 291438 238776
rect 292210 318824 292266 318880
rect 292394 315716 292450 315752
rect 292394 315696 292396 315716
rect 292396 315696 292448 315716
rect 292448 315696 292450 315716
rect 292670 317464 292726 317520
rect 293176 320048 293232 320104
rect 292854 317600 292910 317656
rect 292578 312024 292634 312080
rect 290462 221448 290518 221504
rect 289082 220088 289138 220144
rect 286506 218456 286562 218512
rect 289174 211792 289230 211848
rect 293038 315716 293094 315752
rect 293038 315696 293040 315716
rect 293040 315696 293092 315716
rect 293092 315696 293094 315716
rect 293728 320048 293784 320104
rect 293222 319368 293278 319424
rect 293222 318824 293278 318880
rect 294280 320048 294336 320104
rect 293590 318416 293646 318472
rect 293498 318144 293554 318200
rect 293498 310936 293554 310992
rect 294234 318824 294290 318880
rect 294602 319368 294658 319424
rect 294602 318824 294658 318880
rect 295016 320048 295072 320104
rect 294786 317872 294842 317928
rect 295568 320048 295624 320104
rect 295936 320048 295992 320104
rect 295338 319404 295340 319424
rect 295340 319404 295392 319424
rect 295392 319404 295394 319424
rect 295338 319368 295394 319404
rect 294970 317328 295026 317384
rect 294326 224712 294382 224768
rect 291934 222672 291990 222728
rect 296212 320048 296268 320104
rect 292578 208256 292634 208312
rect 293958 166232 294014 166288
rect 296166 317464 296222 317520
rect 296442 318824 296498 318880
rect 296718 318824 296774 318880
rect 296902 318416 296958 318472
rect 297316 320048 297372 320104
rect 297178 318824 297234 318880
rect 297086 317464 297142 317520
rect 297914 318688 297970 318744
rect 298098 317328 298154 317384
rect 298098 312840 298154 312896
rect 299064 320048 299120 320104
rect 299018 318824 299074 318880
rect 298926 318688 298982 318744
rect 298558 312704 298614 312760
rect 298282 241712 298338 241768
rect 297454 235592 297510 235648
rect 298098 188264 298154 188320
rect 299202 318688 299258 318744
rect 299708 320048 299764 320104
rect 299478 317872 299534 317928
rect 299662 318824 299718 318880
rect 300260 320048 300316 320104
rect 299846 319368 299902 319424
rect 299754 305632 299810 305688
rect 300720 320048 300776 320104
rect 300398 319368 300454 319424
rect 300582 317464 300638 317520
rect 300766 312568 300822 312624
rect 300490 300056 300546 300112
rect 301042 318824 301098 318880
rect 300950 317464 301006 317520
rect 300858 291760 300914 291816
rect 302100 320048 302156 320104
rect 301502 312976 301558 313032
rect 301410 312296 301466 312352
rect 302146 319368 302202 319424
rect 301318 300328 301374 300384
rect 302744 320048 302800 320104
rect 302330 318280 302386 318336
rect 302514 319368 302570 319424
rect 302974 318688 303030 318744
rect 302974 318416 303030 318472
rect 302238 231104 302294 231160
rect 302054 227568 302110 227624
rect 302974 312160 303030 312216
rect 302974 229880 303030 229936
rect 303848 320048 303904 320104
rect 303710 318144 303766 318200
rect 304400 320048 304456 320104
rect 303342 315424 303398 315480
rect 303710 233144 303766 233200
rect 303434 219136 303490 219192
rect 304170 319368 304226 319424
rect 305136 320048 305192 320104
rect 304722 317600 304778 317656
rect 304998 318824 305054 318880
rect 305090 317600 305146 317656
rect 305274 317736 305330 317792
rect 305182 317464 305238 317520
rect 306056 320048 306112 320104
rect 306240 320048 306296 320104
rect 305550 317464 305606 317520
rect 305734 319368 305790 319424
rect 305918 317872 305974 317928
rect 306884 320048 306940 320104
rect 306102 318960 306158 319016
rect 306286 319368 306342 319424
rect 306102 229200 306158 229256
rect 305274 226208 305330 226264
rect 304998 213152 305054 213208
rect 307160 320048 307216 320104
rect 306838 319368 306894 319424
rect 306746 319232 306802 319288
rect 307022 317464 307078 317520
rect 307114 311344 307170 311400
rect 307620 320048 307676 320104
rect 307482 319540 307484 319560
rect 307484 319540 307536 319560
rect 307536 319540 307538 319560
rect 307482 319504 307538 319540
rect 307574 317600 307630 317656
rect 308172 320048 308228 320104
rect 307850 318552 307906 318608
rect 308494 319368 308550 319424
rect 308494 317736 308550 317792
rect 308034 311208 308090 311264
rect 308770 319504 308826 319560
rect 308678 317872 308734 317928
rect 309736 320048 309792 320104
rect 310104 320048 310160 320104
rect 309322 319368 309378 319424
rect 309230 319232 309286 319288
rect 308678 311752 308734 311808
rect 308770 311616 308826 311672
rect 309506 319504 309562 319560
rect 309690 319504 309746 319560
rect 309782 318960 309838 319016
rect 308862 223216 308918 223272
rect 308586 222808 308642 222864
rect 309966 311480 310022 311536
rect 309874 253952 309930 254008
rect 309874 230016 309930 230072
rect 310472 320048 310528 320104
rect 310748 320048 310804 320104
rect 310150 319232 310206 319288
rect 310610 319232 310666 319288
rect 310794 319776 310850 319832
rect 310886 319368 310942 319424
rect 310794 318960 310850 319016
rect 310242 311072 310298 311128
rect 311162 312024 311218 312080
rect 311346 319504 311402 319560
rect 311346 319232 311402 319288
rect 311162 235320 311218 235376
rect 310058 222944 310114 223000
rect 312496 320048 312552 320104
rect 312266 319796 312322 319832
rect 312266 319776 312268 319796
rect 312268 319776 312320 319796
rect 312320 319776 312322 319796
rect 311990 318824 312046 318880
rect 311714 317464 311770 317520
rect 311714 314744 311770 314800
rect 313186 319776 313242 319832
rect 312450 319504 312506 319560
rect 312634 319640 312690 319696
rect 312634 318960 312690 319016
rect 313002 319504 313058 319560
rect 313002 318280 313058 318336
rect 312910 315560 312966 315616
rect 312726 309440 312782 309496
rect 312634 233824 312690 233880
rect 313278 319640 313334 319696
rect 313462 319640 313518 319696
rect 313186 300192 313242 300248
rect 313830 319640 313886 319696
rect 314106 315016 314162 315072
rect 313554 294480 313610 294536
rect 313278 222964 313334 223000
rect 313278 222944 313280 222964
rect 313280 222944 313332 222964
rect 313332 222944 313334 222964
rect 311438 221584 311494 221640
rect 311162 192480 311218 192536
rect 314382 317464 314438 317520
rect 314198 310120 314254 310176
rect 314290 309984 314346 310040
rect 314106 232464 314162 232520
rect 314750 319640 314806 319696
rect 314658 319232 314714 319288
rect 314566 317736 314622 317792
rect 315808 320048 315864 320104
rect 315992 320048 316048 320104
rect 316176 320048 316232 320104
rect 315578 310256 315634 310312
rect 315578 238040 315634 238096
rect 315302 232872 315358 232928
rect 315946 319504 316002 319560
rect 316314 319640 316370 319696
rect 316314 318960 316370 319016
rect 317188 320048 317244 320104
rect 317464 320048 317520 320104
rect 317050 319776 317106 319832
rect 316498 319504 316554 319560
rect 316774 319504 316830 319560
rect 316406 287680 316462 287736
rect 316682 235728 316738 235784
rect 317234 319504 317290 319560
rect 317326 318572 317382 318608
rect 317326 318552 317328 318572
rect 317328 318552 317380 318572
rect 317380 318552 317382 318572
rect 317740 319878 317796 319934
rect 317602 319640 317658 319696
rect 318108 320048 318164 320104
rect 318568 320048 318624 320104
rect 317878 319504 317934 319560
rect 318062 319640 318118 319696
rect 318062 319368 318118 319424
rect 317694 308488 317750 308544
rect 317602 290400 317658 290456
rect 318430 319640 318486 319696
rect 318522 319368 318578 319424
rect 318338 317464 318394 317520
rect 318062 224576 318118 224632
rect 318246 224304 318302 224360
rect 318706 319640 318762 319696
rect 318614 318280 318670 318336
rect 319212 320048 319268 320104
rect 319396 320048 319452 320104
rect 318982 319504 319038 319560
rect 318614 304000 318670 304056
rect 319166 319504 319222 319560
rect 319074 318960 319130 319016
rect 319258 318416 319314 318472
rect 319166 318144 319222 318200
rect 319856 320048 319912 320104
rect 320040 320048 320096 320104
rect 319672 319776 319728 319832
rect 319534 319640 319590 319696
rect 319626 319368 319682 319424
rect 319810 319640 319866 319696
rect 319810 319504 319866 319560
rect 319994 319776 320050 319832
rect 319902 308352 319958 308408
rect 316130 152360 316186 152416
rect 319626 244024 319682 244080
rect 320408 320048 320464 320104
rect 320638 319660 320694 319696
rect 320638 319640 320640 319660
rect 320640 319640 320692 319660
rect 320692 319640 320694 319660
rect 320638 319504 320694 319560
rect 320638 316784 320694 316840
rect 320638 290808 320694 290864
rect 321144 320048 321200 320104
rect 321512 320048 321568 320104
rect 321098 319504 321154 319560
rect 321282 319640 321338 319696
rect 320914 236680 320970 236736
rect 320822 232736 320878 232792
rect 322156 320048 322212 320104
rect 322248 319878 322304 319934
rect 322110 319640 322166 319696
rect 322018 319504 322074 319560
rect 322616 320048 322672 320104
rect 321374 241984 321430 242040
rect 322386 319504 322442 319560
rect 322662 319776 322718 319832
rect 322202 239264 322258 239320
rect 322478 317872 322534 317928
rect 322294 227432 322350 227488
rect 322386 226072 322442 226128
rect 322846 319504 322902 319560
rect 323628 320048 323684 320104
rect 323398 319504 323454 319560
rect 324088 320048 324144 320104
rect 323214 244840 323270 244896
rect 323122 243616 323178 243672
rect 322662 230152 322718 230208
rect 323674 319640 323730 319696
rect 323950 319368 324006 319424
rect 323674 316104 323730 316160
rect 324226 319232 324282 319288
rect 323582 241168 323638 241224
rect 324502 319640 324558 319696
rect 324318 243888 324374 243944
rect 323950 241848 324006 241904
rect 324686 318960 324742 319016
rect 325192 319878 325248 319934
rect 324686 258712 324742 258768
rect 324594 246200 324650 246256
rect 325238 319368 325294 319424
rect 325146 241032 325202 241088
rect 325054 239128 325110 239184
rect 324962 237904 325018 237960
rect 325422 318280 325478 318336
rect 325422 318008 325478 318064
rect 325974 317736 326030 317792
rect 326388 320048 326444 320104
rect 326940 320048 326996 320104
rect 326986 319776 327042 319832
rect 326710 319504 326766 319560
rect 326526 318552 326582 318608
rect 326618 318416 326674 318472
rect 326618 317600 326674 317656
rect 326802 317600 326858 317656
rect 326894 317192 326950 317248
rect 326894 316648 326950 316704
rect 326986 272448 327042 272504
rect 326618 271088 326674 271144
rect 325974 250416 326030 250472
rect 325882 244976 325938 245032
rect 325790 243752 325846 243808
rect 327078 224168 327134 224224
rect 324962 199280 325018 199336
rect 327262 318552 327318 318608
rect 327722 317736 327778 317792
rect 327354 317464 327410 317520
rect 327262 258848 327318 258904
rect 327722 240896 327778 240952
rect 327998 247560 328054 247616
rect 327906 240760 327962 240816
rect 327446 234096 327502 234152
rect 327722 234096 327778 234152
rect 328366 231784 328422 231840
rect 328366 231104 328422 231160
rect 328642 319912 328698 319968
rect 328734 231784 328790 231840
rect 331862 370232 331918 370288
rect 330206 320456 330262 320512
rect 329194 318008 329250 318064
rect 329286 231784 329342 231840
rect 328918 231648 328974 231704
rect 328734 231376 328790 231432
rect 328642 226888 328698 226944
rect 330482 234368 330538 234424
rect 330114 234232 330170 234288
rect 330022 232600 330078 232656
rect 329838 186904 329894 186960
rect 331494 319368 331550 319424
rect 331678 318144 331734 318200
rect 331402 233960 331458 234016
rect 331494 231512 331550 231568
rect 334622 369824 334678 369880
rect 332782 321000 332838 321056
rect 332690 318824 332746 318880
rect 332046 317464 332102 317520
rect 334438 320592 334494 320648
rect 334346 320184 334402 320240
rect 334254 319232 334310 319288
rect 334162 318960 334218 319016
rect 333058 231104 333114 231160
rect 334346 232328 334402 232384
rect 334254 230288 334310 230344
rect 335358 321544 335414 321600
rect 334714 318416 334770 318472
rect 334806 230288 334862 230344
rect 334806 229744 334862 229800
rect 335450 321136 335506 321192
rect 335634 319096 335690 319152
rect 335634 228928 335690 228984
rect 335910 234504 335966 234560
rect 335726 228248 335782 228304
rect 335450 225528 335506 225584
rect 333886 6024 333942 6080
rect 336646 234504 336702 234560
rect 336646 233824 336702 233880
rect 336922 229880 336978 229936
rect 336738 197920 336794 197976
rect 338394 320048 338450 320104
rect 338670 320320 338726 320376
rect 347778 167592 347834 167648
rect 358082 314880 358138 314936
rect 354678 236680 354734 236736
rect 355322 236680 355378 236736
rect 350538 178608 350594 178664
rect 354678 202136 354734 202192
rect 475382 317464 475438 317520
rect 365810 138624 365866 138680
rect 373998 314744 374054 314800
rect 378138 312024 378194 312080
rect 379978 3576 380034 3632
rect 383566 3440 383622 3496
rect 401322 6840 401378 6896
rect 404818 6704 404874 6760
rect 418802 283464 418858 283520
rect 418158 156576 418214 156632
rect 434718 253952 434774 254008
rect 426162 6568 426218 6624
rect 436650 6432 436706 6488
rect 440238 229880 440294 229936
rect 440330 6296 440386 6352
rect 447138 168952 447194 169008
rect 449898 151000 449954 151056
rect 456890 15816 456946 15872
rect 465170 6160 465226 6216
rect 471978 146920 472034 146976
rect 474738 25472 474794 25528
rect 488538 316784 488594 316840
rect 483018 234096 483074 234152
rect 486422 3304 486478 3360
rect 569958 316648 570014 316704
rect 490010 231104 490066 231160
rect 508502 311888 508558 311944
rect 502982 233960 503038 234016
rect 507858 232600 507914 232656
rect 514850 190984 514906 191040
rect 517518 189624 517574 189680
rect 523130 228384 523186 228440
rect 525798 225528 525854 225584
rect 528558 10240 528614 10296
rect 532698 233824 532754 233880
rect 538218 316104 538274 316160
rect 536102 229744 536158 229800
rect 546498 182824 546554 182880
rect 555422 232464 555478 232520
rect 557538 228248 557594 228304
rect 562322 226888 562378 226944
rect 574742 302232 574798 302288
rect 580262 371728 580318 371784
rect 580170 365064 580226 365120
rect 579618 351872 579674 351928
rect 580170 325216 580226 325272
rect 580170 272176 580226 272232
rect 579802 258848 579858 258904
rect 579986 232328 580042 232384
rect 580170 205672 580226 205728
rect 579618 192480 579674 192536
rect 579710 179152 579766 179208
rect 580170 152632 580226 152688
rect 580446 312024 580502 312080
rect 580446 298696 580502 298752
rect 580446 289040 580502 289096
rect 580354 139304 580410 139360
rect 580262 112784 580318 112840
rect 579618 99456 579674 99512
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 19760 580226 19816
rect 580630 286320 580686 286376
rect 580538 219000 580594 219056
rect 580722 245520 580778 245576
rect 580630 165824 580686 165880
rect 580446 86128 580502 86184
rect 580354 46280 580410 46336
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2773 527914 2839 527917
rect -960 527912 2839 527914
rect -960 527856 2778 527912
rect 2834 527856 2839 527912
rect -960 527854 2839 527856
rect -960 527764 480 527854
rect 2773 527851 2839 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 90357 403610 90423 403613
rect 309174 403610 309180 403612
rect 90357 403608 309180 403610
rect 90357 403552 90362 403608
rect 90418 403552 309180 403608
rect 90357 403550 309180 403552
rect 90357 403547 90423 403550
rect 309174 403548 309180 403550
rect 309244 403548 309250 403612
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect 46197 389874 46263 389877
rect 313406 389874 313412 389876
rect 46197 389872 313412 389874
rect 46197 389816 46202 389872
rect 46258 389816 313412 389872
rect 46197 389814 313412 389816
rect 46197 389811 46263 389814
rect 313406 389812 313412 389814
rect 313476 389812 313482 389876
rect 299565 386338 299631 386341
rect 305494 386338 305500 386340
rect 299565 386336 305500 386338
rect 299565 386280 299570 386336
rect 299626 386280 305500 386336
rect 299565 386278 305500 386280
rect 299565 386275 299631 386278
rect 305494 386276 305500 386278
rect 305564 386276 305570 386340
rect 305637 385658 305703 385661
rect 316718 385658 316724 385660
rect 305637 385656 316724 385658
rect 305637 385600 305642 385656
rect 305698 385600 316724 385656
rect 305637 385598 316724 385600
rect 305637 385595 305703 385598
rect 316718 385596 316724 385598
rect 316788 385596 316794 385660
rect -960 384284 480 384524
rect 7557 381578 7623 381581
rect 314694 381578 314700 381580
rect 7557 381576 314700 381578
rect 7557 381520 7562 381576
rect 7618 381520 314700 381576
rect 7557 381518 314700 381520
rect 7557 381515 7623 381518
rect 314694 381516 314700 381518
rect 314764 381516 314770 381580
rect 4797 380218 4863 380221
rect 313222 380218 313228 380220
rect 4797 380216 313228 380218
rect 4797 380160 4802 380216
rect 4858 380160 313228 380216
rect 4797 380158 313228 380160
rect 4797 380155 4863 380158
rect 313222 380156 313228 380158
rect 313292 380156 313298 380220
rect 40033 378722 40099 378725
rect 309358 378722 309364 378724
rect 40033 378720 309364 378722
rect 40033 378664 40038 378720
rect 40094 378664 309364 378720
rect 40033 378662 309364 378664
rect 40033 378659 40099 378662
rect 309358 378660 309364 378662
rect 309428 378660 309434 378724
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 169753 377362 169819 377365
rect 306414 377362 306420 377364
rect 169753 377360 306420 377362
rect 169753 377304 169758 377360
rect 169814 377304 306420 377360
rect 169753 377302 306420 377304
rect 169753 377299 169819 377302
rect 306414 377300 306420 377302
rect 306484 377300 306490 377364
rect 277894 375668 277900 375732
rect 277964 375730 277970 375732
rect 301497 375730 301563 375733
rect 277964 375728 301563 375730
rect 277964 375672 301502 375728
rect 301558 375672 301563 375728
rect 277964 375670 301563 375672
rect 277964 375668 277970 375670
rect 301497 375667 301563 375670
rect 275318 375532 275324 375596
rect 275388 375594 275394 375596
rect 302601 375594 302667 375597
rect 302969 375594 303035 375597
rect 275388 375592 303035 375594
rect 275388 375536 302606 375592
rect 302662 375536 302974 375592
rect 303030 375536 303035 375592
rect 275388 375534 303035 375536
rect 275388 375532 275394 375534
rect 302601 375531 302667 375534
rect 302969 375531 303035 375534
rect 275134 375396 275140 375460
rect 275204 375458 275210 375460
rect 311893 375458 311959 375461
rect 312445 375458 312511 375461
rect 275204 375456 312511 375458
rect 275204 375400 311898 375456
rect 311954 375400 312450 375456
rect 312506 375400 312511 375456
rect 275204 375398 312511 375400
rect 275204 375396 275210 375398
rect 311893 375395 311959 375398
rect 312445 375395 312511 375398
rect 104893 374642 104959 374645
rect 307702 374642 307708 374644
rect 104893 374640 307708 374642
rect 104893 374584 104898 374640
rect 104954 374584 307708 374640
rect 104893 374582 307708 374584
rect 104893 374579 104959 374582
rect 307702 374580 307708 374582
rect 307772 374580 307778 374644
rect 278078 374172 278084 374236
rect 278148 374234 278154 374236
rect 299105 374234 299171 374237
rect 278148 374232 299171 374234
rect 278148 374176 299110 374232
rect 299166 374176 299171 374232
rect 278148 374174 299171 374176
rect 278148 374172 278154 374174
rect 299105 374171 299171 374174
rect 251173 374098 251239 374101
rect 310973 374098 311039 374101
rect 251173 374096 311039 374098
rect 251173 374040 251178 374096
rect 251234 374040 310978 374096
rect 311034 374040 311039 374096
rect 251173 374038 311039 374040
rect 251173 374035 251239 374038
rect 310973 374035 311039 374038
rect 289077 373282 289143 373285
rect 311709 373282 311775 373285
rect 289077 373280 311775 373282
rect 289077 373224 289082 373280
rect 289138 373224 311714 373280
rect 311770 373224 311775 373280
rect 289077 373222 311775 373224
rect 289077 373219 289143 373222
rect 311709 373219 311775 373222
rect 263593 372874 263659 372877
rect 319529 372874 319595 372877
rect 263593 372872 319595 372874
rect 263593 372816 263598 372872
rect 263654 372816 319534 372872
rect 319590 372816 319595 372872
rect 263593 372814 319595 372816
rect 263593 372811 263659 372814
rect 319529 372811 319595 372814
rect 264973 372738 265039 372741
rect 324957 372738 325023 372741
rect 264973 372736 325023 372738
rect 264973 372680 264978 372736
rect 265034 372680 324962 372736
rect 325018 372680 325023 372736
rect 264973 372678 325023 372680
rect 264973 372675 265039 372678
rect 324957 372675 325023 372678
rect 307518 372540 307524 372604
rect 307588 372602 307594 372604
rect 307937 372602 308003 372605
rect 307588 372600 308003 372602
rect 307588 372544 307942 372600
rect 307998 372544 308003 372600
rect 307588 372542 308003 372544
rect 307588 372540 307594 372542
rect 307937 372539 308003 372542
rect 309358 372540 309364 372604
rect 309428 372602 309434 372604
rect 309593 372602 309659 372605
rect 309428 372600 309659 372602
rect 309428 372544 309598 372600
rect 309654 372544 309659 372600
rect 309428 372542 309659 372544
rect 309428 372540 309434 372542
rect 309593 372539 309659 372542
rect 310697 372602 310763 372605
rect 311341 372602 311407 372605
rect 310697 372600 311407 372602
rect 310697 372544 310702 372600
rect 310758 372544 311346 372600
rect 311402 372544 311407 372600
rect 310697 372542 311407 372544
rect 310697 372539 310763 372542
rect 311341 372539 311407 372542
rect 285622 371860 285628 371924
rect 285692 371922 285698 371924
rect 311341 371922 311407 371925
rect 285692 371920 311407 371922
rect 285692 371864 311346 371920
rect 311402 371864 311407 371920
rect 285692 371862 311407 371864
rect 285692 371860 285698 371862
rect 311341 371859 311407 371862
rect 286777 371786 286843 371789
rect 580257 371786 580323 371789
rect 282870 371784 580323 371786
rect 282870 371728 286782 371784
rect 286838 371728 580262 371784
rect 580318 371728 580323 371784
rect 282870 371726 580323 371728
rect 231117 371650 231183 371653
rect 282870 371650 282930 371726
rect 286777 371723 286843 371726
rect 580257 371723 580323 371726
rect 231117 371648 282930 371650
rect 231117 371592 231122 371648
rect 231178 371592 282930 371648
rect 231117 371590 282930 371592
rect 288249 371650 288315 371653
rect 302325 371650 302391 371653
rect 288249 371648 302391 371650
rect 288249 371592 288254 371648
rect 288310 371592 302330 371648
rect 302386 371592 302391 371648
rect 288249 371590 302391 371592
rect 231117 371587 231183 371590
rect 288249 371587 288315 371590
rect 302325 371587 302391 371590
rect 281257 371514 281323 371517
rect 287053 371514 287119 371517
rect 281257 371512 287119 371514
rect -960 371378 480 371468
rect 281257 371456 281262 371512
rect 281318 371456 287058 371512
rect 287114 371456 287119 371512
rect 281257 371454 287119 371456
rect 281257 371451 281323 371454
rect 287053 371451 287119 371454
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 282085 371378 282151 371381
rect 286041 371378 286107 371381
rect 282085 371376 286107 371378
rect 282085 371320 282090 371376
rect 282146 371320 286046 371376
rect 286102 371320 286107 371376
rect 282085 371318 286107 371320
rect 282085 371315 282151 371318
rect 286041 371315 286107 371318
rect 296478 371316 296484 371380
rect 296548 371378 296554 371380
rect 298921 371378 298987 371381
rect 296548 371376 298987 371378
rect 296548 371320 298926 371376
rect 298982 371320 298987 371376
rect 296548 371318 298987 371320
rect 296548 371316 296554 371318
rect 298921 371315 298987 371318
rect 301037 370562 301103 370565
rect 292530 370560 301103 370562
rect 292530 370504 301042 370560
rect 301098 370504 301103 370560
rect 292530 370502 301103 370504
rect 240409 370426 240475 370429
rect 292530 370426 292590 370502
rect 301037 370499 301103 370502
rect 240409 370424 292590 370426
rect 240409 370368 240414 370424
rect 240470 370368 292590 370424
rect 240409 370366 292590 370368
rect 295609 370426 295675 370429
rect 299657 370426 299723 370429
rect 295609 370424 299723 370426
rect 295609 370368 295614 370424
rect 295670 370368 299662 370424
rect 299718 370368 299723 370424
rect 295609 370366 299723 370368
rect 240409 370363 240475 370366
rect 295609 370363 295675 370366
rect 299657 370363 299723 370366
rect 286041 370290 286107 370293
rect 331857 370290 331923 370293
rect 286041 370288 331923 370290
rect 286041 370232 286046 370288
rect 286102 370232 331862 370288
rect 331918 370232 331923 370288
rect 286041 370230 331923 370232
rect 286041 370227 286107 370230
rect 331857 370227 331923 370230
rect 240225 370154 240291 370157
rect 295609 370154 295675 370157
rect 296713 370154 296779 370157
rect 297955 370154 298021 370157
rect 240225 370152 295675 370154
rect 240225 370096 240230 370152
rect 240286 370096 295614 370152
rect 295670 370096 295675 370152
rect 240225 370094 295675 370096
rect 240225 370091 240291 370094
rect 295609 370091 295675 370094
rect 295750 370152 298021 370154
rect 295750 370096 296718 370152
rect 296774 370096 297960 370152
rect 298016 370096 298021 370152
rect 295750 370094 298021 370096
rect 237373 370018 237439 370021
rect 295750 370018 295810 370094
rect 296713 370091 296779 370094
rect 297955 370091 298021 370094
rect 299657 370154 299723 370157
rect 300163 370154 300229 370157
rect 299657 370152 300229 370154
rect 299657 370096 299662 370152
rect 299718 370096 300168 370152
rect 300224 370096 300229 370152
rect 299657 370094 300229 370096
rect 299657 370091 299723 370094
rect 300163 370091 300229 370094
rect 237373 370016 295810 370018
rect 237373 369960 237378 370016
rect 237434 369960 295810 370016
rect 237373 369958 295810 369960
rect 237373 369955 237439 369958
rect 279969 369882 280035 369885
rect 286179 369882 286245 369885
rect 288019 369884 288085 369885
rect 288014 369882 288020 369884
rect 279969 369880 286245 369882
rect 279969 369824 279974 369880
rect 280030 369824 286184 369880
rect 286240 369824 286245 369880
rect 279969 369822 286245 369824
rect 287892 369822 288020 369882
rect 288084 369882 288090 369884
rect 334617 369882 334683 369885
rect 288084 369880 334683 369882
rect 288084 369824 334622 369880
rect 334678 369824 334683 369880
rect 279969 369819 280035 369822
rect 286179 369819 286245 369822
rect 288014 369820 288020 369822
rect 288084 369822 334683 369824
rect 288084 369820 288090 369822
rect 288019 369819 288085 369820
rect 334617 369819 334683 369822
rect 302877 369746 302943 369749
rect 303475 369746 303541 369749
rect 302877 369744 303541 369746
rect 302877 369688 302882 369744
rect 302938 369688 303480 369744
rect 303536 369688 303541 369744
rect 302877 369686 303541 369688
rect 302877 369683 302943 369686
rect 303475 369683 303541 369686
rect 308070 369684 308076 369748
rect 308140 369746 308146 369748
rect 308397 369746 308463 369749
rect 309363 369748 309429 369749
rect 309358 369746 309364 369748
rect 308140 369744 308463 369746
rect 308140 369688 308402 369744
rect 308458 369688 308463 369744
rect 308140 369686 308463 369688
rect 309272 369686 309364 369746
rect 308140 369684 308146 369686
rect 308397 369683 308463 369686
rect 309358 369684 309364 369686
rect 309428 369684 309434 369748
rect 311566 369684 311572 369748
rect 311636 369746 311642 369748
rect 311709 369746 311775 369749
rect 311636 369744 311775 369746
rect 311636 369688 311714 369744
rect 311770 369688 311775 369744
rect 311636 369686 311775 369688
rect 311636 369684 311642 369686
rect 309363 369683 309429 369684
rect 311709 369683 311775 369686
rect 283782 369548 283788 369612
rect 283852 369610 283858 369612
rect 285213 369610 285279 369613
rect 312813 369610 312879 369613
rect 313273 369610 313339 369613
rect 314515 369610 314581 369613
rect 283852 369608 285279 369610
rect 283852 369552 285218 369608
rect 285274 369552 285279 369608
rect 283852 369550 285279 369552
rect 283852 369548 283858 369550
rect 285213 369547 285279 369550
rect 311942 369608 312879 369610
rect 311942 369552 312818 369608
rect 312874 369552 312879 369608
rect 311942 369550 312879 369552
rect 283046 369412 283052 369476
rect 283116 369474 283122 369476
rect 283649 369474 283715 369477
rect 283116 369472 283715 369474
rect 283116 369416 283654 369472
rect 283710 369416 283715 369472
rect 283116 369414 283715 369416
rect 283116 369412 283122 369414
rect 283649 369411 283715 369414
rect 283966 369412 283972 369476
rect 284036 369474 284042 369476
rect 284477 369474 284543 369477
rect 284937 369476 285003 369477
rect 284036 369472 284543 369474
rect 284036 369416 284482 369472
rect 284538 369416 284543 369472
rect 284036 369414 284543 369416
rect 284036 369412 284042 369414
rect 284477 369411 284543 369414
rect 284886 369412 284892 369476
rect 284956 369474 285003 369476
rect 284956 369472 285048 369474
rect 284998 369416 285048 369472
rect 284956 369414 285048 369416
rect 284956 369412 285003 369414
rect 287278 369412 287284 369476
rect 287348 369474 287354 369476
rect 287421 369474 287487 369477
rect 299289 369474 299355 369477
rect 287348 369472 287487 369474
rect 287348 369416 287426 369472
rect 287482 369416 287487 369472
rect 287348 369414 287487 369416
rect 287348 369412 287354 369414
rect 284937 369411 285003 369412
rect 287421 369411 287487 369414
rect 292530 369472 299355 369474
rect 292530 369416 299294 369472
rect 299350 369416 299355 369472
rect 292530 369414 299355 369416
rect 286547 369338 286613 369341
rect 282870 369336 286613 369338
rect 282870 369280 286552 369336
rect 286608 369280 286613 369336
rect 282870 369278 286613 369280
rect 282678 369140 282684 369204
rect 282748 369202 282754 369204
rect 282870 369202 282930 369278
rect 286547 369275 286613 369278
rect 282748 369142 282930 369202
rect 282748 369140 282754 369142
rect 253933 369066 253999 369069
rect 292530 369066 292590 369414
rect 299289 369411 299355 369414
rect 299974 369412 299980 369476
rect 300044 369474 300050 369476
rect 301773 369474 301839 369477
rect 300044 369472 301839 369474
rect 300044 369416 301778 369472
rect 301834 369416 301839 369472
rect 300044 369414 301839 369416
rect 300044 369412 300050 369414
rect 301773 369411 301839 369414
rect 302734 369412 302740 369476
rect 302804 369474 302810 369476
rect 302877 369474 302943 369477
rect 302804 369472 302943 369474
rect 302804 369416 302882 369472
rect 302938 369416 302943 369472
rect 302804 369414 302943 369416
rect 302804 369412 302810 369414
rect 302877 369411 302943 369414
rect 303654 369412 303660 369476
rect 303724 369474 303730 369476
rect 303981 369474 304047 369477
rect 305453 369476 305519 369477
rect 305453 369474 305500 369476
rect 303724 369472 304047 369474
rect 303724 369416 303986 369472
rect 304042 369416 304047 369472
rect 303724 369414 304047 369416
rect 305408 369472 305500 369474
rect 305408 369416 305458 369472
rect 305408 369414 305500 369416
rect 303724 369412 303730 369414
rect 303981 369411 304047 369414
rect 305453 369412 305500 369414
rect 305564 369412 305570 369476
rect 306414 369412 306420 369476
rect 306484 369474 306490 369476
rect 307293 369474 307359 369477
rect 309869 369476 309935 369477
rect 309869 369474 309916 369476
rect 306484 369472 307359 369474
rect 306484 369416 307298 369472
rect 307354 369416 307359 369472
rect 306484 369414 307359 369416
rect 309824 369472 309916 369474
rect 309824 369416 309874 369472
rect 309824 369414 309916 369416
rect 306484 369412 306490 369414
rect 305453 369411 305519 369412
rect 307293 369411 307359 369414
rect 309869 369412 309916 369414
rect 309980 369412 309986 369476
rect 310099 369472 310165 369477
rect 310973 369476 311039 369477
rect 310973 369474 311020 369476
rect 310099 369416 310104 369472
rect 310160 369416 310165 369472
rect 309869 369411 309935 369412
rect 310099 369411 310165 369416
rect 310928 369472 311020 369474
rect 310928 369416 310978 369472
rect 310928 369414 311020 369416
rect 310973 369412 311020 369414
rect 311084 369412 311090 369476
rect 311750 369412 311756 369476
rect 311820 369474 311826 369476
rect 311942 369474 312002 369550
rect 312813 369547 312879 369550
rect 313046 369608 314581 369610
rect 313046 369552 313278 369608
rect 313334 369552 314520 369608
rect 314576 369552 314581 369608
rect 313046 369550 314581 369552
rect 311820 369414 312002 369474
rect 312077 369474 312143 369477
rect 312077 369472 312370 369474
rect 312077 369416 312082 369472
rect 312138 369416 312370 369472
rect 312077 369414 312370 369416
rect 311820 369412 311826 369414
rect 310973 369411 311039 369412
rect 312077 369411 312143 369414
rect 310102 369341 310162 369411
rect 312310 369341 312370 369414
rect 307518 369276 307524 369340
rect 307588 369338 307594 369340
rect 308995 369338 309061 369341
rect 310099 369340 310165 369341
rect 310094 369338 310100 369340
rect 307588 369336 309061 369338
rect 307588 369280 309000 369336
rect 309056 369280 309061 369336
rect 307588 369278 309061 369280
rect 310008 369278 310100 369338
rect 307588 369276 307594 369278
rect 308995 369275 309061 369278
rect 310094 369276 310100 369278
rect 310164 369276 310170 369340
rect 312307 369336 312373 369341
rect 312307 369280 312312 369336
rect 312368 369280 312373 369336
rect 310099 369275 310165 369276
rect 312307 369275 312373 369280
rect 253933 369064 292590 369066
rect 253933 369008 253938 369064
rect 253994 369008 292590 369064
rect 253933 369006 292590 369008
rect 253933 369003 253999 369006
rect 251265 368930 251331 368933
rect 312310 368930 312370 369275
rect 251265 368928 312370 368930
rect 251265 368872 251270 368928
rect 251326 368872 312370 368928
rect 251265 368870 312370 368872
rect 251265 368867 251331 368870
rect 254117 368794 254183 368797
rect 313046 368794 313106 369550
rect 313273 369547 313339 369550
rect 314515 369547 314581 369550
rect 313222 369412 313228 369476
rect 313292 369474 313298 369476
rect 313917 369474 313983 369477
rect 313292 369472 313983 369474
rect 313292 369416 313922 369472
rect 313978 369416 313983 369472
rect 313292 369414 313983 369416
rect 313292 369412 313298 369414
rect 313917 369411 313983 369414
rect 314694 369412 314700 369476
rect 314764 369474 314770 369476
rect 315021 369474 315087 369477
rect 314764 369472 315087 369474
rect 314764 369416 315026 369472
rect 315082 369416 315087 369472
rect 314764 369414 315087 369416
rect 314764 369412 314770 369414
rect 315021 369411 315087 369414
rect 320214 369412 320220 369476
rect 320284 369474 320290 369476
rect 320909 369474 320975 369477
rect 320284 369472 320975 369474
rect 320284 369416 320914 369472
rect 320970 369416 320975 369472
rect 320284 369414 320975 369416
rect 320284 369412 320290 369414
rect 320909 369411 320975 369414
rect 322790 369412 322796 369476
rect 322860 369474 322866 369476
rect 324221 369474 324287 369477
rect 322860 369472 324287 369474
rect 322860 369416 324226 369472
rect 324282 369416 324287 369472
rect 322860 369414 324287 369416
rect 322860 369412 322866 369414
rect 324221 369411 324287 369414
rect 313411 369340 313477 369341
rect 316723 369340 316789 369341
rect 313406 369338 313412 369340
rect 313320 369278 313412 369338
rect 313406 369276 313412 369278
rect 313476 369276 313482 369340
rect 316718 369338 316724 369340
rect 316632 369278 316724 369338
rect 316718 369276 316724 369278
rect 316788 369276 316794 369340
rect 313411 369275 313477 369276
rect 316723 369275 316789 369276
rect 254117 368792 313106 368794
rect 254117 368736 254122 368792
rect 254178 368736 313106 368792
rect 254117 368734 313106 368736
rect 254117 368731 254183 368734
rect 249885 368658 249951 368661
rect 310094 368658 310100 368660
rect 249885 368656 310100 368658
rect 249885 368600 249890 368656
rect 249946 368600 310100 368656
rect 249885 368598 310100 368600
rect 249885 368595 249951 368598
rect 310094 368596 310100 368598
rect 310164 368596 310170 368660
rect 251357 367842 251423 367845
rect 285622 367842 285628 367844
rect 251357 367840 285628 367842
rect 251357 367784 251362 367840
rect 251418 367784 285628 367840
rect 251357 367782 285628 367784
rect 251357 367779 251423 367782
rect 285622 367780 285628 367782
rect 285692 367780 285698 367844
rect 227713 367706 227779 367709
rect 288014 367706 288020 367708
rect 227713 367704 288020 367706
rect 227713 367648 227718 367704
rect 227774 367648 288020 367704
rect 227713 367646 288020 367648
rect 227713 367643 227779 367646
rect 288014 367644 288020 367646
rect 288084 367644 288090 367708
rect 226977 367570 227043 367573
rect 284886 367570 284892 367572
rect 226977 367568 284892 367570
rect 226977 367512 226982 367568
rect 227038 367512 284892 367568
rect 226977 367510 284892 367512
rect 226977 367507 227043 367510
rect 284886 367508 284892 367510
rect 284956 367508 284962 367572
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 224217 363626 224283 363629
rect 282361 363626 282427 363629
rect 224217 363624 282427 363626
rect 224217 363568 224222 363624
rect 224278 363568 282366 363624
rect 282422 363568 282427 363624
rect 224217 363566 282427 363568
rect 224217 363563 224283 363566
rect 282361 363563 282427 363566
rect 225597 362266 225663 362269
rect 283782 362266 283788 362268
rect 225597 362264 283788 362266
rect 225597 362208 225602 362264
rect 225658 362208 283788 362264
rect 225597 362206 283788 362208
rect 225597 362203 225663 362206
rect 283782 362204 283788 362206
rect 283852 362204 283858 362268
rect 280705 360226 280771 360229
rect 281390 360226 281396 360228
rect 280705 360224 281396 360226
rect 280705 360168 280710 360224
rect 280766 360168 281396 360224
rect 280705 360166 281396 360168
rect 280705 360163 280771 360166
rect 281390 360164 281396 360166
rect 281460 360226 281466 360228
rect 283966 360226 283972 360228
rect 281460 360166 283972 360226
rect 281460 360164 281466 360166
rect 283966 360164 283972 360166
rect 284036 360164 284042 360228
rect 280705 358866 280771 358869
rect 281257 358866 281323 358869
rect 280705 358864 281323 358866
rect 280705 358808 280710 358864
rect 280766 358808 281262 358864
rect 281318 358808 281323 358864
rect 280705 358806 281323 358808
rect 280705 358803 280771 358806
rect 281257 358803 281323 358806
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 583520 351780 584960 351870
rect 256785 345674 256851 345677
rect 282269 345674 282335 345677
rect 256785 345672 282335 345674
rect 256785 345616 256790 345672
rect 256846 345616 282274 345672
rect 282330 345616 282335 345672
rect 256785 345614 282335 345616
rect 256785 345611 256851 345614
rect 282269 345611 282335 345614
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 225229 329082 225295 329085
rect 282177 329082 282243 329085
rect 225229 329080 282243 329082
rect 225229 329024 225234 329080
rect 225290 329024 282182 329080
rect 282238 329024 282243 329080
rect 225229 329022 282243 329024
rect 225229 329019 225295 329022
rect 282177 329019 282243 329022
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 220721 322146 220787 322149
rect 282269 322146 282335 322149
rect 220721 322144 282335 322146
rect 220721 322088 220726 322144
rect 220782 322088 282274 322144
rect 282330 322088 282335 322144
rect 220721 322086 282335 322088
rect 220721 322083 220787 322086
rect 282269 322083 282335 322086
rect 217961 322010 218027 322013
rect 281993 322010 282059 322013
rect 217961 322008 282059 322010
rect 217961 321952 217966 322008
rect 218022 321952 281998 322008
rect 282054 321952 282059 322008
rect 217961 321950 282059 321952
rect 217961 321947 218027 321950
rect 281993 321947 282059 321950
rect 213729 321874 213795 321877
rect 283966 321874 283972 321876
rect 213729 321872 283972 321874
rect 213729 321816 213734 321872
rect 213790 321816 283972 321872
rect 213729 321814 283972 321816
rect 213729 321811 213795 321814
rect 283966 321812 283972 321814
rect 284036 321812 284042 321876
rect 220629 321738 220695 321741
rect 293166 321738 293172 321740
rect 220629 321736 293172 321738
rect 220629 321680 220634 321736
rect 220690 321680 293172 321736
rect 220629 321678 293172 321680
rect 220629 321675 220695 321678
rect 293166 321676 293172 321678
rect 293236 321676 293242 321740
rect 213637 321602 213703 321605
rect 288014 321602 288020 321604
rect 213637 321600 288020 321602
rect 213637 321544 213642 321600
rect 213698 321544 288020 321600
rect 213637 321542 288020 321544
rect 213637 321539 213703 321542
rect 288014 321540 288020 321542
rect 288084 321540 288090 321604
rect 319294 321540 319300 321604
rect 319364 321602 319370 321604
rect 335353 321602 335419 321605
rect 319364 321600 335419 321602
rect 319364 321544 335358 321600
rect 335414 321544 335419 321600
rect 319364 321542 335419 321544
rect 319364 321540 319370 321542
rect 335353 321539 335419 321542
rect 247125 321330 247191 321333
rect 306414 321330 306420 321332
rect 247125 321328 306420 321330
rect 247125 321272 247130 321328
rect 247186 321272 306420 321328
rect 247125 321270 306420 321272
rect 247125 321267 247191 321270
rect 306414 321268 306420 321270
rect 306484 321268 306490 321332
rect 317454 321268 317460 321332
rect 317524 321330 317530 321332
rect 327717 321330 327783 321333
rect 317524 321328 327783 321330
rect 317524 321272 327722 321328
rect 327778 321272 327783 321328
rect 317524 321270 327783 321272
rect 317524 321268 317530 321270
rect 327717 321267 327783 321270
rect 248413 321194 248479 321197
rect 307702 321194 307708 321196
rect 248413 321192 307708 321194
rect 248413 321136 248418 321192
rect 248474 321136 307708 321192
rect 248413 321134 307708 321136
rect 248413 321131 248479 321134
rect 307702 321132 307708 321134
rect 307772 321132 307778 321196
rect 310646 321132 310652 321196
rect 310716 321194 310722 321196
rect 314694 321194 314700 321196
rect 310716 321134 314700 321194
rect 310716 321132 310722 321134
rect 314694 321132 314700 321134
rect 314764 321132 314770 321196
rect 335445 321194 335511 321197
rect 323350 321192 335511 321194
rect 323350 321136 335450 321192
rect 335506 321136 335511 321192
rect 323350 321134 335511 321136
rect 242985 321058 243051 321061
rect 303654 321058 303660 321060
rect 242985 321056 303660 321058
rect 242985 321000 242990 321056
rect 243046 321000 303660 321056
rect 242985 320998 303660 321000
rect 242985 320995 243051 320998
rect 303654 320996 303660 320998
rect 303724 320996 303730 321060
rect 252645 320922 252711 320925
rect 313406 320922 313412 320924
rect 252645 320920 313412 320922
rect 252645 320864 252650 320920
rect 252706 320864 313412 320920
rect 252645 320862 313412 320864
rect 252645 320859 252711 320862
rect 313406 320860 313412 320862
rect 313476 320860 313482 320924
rect 323350 320789 323410 321134
rect 335445 321131 335511 321134
rect 332777 321058 332843 321061
rect 324454 321056 332843 321058
rect 324454 321000 332782 321056
rect 332838 321000 332843 321056
rect 324454 320998 332843 321000
rect 324454 320789 324514 320998
rect 332777 320995 332843 320998
rect 325366 320860 325372 320924
rect 325436 320922 325442 320924
rect 327533 320922 327599 320925
rect 325436 320920 327599 320922
rect 325436 320864 327538 320920
rect 327594 320864 327599 320920
rect 325436 320862 327599 320864
rect 325436 320860 325442 320862
rect 327533 320859 327599 320862
rect 226425 320786 226491 320789
rect 288019 320788 288085 320789
rect 287278 320786 287284 320788
rect 226425 320784 287284 320786
rect 226425 320728 226430 320784
rect 226486 320728 287284 320784
rect 226425 320726 287284 320728
rect 226425 320723 226491 320726
rect 287278 320724 287284 320726
rect 287348 320724 287354 320788
rect 288014 320786 288020 320788
rect 287928 320726 288020 320786
rect 288014 320724 288020 320726
rect 288084 320724 288090 320788
rect 290135 320786 290201 320789
rect 291878 320786 291884 320788
rect 290135 320784 291884 320786
rect 290135 320728 290140 320784
rect 290196 320728 291884 320784
rect 290135 320726 291884 320728
rect 288019 320723 288085 320724
rect 290135 320723 290201 320726
rect 291878 320724 291884 320726
rect 291948 320724 291954 320788
rect 292614 320724 292620 320788
rect 292684 320786 292690 320788
rect 293447 320786 293513 320789
rect 292684 320784 293513 320786
rect 292684 320728 293452 320784
rect 293508 320728 293513 320784
rect 292684 320726 293513 320728
rect 292684 320724 292690 320726
rect 293447 320723 293513 320726
rect 294091 320786 294157 320789
rect 294454 320786 294460 320788
rect 294091 320784 294460 320786
rect 294091 320728 294096 320784
rect 294152 320728 294460 320784
rect 294091 320726 294460 320728
rect 294091 320723 294157 320726
rect 294454 320724 294460 320726
rect 294524 320724 294530 320788
rect 295379 320786 295445 320789
rect 295742 320786 295748 320788
rect 295379 320784 295748 320786
rect 295379 320728 295384 320784
rect 295440 320728 295748 320784
rect 295379 320726 295748 320728
rect 295379 320723 295445 320726
rect 295742 320724 295748 320726
rect 295812 320724 295818 320788
rect 299238 320724 299244 320788
rect 299308 320786 299314 320788
rect 299427 320786 299493 320789
rect 299308 320784 299493 320786
rect 299308 320728 299432 320784
rect 299488 320728 299493 320784
rect 299308 320726 299493 320728
rect 299308 320724 299314 320726
rect 299427 320723 299493 320726
rect 311203 320786 311269 320789
rect 322238 320786 322244 320788
rect 311203 320784 322244 320786
rect 311203 320728 311208 320784
rect 311264 320728 322244 320784
rect 311203 320726 322244 320728
rect 311203 320723 311269 320726
rect 322238 320724 322244 320726
rect 322308 320724 322314 320788
rect 323347 320784 323413 320789
rect 323347 320728 323352 320784
rect 323408 320728 323413 320784
rect 323347 320723 323413 320728
rect 324451 320784 324517 320789
rect 328545 320786 328611 320789
rect 324451 320728 324456 320784
rect 324512 320728 324517 320784
rect 324451 320723 324517 320728
rect 324822 320784 328611 320786
rect 324822 320728 328550 320784
rect 328606 320728 328611 320784
rect 324822 320726 328611 320728
rect 241605 320650 241671 320653
rect 299974 320650 299980 320652
rect 241605 320648 299980 320650
rect 241605 320592 241610 320648
rect 241666 320592 299980 320648
rect 241605 320590 299980 320592
rect 241605 320587 241671 320590
rect 299974 320588 299980 320590
rect 300044 320588 300050 320652
rect 311939 320650 312005 320653
rect 312854 320650 312860 320652
rect 311939 320648 312860 320650
rect 311939 320592 311944 320648
rect 312000 320592 312860 320648
rect 311939 320590 312860 320592
rect 311939 320587 312005 320590
rect 312854 320588 312860 320590
rect 312924 320588 312930 320652
rect 313135 320650 313201 320653
rect 313406 320650 313412 320652
rect 313135 320648 313412 320650
rect 313135 320592 313140 320648
rect 313196 320592 313412 320648
rect 313135 320590 313412 320592
rect 313135 320587 313201 320590
rect 313406 320588 313412 320590
rect 313476 320588 313482 320652
rect 322795 320650 322861 320653
rect 324822 320650 324882 320726
rect 328545 320723 328611 320726
rect 322795 320648 324882 320650
rect 322795 320592 322800 320648
rect 322856 320592 324882 320648
rect 322795 320590 324882 320592
rect 325003 320650 325069 320653
rect 334433 320650 334499 320653
rect 325003 320648 334499 320650
rect 325003 320592 325008 320648
rect 325064 320592 334438 320648
rect 334494 320592 334499 320648
rect 325003 320590 334499 320592
rect 322795 320587 322861 320590
rect 325003 320587 325069 320590
rect 334433 320587 334499 320590
rect 254025 320514 254091 320517
rect 313222 320514 313228 320516
rect 254025 320512 313228 320514
rect 254025 320456 254030 320512
rect 254086 320456 313228 320512
rect 254025 320454 313228 320456
rect 254025 320451 254091 320454
rect 313222 320452 313228 320454
rect 313292 320452 313298 320516
rect 315067 320514 315133 320517
rect 317454 320514 317460 320516
rect 315067 320512 317460 320514
rect 315067 320456 315072 320512
rect 315128 320456 317460 320512
rect 315067 320454 317460 320456
rect 315067 320451 315133 320454
rect 317454 320452 317460 320454
rect 317524 320452 317530 320516
rect 317643 320514 317709 320517
rect 318558 320514 318564 320516
rect 317643 320512 318564 320514
rect 317643 320456 317648 320512
rect 317704 320456 318564 320512
rect 317643 320454 318564 320456
rect 317643 320451 317709 320454
rect 318558 320452 318564 320454
rect 318628 320452 318634 320516
rect 318839 320514 318905 320517
rect 319110 320514 319116 320516
rect 318839 320512 319116 320514
rect 318839 320456 318844 320512
rect 318900 320456 319116 320512
rect 318839 320454 319116 320456
rect 318839 320451 318905 320454
rect 319110 320452 319116 320454
rect 319180 320452 319186 320516
rect 323899 320514 323965 320517
rect 325366 320514 325372 320516
rect 323899 320512 325372 320514
rect 323899 320456 323904 320512
rect 323960 320456 325372 320512
rect 323899 320454 325372 320456
rect 323899 320451 323965 320454
rect 325366 320452 325372 320454
rect 325436 320452 325442 320516
rect 325555 320514 325621 320517
rect 330201 320514 330267 320517
rect 325555 320512 330267 320514
rect 325555 320456 325560 320512
rect 325616 320456 330206 320512
rect 330262 320456 330267 320512
rect 325555 320454 330267 320456
rect 325555 320451 325621 320454
rect 330201 320451 330267 320454
rect 280153 320378 280219 320381
rect 282959 320378 283025 320381
rect 280153 320376 283025 320378
rect 280153 320320 280158 320376
rect 280214 320320 282964 320376
rect 283020 320320 283025 320376
rect 280153 320318 283025 320320
rect 280153 320315 280219 320318
rect 282959 320315 283025 320318
rect 283235 320378 283301 320381
rect 283787 320380 283853 320381
rect 283414 320378 283420 320380
rect 283235 320376 283420 320378
rect 283235 320320 283240 320376
rect 283296 320320 283420 320376
rect 283235 320318 283420 320320
rect 283235 320315 283301 320318
rect 283414 320316 283420 320318
rect 283484 320316 283490 320380
rect 283782 320378 283788 320380
rect 283696 320318 283788 320378
rect 283782 320316 283788 320318
rect 283852 320316 283858 320380
rect 288934 320316 288940 320380
rect 289004 320378 289010 320380
rect 289675 320378 289741 320381
rect 289004 320376 289741 320378
rect 289004 320320 289680 320376
rect 289736 320320 289741 320376
rect 289004 320318 289741 320320
rect 289004 320316 289010 320318
rect 283787 320315 283853 320316
rect 289675 320315 289741 320318
rect 290774 320316 290780 320380
rect 290844 320378 290850 320380
rect 291055 320378 291121 320381
rect 290844 320376 291121 320378
rect 290844 320320 291060 320376
rect 291116 320320 291121 320376
rect 290844 320318 291121 320320
rect 290844 320316 290850 320318
rect 291055 320315 291121 320318
rect 292798 320316 292804 320380
rect 292868 320378 292874 320380
rect 297679 320378 297745 320381
rect 292868 320376 297745 320378
rect 292868 320320 297684 320376
rect 297740 320320 297745 320376
rect 292868 320318 297745 320320
rect 292868 320316 292874 320318
rect 297679 320315 297745 320318
rect 298047 320378 298113 320381
rect 298599 320378 298665 320381
rect 299606 320378 299612 320380
rect 298047 320376 298156 320378
rect 298047 320320 298052 320376
rect 298108 320320 298156 320376
rect 298047 320315 298156 320320
rect 298599 320376 299612 320378
rect 298599 320320 298604 320376
rect 298660 320320 299612 320376
rect 298599 320318 299612 320320
rect 298599 320315 298665 320318
rect 299606 320316 299612 320318
rect 299676 320316 299682 320380
rect 299790 320316 299796 320380
rect 299860 320378 299866 320380
rect 300623 320378 300689 320381
rect 299860 320376 300689 320378
rect 299860 320320 300628 320376
rect 300684 320320 300689 320376
rect 299860 320318 300689 320320
rect 299860 320316 299866 320318
rect 300623 320315 300689 320318
rect 307702 320316 307708 320380
rect 307772 320378 307778 320380
rect 308903 320378 308969 320381
rect 312215 320378 312281 320381
rect 313227 320380 313293 320381
rect 317091 320380 317157 320381
rect 318747 320380 318813 320381
rect 313222 320378 313228 320380
rect 307772 320376 308969 320378
rect 307772 320320 308908 320376
rect 308964 320320 308969 320376
rect 307772 320318 308969 320320
rect 307772 320316 307778 320318
rect 308903 320315 308969 320318
rect 311942 320376 312281 320378
rect 311942 320320 312220 320376
rect 312276 320320 312281 320376
rect 311942 320318 312281 320320
rect 313136 320318 313228 320378
rect 281901 320242 281967 320245
rect 285167 320242 285233 320245
rect 281901 320240 285233 320242
rect 281901 320184 281906 320240
rect 281962 320184 285172 320240
rect 285228 320184 285233 320240
rect 281901 320182 285233 320184
rect 281901 320179 281967 320182
rect 285167 320179 285233 320182
rect 285622 320180 285628 320244
rect 285692 320242 285698 320244
rect 286455 320242 286521 320245
rect 286639 320242 286705 320245
rect 285692 320240 286521 320242
rect 285692 320184 286460 320240
rect 286516 320184 286521 320240
rect 285692 320182 286521 320184
rect 285692 320180 285698 320182
rect 286455 320179 286521 320182
rect 286596 320240 286705 320242
rect 286596 320184 286644 320240
rect 286700 320184 286705 320240
rect 286596 320179 286705 320184
rect 287375 320242 287441 320245
rect 287830 320242 287836 320244
rect 287375 320240 287836 320242
rect 287375 320184 287380 320240
rect 287436 320184 287836 320240
rect 287375 320182 287836 320184
rect 287375 320179 287441 320182
rect 287830 320180 287836 320182
rect 287900 320180 287906 320244
rect 288111 320242 288177 320245
rect 288068 320240 288177 320242
rect 288068 320184 288116 320240
rect 288172 320184 288177 320240
rect 288068 320179 288177 320184
rect 288750 320180 288756 320244
rect 288820 320242 288826 320244
rect 289031 320242 289097 320245
rect 288820 320240 289097 320242
rect 288820 320184 289036 320240
rect 289092 320184 289097 320240
rect 288820 320182 289097 320184
rect 288820 320180 288826 320182
rect 289031 320179 289097 320182
rect 289486 320180 289492 320244
rect 289556 320242 289562 320244
rect 290319 320242 290385 320245
rect 290963 320244 291029 320245
rect 291331 320244 291397 320245
rect 290958 320242 290964 320244
rect 289556 320240 290385 320242
rect 289556 320184 290324 320240
rect 290380 320184 290385 320240
rect 289556 320182 290385 320184
rect 290872 320182 290964 320242
rect 289556 320180 289562 320182
rect 290319 320179 290385 320182
rect 290958 320180 290964 320182
rect 291028 320180 291034 320244
rect 291326 320242 291332 320244
rect 291240 320182 291332 320242
rect 291326 320180 291332 320182
rect 291396 320180 291402 320244
rect 293350 320180 293356 320244
rect 293420 320242 293426 320244
rect 293539 320242 293605 320245
rect 293420 320240 293605 320242
rect 293420 320184 293544 320240
rect 293600 320184 293605 320240
rect 293420 320182 293605 320184
rect 293420 320180 293426 320182
rect 290963 320179 291029 320180
rect 291331 320179 291397 320180
rect 293539 320179 293605 320182
rect 294183 320242 294249 320245
rect 294638 320242 294644 320244
rect 294183 320240 294644 320242
rect 294183 320184 294188 320240
rect 294244 320184 294644 320240
rect 294183 320182 294644 320184
rect 294183 320179 294249 320182
rect 294638 320180 294644 320182
rect 294708 320180 294714 320244
rect 294822 320180 294828 320244
rect 294892 320242 294898 320244
rect 296851 320242 296917 320245
rect 294892 320240 296917 320242
rect 294892 320184 296856 320240
rect 296912 320184 296917 320240
rect 294892 320182 296917 320184
rect 294892 320180 294898 320182
rect 296851 320179 296917 320182
rect 297771 320242 297837 320245
rect 297950 320242 297956 320244
rect 297771 320240 297956 320242
rect 297771 320184 297776 320240
rect 297832 320184 297956 320240
rect 297771 320182 297956 320184
rect 297771 320179 297837 320182
rect 297950 320180 297956 320182
rect 298020 320180 298026 320244
rect 282269 320106 282335 320109
rect 282867 320106 282933 320109
rect 282269 320104 282933 320106
rect 282269 320048 282274 320104
rect 282330 320048 282872 320104
rect 282928 320048 282933 320104
rect 282269 320046 282933 320048
rect 282269 320043 282335 320046
rect 282867 320043 282933 320046
rect 283051 320104 283117 320109
rect 283051 320048 283056 320104
rect 283112 320048 283117 320104
rect 283051 320043 283117 320048
rect 283230 320044 283236 320108
rect 283300 320106 283306 320108
rect 284155 320106 284221 320109
rect 283300 320104 284221 320106
rect 283300 320048 284160 320104
rect 284216 320048 284221 320104
rect 283300 320046 284221 320048
rect 283300 320044 283306 320046
rect 284155 320043 284221 320046
rect 284334 320044 284340 320108
rect 284404 320106 284410 320108
rect 284707 320106 284773 320109
rect 285535 320106 285601 320109
rect 284404 320104 284773 320106
rect 284404 320048 284712 320104
rect 284768 320048 284773 320104
rect 284404 320046 284773 320048
rect 284404 320044 284410 320046
rect 284707 320043 284773 320046
rect 285400 320104 285601 320106
rect 285400 320048 285540 320104
rect 285596 320048 285601 320104
rect 285400 320046 285601 320048
rect 283054 319970 283114 320043
rect 285400 319972 285460 320046
rect 285535 320043 285601 320046
rect 285806 320044 285812 320108
rect 285876 320106 285882 320108
rect 286087 320106 286153 320109
rect 285876 320104 286153 320106
rect 285876 320048 286092 320104
rect 286148 320048 286153 320104
rect 285876 320046 286153 320048
rect 286596 320106 286656 320179
rect 287651 320108 287717 320109
rect 288068 320108 288128 320179
rect 286726 320106 286732 320108
rect 286596 320046 286732 320106
rect 285876 320044 285882 320046
rect 286087 320043 286153 320046
rect 286726 320044 286732 320046
rect 286796 320044 286802 320108
rect 287646 320106 287652 320108
rect 287560 320046 287652 320106
rect 287646 320044 287652 320046
rect 287716 320044 287722 320108
rect 288014 320044 288020 320108
rect 288084 320046 288128 320108
rect 288084 320044 288090 320046
rect 288198 320044 288204 320108
rect 288268 320106 288274 320108
rect 288387 320106 288453 320109
rect 288268 320104 288453 320106
rect 288268 320048 288392 320104
rect 288448 320048 288453 320104
rect 288268 320046 288453 320048
rect 288268 320044 288274 320046
rect 287651 320043 287717 320044
rect 288387 320043 288453 320046
rect 288566 320044 288572 320108
rect 288636 320106 288642 320108
rect 288847 320106 288913 320109
rect 288636 320104 288913 320106
rect 288636 320048 288852 320104
rect 288908 320048 288913 320104
rect 288636 320046 288913 320048
rect 288636 320044 288642 320046
rect 288847 320043 288913 320046
rect 289118 320044 289124 320108
rect 289188 320106 289194 320108
rect 289399 320106 289465 320109
rect 289188 320104 289465 320106
rect 289188 320048 289404 320104
rect 289460 320048 289465 320104
rect 289188 320046 289465 320048
rect 289188 320044 289194 320046
rect 289399 320043 289465 320046
rect 289859 320104 289925 320109
rect 289859 320048 289864 320104
rect 289920 320048 289925 320104
rect 289859 320043 289925 320048
rect 290411 320104 290477 320109
rect 290411 320048 290416 320104
rect 290472 320048 290477 320104
rect 290411 320043 290477 320048
rect 290590 320044 290596 320108
rect 290660 320106 290666 320108
rect 290871 320106 290937 320109
rect 291515 320108 291581 320109
rect 291699 320108 291765 320109
rect 291510 320106 291516 320108
rect 290660 320104 290937 320106
rect 290660 320048 290876 320104
rect 290932 320048 290937 320104
rect 290660 320046 290937 320048
rect 291424 320046 291516 320106
rect 290660 320044 290666 320046
rect 290871 320043 290937 320046
rect 291510 320044 291516 320046
rect 291580 320044 291586 320108
rect 291694 320044 291700 320108
rect 291764 320106 291770 320108
rect 291764 320046 291856 320106
rect 291764 320044 291770 320046
rect 292062 320044 292068 320108
rect 292132 320106 292138 320108
rect 292343 320106 292409 320109
rect 292132 320104 292409 320106
rect 292132 320048 292348 320104
rect 292404 320048 292409 320104
rect 292132 320046 292409 320048
rect 292132 320044 292138 320046
rect 291515 320043 291581 320044
rect 291699 320043 291765 320044
rect 292343 320043 292409 320046
rect 292982 320044 292988 320108
rect 293052 320106 293058 320108
rect 293171 320106 293237 320109
rect 293052 320104 293237 320106
rect 293052 320048 293176 320104
rect 293232 320048 293237 320104
rect 293052 320046 293237 320048
rect 293052 320044 293058 320046
rect 293171 320043 293237 320046
rect 293723 320104 293789 320109
rect 294275 320108 294341 320109
rect 295011 320108 295077 320109
rect 295563 320108 295629 320109
rect 295931 320108 295997 320109
rect 294270 320106 294276 320108
rect 293723 320048 293728 320104
rect 293784 320048 293789 320104
rect 293723 320043 293789 320048
rect 294184 320046 294276 320106
rect 294270 320044 294276 320046
rect 294340 320044 294346 320108
rect 295006 320106 295012 320108
rect 294920 320046 295012 320106
rect 295006 320044 295012 320046
rect 295076 320044 295082 320108
rect 295558 320106 295564 320108
rect 295472 320046 295564 320106
rect 295558 320044 295564 320046
rect 295628 320044 295634 320108
rect 295926 320106 295932 320108
rect 295840 320046 295932 320106
rect 295926 320044 295932 320046
rect 295996 320044 296002 320108
rect 296207 320106 296273 320109
rect 296164 320104 296273 320106
rect 296164 320048 296212 320104
rect 296268 320048 296273 320104
rect 294275 320043 294341 320044
rect 295011 320043 295077 320044
rect 295563 320043 295629 320044
rect 295931 320043 295997 320044
rect 296164 320043 296273 320048
rect 297030 320044 297036 320108
rect 297100 320106 297106 320108
rect 297311 320106 297377 320109
rect 297100 320104 297377 320106
rect 297100 320048 297316 320104
rect 297372 320048 297377 320104
rect 297100 320046 297377 320048
rect 297100 320044 297106 320046
rect 297311 320043 297377 320046
rect 283414 319970 283420 319972
rect 283054 319910 283420 319970
rect 283414 319908 283420 319910
rect 283484 319908 283490 319972
rect 285400 319910 285444 319972
rect 285438 319908 285444 319910
rect 285508 319908 285514 319972
rect 289302 319908 289308 319972
rect 289372 319970 289378 319972
rect 289862 319970 289922 320043
rect 289372 319910 289922 319970
rect 290414 319970 290474 320043
rect 291142 319970 291148 319972
rect 290414 319910 291148 319970
rect 289372 319908 289378 319910
rect 291142 319908 291148 319910
rect 291212 319908 291218 319972
rect 292430 319908 292436 319972
rect 292500 319970 292506 319972
rect 293726 319970 293786 320043
rect 292500 319910 293786 319970
rect 292500 319908 292506 319910
rect 295374 319908 295380 319972
rect 295444 319970 295450 319972
rect 296164 319970 296224 320043
rect 295444 319910 296224 319970
rect 295444 319908 295450 319910
rect 296846 319908 296852 319972
rect 296916 319970 296922 319972
rect 298096 319970 298156 320315
rect 299054 320180 299060 320244
rect 299124 320242 299130 320244
rect 299335 320242 299401 320245
rect 299124 320240 299401 320242
rect 299124 320184 299340 320240
rect 299396 320184 299401 320240
rect 299124 320182 299401 320184
rect 299124 320180 299130 320182
rect 299335 320179 299401 320182
rect 300526 320180 300532 320244
rect 300596 320242 300602 320244
rect 300991 320242 301057 320245
rect 300596 320240 301057 320242
rect 300596 320184 300996 320240
rect 301052 320184 301057 320240
rect 300596 320182 301057 320184
rect 300596 320180 300602 320182
rect 300991 320179 301057 320182
rect 303654 320180 303660 320244
rect 303724 320242 303730 320244
rect 304211 320242 304277 320245
rect 303724 320240 304277 320242
rect 303724 320184 304216 320240
rect 304272 320184 304277 320240
rect 303724 320182 304277 320184
rect 303724 320180 303730 320182
rect 304211 320179 304277 320182
rect 308070 320180 308076 320244
rect 308140 320242 308146 320244
rect 308443 320242 308509 320245
rect 308140 320240 308509 320242
rect 308140 320184 308448 320240
rect 308504 320184 308509 320240
rect 308140 320182 308509 320184
rect 308140 320180 308146 320182
rect 308443 320179 308509 320182
rect 309915 320242 309981 320245
rect 310835 320244 310901 320245
rect 310278 320242 310284 320244
rect 309915 320240 310284 320242
rect 309915 320184 309920 320240
rect 309976 320184 310284 320240
rect 309915 320182 310284 320184
rect 309915 320179 309981 320182
rect 310278 320180 310284 320182
rect 310348 320180 310354 320244
rect 310830 320242 310836 320244
rect 310744 320182 310836 320242
rect 310830 320180 310836 320182
rect 310900 320180 310906 320244
rect 311382 320180 311388 320244
rect 311452 320242 311458 320244
rect 311663 320242 311729 320245
rect 311452 320240 311729 320242
rect 311452 320184 311668 320240
rect 311724 320184 311729 320240
rect 311452 320182 311729 320184
rect 311452 320180 311458 320182
rect 310835 320179 310901 320180
rect 311663 320179 311729 320182
rect 298318 320044 298324 320108
rect 298388 320106 298394 320108
rect 299059 320106 299125 320109
rect 298388 320104 299125 320106
rect 298388 320048 299064 320104
rect 299120 320048 299125 320104
rect 298388 320046 299125 320048
rect 298388 320044 298394 320046
rect 299059 320043 299125 320046
rect 299422 320044 299428 320108
rect 299492 320106 299498 320108
rect 299703 320106 299769 320109
rect 299492 320104 299769 320106
rect 299492 320048 299708 320104
rect 299764 320048 299769 320104
rect 299492 320046 299769 320048
rect 299492 320044 299498 320046
rect 299703 320043 299769 320046
rect 299974 320044 299980 320108
rect 300044 320106 300050 320108
rect 300255 320106 300321 320109
rect 300715 320108 300781 320109
rect 300710 320106 300716 320108
rect 300044 320104 300321 320106
rect 300044 320048 300260 320104
rect 300316 320048 300321 320104
rect 300044 320046 300321 320048
rect 300624 320046 300716 320106
rect 300044 320044 300050 320046
rect 300255 320043 300321 320046
rect 300710 320044 300716 320046
rect 300780 320044 300786 320108
rect 301814 320044 301820 320108
rect 301884 320106 301890 320108
rect 302095 320106 302161 320109
rect 301884 320104 302161 320106
rect 301884 320048 302100 320104
rect 302156 320048 302161 320104
rect 301884 320046 302161 320048
rect 301884 320044 301890 320046
rect 300715 320043 300781 320044
rect 302095 320043 302161 320046
rect 302366 320044 302372 320108
rect 302436 320106 302442 320108
rect 302739 320106 302805 320109
rect 303843 320108 303909 320109
rect 304395 320108 304461 320109
rect 303838 320106 303844 320108
rect 302436 320104 302805 320106
rect 302436 320048 302744 320104
rect 302800 320048 302805 320104
rect 302436 320046 302805 320048
rect 303752 320046 303844 320106
rect 302436 320044 302442 320046
rect 302739 320043 302805 320046
rect 303838 320044 303844 320046
rect 303908 320044 303914 320108
rect 304390 320106 304396 320108
rect 304304 320046 304396 320106
rect 304390 320044 304396 320046
rect 304460 320044 304466 320108
rect 305131 320106 305197 320109
rect 306051 320108 306117 320109
rect 306235 320108 306301 320109
rect 305678 320106 305684 320108
rect 305131 320104 305684 320106
rect 305131 320048 305136 320104
rect 305192 320048 305684 320104
rect 305131 320046 305684 320048
rect 303843 320043 303909 320044
rect 304395 320043 304461 320044
rect 305131 320043 305197 320046
rect 305678 320044 305684 320046
rect 305748 320044 305754 320108
rect 306046 320106 306052 320108
rect 305960 320046 306052 320106
rect 306046 320044 306052 320046
rect 306116 320044 306122 320108
rect 306230 320044 306236 320108
rect 306300 320106 306306 320108
rect 306300 320046 306392 320106
rect 306300 320044 306306 320046
rect 306598 320044 306604 320108
rect 306668 320106 306674 320108
rect 306879 320106 306945 320109
rect 307155 320108 307221 320109
rect 307150 320106 307156 320108
rect 306668 320104 306945 320106
rect 306668 320048 306884 320104
rect 306940 320048 306945 320104
rect 306668 320046 306945 320048
rect 307064 320046 307156 320106
rect 306668 320044 306674 320046
rect 306051 320043 306117 320044
rect 306235 320043 306301 320044
rect 306879 320043 306945 320046
rect 307150 320044 307156 320046
rect 307220 320044 307226 320108
rect 307334 320044 307340 320108
rect 307404 320106 307410 320108
rect 307615 320106 307681 320109
rect 307404 320104 307681 320106
rect 307404 320048 307620 320104
rect 307676 320048 307681 320104
rect 307404 320046 307681 320048
rect 307404 320044 307410 320046
rect 307155 320043 307221 320044
rect 307615 320043 307681 320046
rect 307886 320044 307892 320108
rect 307956 320106 307962 320108
rect 308167 320106 308233 320109
rect 307956 320104 308233 320106
rect 307956 320048 308172 320104
rect 308228 320048 308233 320104
rect 307956 320046 308233 320048
rect 307956 320044 307962 320046
rect 308167 320043 308233 320046
rect 309542 320044 309548 320108
rect 309612 320106 309618 320108
rect 309731 320106 309797 320109
rect 309612 320104 309797 320106
rect 309612 320048 309736 320104
rect 309792 320048 309797 320104
rect 309612 320046 309797 320048
rect 309612 320044 309618 320046
rect 309731 320043 309797 320046
rect 309910 320044 309916 320108
rect 309980 320106 309986 320108
rect 310099 320106 310165 320109
rect 310467 320108 310533 320109
rect 310462 320106 310468 320108
rect 309980 320104 310165 320106
rect 309980 320048 310104 320104
rect 310160 320048 310165 320104
rect 309980 320046 310165 320048
rect 310376 320046 310468 320106
rect 309980 320044 309986 320046
rect 310099 320043 310165 320046
rect 310462 320044 310468 320046
rect 310532 320044 310538 320108
rect 310743 320106 310809 320109
rect 311198 320106 311204 320108
rect 310743 320104 311204 320106
rect 310743 320048 310748 320104
rect 310804 320048 311204 320104
rect 310743 320046 311204 320048
rect 310467 320043 310533 320044
rect 310743 320043 310809 320046
rect 311198 320044 311204 320046
rect 311268 320044 311274 320108
rect 311942 320106 312002 320318
rect 312215 320315 312281 320318
rect 313222 320316 313228 320318
rect 313292 320316 313298 320380
rect 317086 320378 317092 320380
rect 317000 320318 317092 320378
rect 317086 320316 317092 320318
rect 317156 320316 317162 320380
rect 318742 320378 318748 320380
rect 318656 320318 318748 320378
rect 318742 320316 318748 320318
rect 318812 320316 318818 320380
rect 318931 320378 318997 320381
rect 323163 320380 323229 320381
rect 323158 320378 323164 320380
rect 318931 320376 320696 320378
rect 318931 320320 318936 320376
rect 318992 320320 320696 320376
rect 318931 320318 320696 320320
rect 323072 320318 323164 320378
rect 313227 320315 313293 320316
rect 317091 320315 317157 320316
rect 318747 320315 318813 320316
rect 318931 320315 318997 320318
rect 312399 320242 312465 320245
rect 312951 320242 313017 320245
rect 314331 320244 314397 320245
rect 314326 320242 314332 320244
rect 312399 320240 312692 320242
rect 312399 320184 312404 320240
rect 312460 320184 312692 320240
rect 312399 320182 312692 320184
rect 312399 320179 312465 320182
rect 311942 320046 312186 320106
rect 296916 319910 298156 319970
rect 296916 319908 296922 319910
rect 306966 319908 306972 319972
rect 307036 319970 307042 319972
rect 310646 319970 310652 319972
rect 307036 319910 310652 319970
rect 307036 319908 307042 319910
rect 310646 319908 310652 319910
rect 310716 319908 310722 319972
rect 260925 319834 260991 319837
rect 310789 319834 310855 319837
rect 260925 319832 310855 319834
rect 260925 319776 260930 319832
rect 260986 319776 310794 319832
rect 310850 319776 310855 319832
rect 260925 319774 310855 319776
rect 312126 319834 312186 320046
rect 312491 320104 312557 320109
rect 312491 320048 312496 320104
rect 312552 320048 312557 320104
rect 312491 320043 312557 320048
rect 312261 319834 312327 319837
rect 312126 319832 312327 319834
rect 312126 319776 312266 319832
rect 312322 319776 312327 319832
rect 312126 319774 312327 319776
rect 260925 319771 260991 319774
rect 310789 319771 310855 319774
rect 312261 319771 312327 319774
rect 256969 319698 257035 319701
rect 256969 319696 312370 319698
rect 256969 319640 256974 319696
rect 257030 319640 312370 319696
rect 256969 319638 312370 319640
rect 256969 319635 257035 319638
rect 254209 319562 254275 319565
rect 307477 319564 307543 319565
rect 306966 319562 306972 319564
rect 254209 319560 306972 319562
rect 254209 319504 254214 319560
rect 254270 319504 306972 319560
rect 254209 319502 306972 319504
rect 254209 319499 254275 319502
rect 306966 319500 306972 319502
rect 307036 319500 307042 319564
rect 307477 319562 307524 319564
rect 307432 319560 307524 319562
rect 307432 319504 307482 319560
rect 307432 319502 307524 319504
rect 307477 319500 307524 319502
rect 307588 319500 307594 319564
rect 307702 319500 307708 319564
rect 307772 319562 307778 319564
rect 308765 319562 308831 319565
rect 309501 319564 309567 319565
rect 309501 319562 309548 319564
rect 307772 319560 308831 319562
rect 307772 319504 308770 319560
rect 308826 319504 308831 319560
rect 307772 319502 308831 319504
rect 309456 319560 309548 319562
rect 309456 319504 309506 319560
rect 309456 319502 309548 319504
rect 307772 319500 307778 319502
rect 307477 319499 307543 319500
rect 308765 319499 308831 319502
rect 309501 319500 309548 319502
rect 309612 319500 309618 319564
rect 309685 319562 309751 319565
rect 311014 319562 311020 319564
rect 309685 319560 311020 319562
rect 309685 319504 309690 319560
rect 309746 319504 311020 319560
rect 309685 319502 311020 319504
rect 309501 319499 309567 319500
rect 309685 319499 309751 319502
rect 311014 319500 311020 319502
rect 311084 319500 311090 319564
rect 311341 319562 311407 319565
rect 311566 319562 311572 319564
rect 311341 319560 311572 319562
rect 311341 319504 311346 319560
rect 311402 319504 311572 319560
rect 311341 319502 311572 319504
rect 311341 319499 311407 319502
rect 311566 319500 311572 319502
rect 311636 319500 311642 319564
rect 244365 319426 244431 319429
rect 293217 319428 293283 319429
rect 244365 319424 292590 319426
rect -960 319290 480 319380
rect 244365 319368 244370 319424
rect 244426 319368 292590 319424
rect 244365 319366 292590 319368
rect 244365 319363 244431 319366
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 282361 319290 282427 319293
rect 283046 319290 283052 319292
rect 282361 319288 283052 319290
rect 282361 319232 282366 319288
rect 282422 319232 283052 319288
rect 282361 319230 283052 319232
rect 282361 319227 282427 319230
rect 283046 319228 283052 319230
rect 283116 319290 283122 319292
rect 283465 319290 283531 319293
rect 284017 319292 284083 319293
rect 283116 319288 283531 319290
rect 283116 319232 283470 319288
rect 283526 319232 283531 319288
rect 283116 319230 283531 319232
rect 283116 319228 283122 319230
rect 283465 319227 283531 319230
rect 283966 319228 283972 319292
rect 284036 319290 284083 319292
rect 284569 319290 284635 319293
rect 285029 319290 285095 319293
rect 285489 319292 285555 319293
rect 284036 319288 284128 319290
rect 284078 319232 284128 319288
rect 284036 319230 284128 319232
rect 284569 319288 285095 319290
rect 284569 319232 284574 319288
rect 284630 319232 285034 319288
rect 285090 319232 285095 319288
rect 284569 319230 285095 319232
rect 284036 319228 284083 319230
rect 284017 319227 284083 319228
rect 284569 319227 284635 319230
rect 285029 319227 285095 319230
rect 285438 319228 285444 319292
rect 285508 319290 285555 319292
rect 285508 319288 285600 319290
rect 285550 319232 285600 319288
rect 285508 319230 285600 319232
rect 285508 319228 285555 319230
rect 287646 319228 287652 319292
rect 287716 319290 287722 319292
rect 288065 319290 288131 319293
rect 287716 319288 288131 319290
rect 287716 319232 288070 319288
rect 288126 319232 288131 319288
rect 287716 319230 288131 319232
rect 287716 319228 287722 319230
rect 285489 319227 285555 319228
rect 288065 319227 288131 319230
rect 289302 319228 289308 319292
rect 289372 319290 289378 319292
rect 289905 319290 289971 319293
rect 289372 319288 289971 319290
rect 289372 319232 289910 319288
rect 289966 319232 289971 319288
rect 289372 319230 289971 319232
rect 289372 319228 289378 319230
rect 289905 319227 289971 319230
rect 290365 319290 290431 319293
rect 290590 319290 290596 319292
rect 290365 319288 290596 319290
rect 290365 319232 290370 319288
rect 290426 319232 290596 319288
rect 290365 319230 290596 319232
rect 290365 319227 290431 319230
rect 290590 319228 290596 319230
rect 290660 319228 290666 319292
rect 290825 319290 290891 319293
rect 290958 319290 290964 319292
rect 290825 319288 290964 319290
rect 290825 319232 290830 319288
rect 290886 319232 290964 319288
rect 290825 319230 290964 319232
rect 290825 319227 290891 319230
rect 290958 319228 290964 319230
rect 291028 319228 291034 319292
rect 291193 319290 291259 319293
rect 291510 319290 291516 319292
rect 291193 319288 291516 319290
rect 291193 319232 291198 319288
rect 291254 319232 291516 319288
rect 291193 319230 291516 319232
rect 291193 319227 291259 319230
rect 291510 319228 291516 319230
rect 291580 319228 291586 319292
rect 292530 319290 292590 319366
rect 293166 319364 293172 319428
rect 293236 319426 293283 319428
rect 294597 319426 294663 319429
rect 294822 319426 294828 319428
rect 293236 319424 293328 319426
rect 293278 319368 293328 319424
rect 293236 319366 293328 319368
rect 294597 319424 294828 319426
rect 294597 319368 294602 319424
rect 294658 319368 294828 319424
rect 294597 319366 294828 319368
rect 293236 319364 293283 319366
rect 293217 319363 293283 319364
rect 294597 319363 294663 319366
rect 294822 319364 294828 319366
rect 294892 319364 294898 319428
rect 295333 319426 295399 319429
rect 296478 319426 296484 319428
rect 295333 319424 296484 319426
rect 295333 319368 295338 319424
rect 295394 319368 296484 319424
rect 295333 319366 296484 319368
rect 295333 319363 295399 319366
rect 296478 319364 296484 319366
rect 296548 319364 296554 319428
rect 299841 319426 299907 319429
rect 299974 319426 299980 319428
rect 299841 319424 299980 319426
rect 299841 319368 299846 319424
rect 299902 319368 299980 319424
rect 299841 319366 299980 319368
rect 299841 319363 299907 319366
rect 299974 319364 299980 319366
rect 300044 319364 300050 319428
rect 300393 319426 300459 319429
rect 300710 319426 300716 319428
rect 300393 319424 300716 319426
rect 300393 319368 300398 319424
rect 300454 319368 300716 319424
rect 300393 319366 300716 319368
rect 300393 319363 300459 319366
rect 300710 319364 300716 319366
rect 300780 319364 300786 319428
rect 301814 319364 301820 319428
rect 301884 319426 301890 319428
rect 302141 319426 302207 319429
rect 301884 319424 302207 319426
rect 301884 319368 302146 319424
rect 302202 319368 302207 319424
rect 301884 319366 302207 319368
rect 301884 319364 301890 319366
rect 302141 319363 302207 319366
rect 302509 319426 302575 319429
rect 302918 319426 302924 319428
rect 302509 319424 302924 319426
rect 302509 319368 302514 319424
rect 302570 319368 302924 319424
rect 302509 319366 302924 319368
rect 302509 319363 302575 319366
rect 302918 319364 302924 319366
rect 302988 319364 302994 319428
rect 304165 319426 304231 319429
rect 304390 319426 304396 319428
rect 304165 319424 304396 319426
rect 304165 319368 304170 319424
rect 304226 319368 304396 319424
rect 304165 319366 304396 319368
rect 304165 319363 304231 319366
rect 304390 319364 304396 319366
rect 304460 319364 304466 319428
rect 305729 319426 305795 319429
rect 306281 319428 306347 319429
rect 306046 319426 306052 319428
rect 305729 319424 306052 319426
rect 305729 319368 305734 319424
rect 305790 319368 306052 319424
rect 305729 319366 306052 319368
rect 305729 319363 305795 319366
rect 306046 319364 306052 319366
rect 306116 319364 306122 319428
rect 306230 319364 306236 319428
rect 306300 319426 306347 319428
rect 306300 319424 306392 319426
rect 306342 319368 306392 319424
rect 306300 319366 306392 319368
rect 306300 319364 306347 319366
rect 306598 319364 306604 319428
rect 306668 319426 306674 319428
rect 306833 319426 306899 319429
rect 306668 319424 306899 319426
rect 306668 319368 306838 319424
rect 306894 319368 306899 319424
rect 306668 319366 306899 319368
rect 306668 319364 306674 319366
rect 306281 319363 306347 319364
rect 306833 319363 306899 319366
rect 308070 319364 308076 319428
rect 308140 319426 308146 319428
rect 308489 319426 308555 319429
rect 308140 319424 308555 319426
rect 308140 319368 308494 319424
rect 308550 319368 308555 319424
rect 308140 319366 308555 319368
rect 308140 319364 308146 319366
rect 308489 319363 308555 319366
rect 309317 319426 309383 319429
rect 310094 319426 310100 319428
rect 309317 319424 310100 319426
rect 309317 319368 309322 319424
rect 309378 319368 310100 319424
rect 309317 319366 310100 319368
rect 309317 319363 309383 319366
rect 310094 319364 310100 319366
rect 310164 319364 310170 319428
rect 310881 319426 310947 319429
rect 311750 319426 311756 319428
rect 310881 319424 311756 319426
rect 310881 319368 310886 319424
rect 310942 319368 311756 319424
rect 310881 319366 311756 319368
rect 310881 319363 310947 319366
rect 311750 319364 311756 319366
rect 311820 319364 311826 319428
rect 312310 319426 312370 319638
rect 312494 319565 312554 320043
rect 312632 319701 312692 320182
rect 312951 320240 313290 320242
rect 312951 320184 312956 320240
rect 313012 320184 313290 320240
rect 312951 320182 313290 320184
rect 314240 320182 314332 320242
rect 312951 320179 313017 320182
rect 313230 319837 313290 320182
rect 314326 320180 314332 320182
rect 314396 320180 314402 320244
rect 314510 320180 314516 320244
rect 314580 320242 314586 320244
rect 316263 320242 316329 320245
rect 316539 320244 316605 320245
rect 316534 320242 316540 320244
rect 314580 320240 316329 320242
rect 314580 320184 316268 320240
rect 316324 320184 316329 320240
rect 314580 320182 316329 320184
rect 316448 320182 316540 320242
rect 314580 320180 314586 320182
rect 314331 320179 314397 320180
rect 316263 320179 316329 320182
rect 316534 320180 316540 320182
rect 316604 320180 316610 320244
rect 317275 320242 317341 320245
rect 316772 320240 317341 320242
rect 316772 320184 317280 320240
rect 317336 320184 317341 320240
rect 316772 320182 317341 320184
rect 316539 320179 316605 320180
rect 315803 320104 315869 320109
rect 315803 320048 315808 320104
rect 315864 320048 315869 320104
rect 315803 320043 315869 320048
rect 315987 320104 316053 320109
rect 315987 320048 315992 320104
rect 316048 320048 316053 320104
rect 315987 320043 316053 320048
rect 316171 320104 316237 320109
rect 316171 320048 316176 320104
rect 316232 320048 316237 320104
rect 316171 320043 316237 320048
rect 313181 319832 313290 319837
rect 313181 319776 313186 319832
rect 313242 319776 313290 319832
rect 313181 319774 313290 319776
rect 313181 319771 313247 319774
rect 312629 319696 312695 319701
rect 312629 319640 312634 319696
rect 312690 319640 312695 319696
rect 312629 319635 312695 319640
rect 313273 319698 313339 319701
rect 313457 319698 313523 319701
rect 313273 319696 313523 319698
rect 313273 319640 313278 319696
rect 313334 319640 313462 319696
rect 313518 319640 313523 319696
rect 313273 319638 313523 319640
rect 313273 319635 313339 319638
rect 313457 319635 313523 319638
rect 313825 319698 313891 319701
rect 314326 319698 314332 319700
rect 313825 319696 314332 319698
rect 313825 319640 313830 319696
rect 313886 319640 314332 319696
rect 313825 319638 314332 319640
rect 313825 319635 313891 319638
rect 314326 319636 314332 319638
rect 314396 319636 314402 319700
rect 314745 319698 314811 319701
rect 315806 319698 315866 320043
rect 314745 319696 315866 319698
rect 314745 319640 314750 319696
rect 314806 319640 315866 319696
rect 314745 319638 315866 319640
rect 314745 319635 314811 319638
rect 315990 319565 316050 320043
rect 312445 319560 312554 319565
rect 312445 319504 312450 319560
rect 312506 319504 312554 319560
rect 312445 319502 312554 319504
rect 312997 319562 313063 319565
rect 313406 319562 313412 319564
rect 312997 319560 313412 319562
rect 312997 319504 313002 319560
rect 313058 319504 313412 319560
rect 312997 319502 313412 319504
rect 312445 319499 312511 319502
rect 312997 319499 313063 319502
rect 313406 319500 313412 319502
rect 313476 319500 313482 319564
rect 315941 319560 316050 319565
rect 315941 319504 315946 319560
rect 316002 319504 316050 319560
rect 315941 319502 316050 319504
rect 316174 319562 316234 320043
rect 316772 319834 316832 320182
rect 317275 320179 317341 320182
rect 318379 320242 318445 320245
rect 319294 320242 319300 320244
rect 318379 320240 318810 320242
rect 318379 320184 318384 320240
rect 318440 320184 318810 320240
rect 318379 320182 318810 320184
rect 318379 320179 318445 320182
rect 316902 320044 316908 320108
rect 316972 320106 316978 320108
rect 317183 320106 317249 320109
rect 316972 320104 317249 320106
rect 316972 320048 317188 320104
rect 317244 320048 317249 320104
rect 316972 320046 317249 320048
rect 316972 320044 316978 320046
rect 317183 320043 317249 320046
rect 317459 320104 317525 320109
rect 317459 320048 317464 320104
rect 317520 320048 317525 320104
rect 317459 320043 317525 320048
rect 318103 320106 318169 320109
rect 318374 320106 318380 320108
rect 318103 320104 318380 320106
rect 318103 320048 318108 320104
rect 318164 320048 318380 320104
rect 318103 320046 318380 320048
rect 318103 320043 318169 320046
rect 318374 320044 318380 320046
rect 318444 320044 318450 320108
rect 318563 320104 318629 320109
rect 318563 320048 318568 320104
rect 318624 320048 318629 320104
rect 318563 320043 318629 320048
rect 317045 319834 317111 319837
rect 316772 319832 317111 319834
rect 316772 319776 317050 319832
rect 317106 319776 317111 319832
rect 316772 319774 317111 319776
rect 317045 319771 317111 319774
rect 316309 319698 316375 319701
rect 316309 319696 317292 319698
rect 316309 319640 316314 319696
rect 316370 319640 317292 319696
rect 316309 319638 317292 319640
rect 316309 319635 316375 319638
rect 317232 319565 317292 319638
rect 316493 319562 316559 319565
rect 316174 319560 316559 319562
rect 316174 319504 316498 319560
rect 316554 319504 316559 319560
rect 316174 319502 316559 319504
rect 315941 319499 316007 319502
rect 316493 319499 316559 319502
rect 316769 319562 316835 319565
rect 316902 319562 316908 319564
rect 316769 319560 316908 319562
rect 316769 319504 316774 319560
rect 316830 319504 316908 319560
rect 316769 319502 316908 319504
rect 316769 319499 316835 319502
rect 316902 319500 316908 319502
rect 316972 319500 316978 319564
rect 317229 319560 317295 319565
rect 317229 319504 317234 319560
rect 317290 319504 317295 319560
rect 317229 319499 317295 319504
rect 316718 319426 316724 319428
rect 312310 319366 316724 319426
rect 316718 319364 316724 319366
rect 316788 319364 316794 319428
rect 317462 319426 317522 320043
rect 317735 319936 317801 319939
rect 317735 319934 317936 319936
rect 317735 319878 317740 319934
rect 317796 319878 317936 319934
rect 317735 319876 317936 319878
rect 317735 319873 317801 319876
rect 317597 319698 317663 319701
rect 317876 319698 317936 319876
rect 317597 319696 317936 319698
rect 317597 319640 317602 319696
rect 317658 319640 317936 319696
rect 317597 319638 317936 319640
rect 318057 319698 318123 319701
rect 318425 319698 318491 319701
rect 318057 319696 318491 319698
rect 318057 319640 318062 319696
rect 318118 319640 318430 319696
rect 318486 319640 318491 319696
rect 318057 319638 318491 319640
rect 317597 319635 317663 319638
rect 318057 319635 318123 319638
rect 318425 319635 318491 319638
rect 317873 319562 317939 319565
rect 318566 319562 318626 320043
rect 318750 319701 318810 320182
rect 319256 320180 319300 320242
rect 319364 320180 319370 320244
rect 319662 320180 319668 320244
rect 319732 320242 319738 320244
rect 320127 320242 320193 320245
rect 319732 320240 320193 320242
rect 319732 320184 320132 320240
rect 320188 320184 320193 320240
rect 319732 320182 320193 320184
rect 319732 320180 319738 320182
rect 319256 320109 319316 320180
rect 320127 320179 320193 320182
rect 319207 320104 319316 320109
rect 319207 320048 319212 320104
rect 319268 320048 319316 320104
rect 319207 320046 319316 320048
rect 319391 320106 319457 320109
rect 319391 320104 319592 320106
rect 319391 320048 319396 320104
rect 319452 320048 319592 320104
rect 319391 320046 319592 320048
rect 319207 320043 319273 320046
rect 319391 320043 319457 320046
rect 319532 319701 319592 320046
rect 319851 320104 319917 320109
rect 319851 320048 319856 320104
rect 319912 320048 319917 320104
rect 319851 320043 319917 320048
rect 320035 320104 320101 320109
rect 320035 320048 320040 320104
rect 320096 320048 320101 320104
rect 320035 320043 320101 320048
rect 320403 320104 320469 320109
rect 320403 320048 320408 320104
rect 320464 320048 320469 320104
rect 320403 320043 320469 320048
rect 319667 319832 319733 319837
rect 319667 319776 319672 319832
rect 319728 319776 319733 319832
rect 319667 319771 319733 319776
rect 318701 319696 318810 319701
rect 318701 319640 318706 319696
rect 318762 319640 318810 319696
rect 318701 319638 318810 319640
rect 319529 319696 319595 319701
rect 319529 319640 319534 319696
rect 319590 319640 319595 319696
rect 318701 319635 318767 319638
rect 319529 319635 319595 319640
rect 317873 319560 318626 319562
rect 317873 319504 317878 319560
rect 317934 319504 318626 319560
rect 317873 319502 318626 319504
rect 318977 319562 319043 319565
rect 319161 319562 319227 319565
rect 318977 319560 319227 319562
rect 318977 319504 318982 319560
rect 319038 319504 319166 319560
rect 319222 319504 319227 319560
rect 318977 319502 319227 319504
rect 319670 319562 319730 319771
rect 319854 319701 319914 320043
rect 320038 319837 320098 320043
rect 319989 319832 320098 319837
rect 319989 319776 319994 319832
rect 320050 319776 320098 319832
rect 319989 319774 320098 319776
rect 319989 319771 320055 319774
rect 319805 319696 319914 319701
rect 319805 319640 319810 319696
rect 319866 319640 319914 319696
rect 319805 319638 319914 319640
rect 319805 319635 319871 319638
rect 319805 319562 319871 319565
rect 319670 319560 319871 319562
rect 319670 319504 319810 319560
rect 319866 319504 319871 319560
rect 319670 319502 319871 319504
rect 320406 319562 320466 320043
rect 320636 319701 320696 320318
rect 323158 320316 323164 320318
rect 323228 320316 323234 320380
rect 326659 320378 326725 320381
rect 338665 320378 338731 320381
rect 326659 320376 338731 320378
rect 326659 320320 326664 320376
rect 326720 320320 338670 320376
rect 338726 320320 338731 320376
rect 326659 320318 338731 320320
rect 323163 320315 323229 320316
rect 326659 320315 326725 320318
rect 338665 320315 338731 320318
rect 321415 320242 321481 320245
rect 322059 320244 322125 320245
rect 321686 320242 321692 320244
rect 321415 320240 321692 320242
rect 321415 320184 321420 320240
rect 321476 320184 321692 320240
rect 321415 320182 321692 320184
rect 321415 320179 321481 320182
rect 321686 320180 321692 320182
rect 321756 320180 321762 320244
rect 322054 320242 322060 320244
rect 321968 320182 322060 320242
rect 322054 320180 322060 320182
rect 322124 320180 322130 320244
rect 323071 320242 323137 320245
rect 324078 320242 324084 320244
rect 323071 320240 324084 320242
rect 323071 320184 323076 320240
rect 323132 320184 324084 320240
rect 323071 320182 324084 320184
rect 322059 320179 322125 320180
rect 323071 320179 323137 320182
rect 324078 320180 324084 320182
rect 324148 320180 324154 320244
rect 324267 320240 324333 320245
rect 324267 320184 324272 320240
rect 324328 320184 324333 320240
rect 324267 320179 324333 320184
rect 326107 320242 326173 320245
rect 334341 320242 334407 320245
rect 326107 320240 334407 320242
rect 326107 320184 326112 320240
rect 326168 320184 334346 320240
rect 334402 320184 334407 320240
rect 326107 320182 334407 320184
rect 326107 320179 326173 320182
rect 334341 320179 334407 320182
rect 321139 320104 321205 320109
rect 321139 320048 321144 320104
rect 321200 320048 321205 320104
rect 321139 320043 321205 320048
rect 321507 320104 321573 320109
rect 322151 320106 322217 320109
rect 321507 320048 321512 320104
rect 321568 320048 321573 320104
rect 321507 320043 321573 320048
rect 321878 320104 322217 320106
rect 321878 320048 322156 320104
rect 322212 320048 322217 320104
rect 321878 320046 322217 320048
rect 320633 319696 320699 319701
rect 320633 319640 320638 319696
rect 320694 319640 320699 319696
rect 320633 319635 320699 319640
rect 321142 319698 321202 320043
rect 321277 319698 321343 319701
rect 321142 319696 321343 319698
rect 321142 319640 321282 319696
rect 321338 319640 321343 319696
rect 321142 319638 321343 319640
rect 321277 319635 321343 319638
rect 320633 319562 320699 319565
rect 320406 319560 320699 319562
rect 320406 319504 320638 319560
rect 320694 319504 320699 319560
rect 320406 319502 320699 319504
rect 317873 319499 317939 319502
rect 318977 319499 319043 319502
rect 319161 319499 319227 319502
rect 319805 319499 319871 319502
rect 320633 319499 320699 319502
rect 321093 319562 321159 319565
rect 321510 319562 321570 320043
rect 321093 319560 321570 319562
rect 321093 319504 321098 319560
rect 321154 319504 321570 319560
rect 321093 319502 321570 319504
rect 321878 319562 321938 320046
rect 322151 320043 322217 320046
rect 322611 320104 322677 320109
rect 322611 320048 322616 320104
rect 322672 320048 322677 320104
rect 322611 320043 322677 320048
rect 323342 320044 323348 320108
rect 323412 320106 323418 320108
rect 323623 320106 323689 320109
rect 323412 320104 323689 320106
rect 323412 320048 323628 320104
rect 323684 320048 323689 320104
rect 323412 320046 323689 320048
rect 323412 320044 323418 320046
rect 323623 320043 323689 320046
rect 323894 320044 323900 320108
rect 323964 320106 323970 320108
rect 324083 320106 324149 320109
rect 323964 320104 324149 320106
rect 323964 320048 324088 320104
rect 324144 320048 324149 320104
rect 323964 320046 324149 320048
rect 323964 320044 323970 320046
rect 324083 320043 324149 320046
rect 322614 319970 322674 320043
rect 322246 319939 322490 319970
rect 322243 319934 322490 319939
rect 322243 319878 322248 319934
rect 322304 319910 322490 319934
rect 322614 319910 322858 319970
rect 322304 319878 322309 319910
rect 322243 319873 322309 319878
rect 322430 319834 322490 319910
rect 322657 319834 322723 319837
rect 322430 319832 322723 319834
rect 322430 319776 322662 319832
rect 322718 319776 322723 319832
rect 322430 319774 322723 319776
rect 322798 319834 322858 319910
rect 322798 319774 323042 319834
rect 322657 319771 322723 319774
rect 322105 319698 322171 319701
rect 322790 319698 322796 319700
rect 322105 319696 322796 319698
rect 322105 319640 322110 319696
rect 322166 319640 322796 319696
rect 322105 319638 322796 319640
rect 322105 319635 322171 319638
rect 322790 319636 322796 319638
rect 322860 319636 322866 319700
rect 322013 319562 322079 319565
rect 321878 319560 322079 319562
rect 321878 319504 322018 319560
rect 322074 319504 322079 319560
rect 321878 319502 322079 319504
rect 321093 319499 321159 319502
rect 322013 319499 322079 319502
rect 322238 319500 322244 319564
rect 322308 319562 322314 319564
rect 322381 319562 322447 319565
rect 322308 319560 322447 319562
rect 322308 319504 322386 319560
rect 322442 319504 322447 319560
rect 322308 319502 322447 319504
rect 322308 319500 322314 319502
rect 322381 319499 322447 319502
rect 322841 319562 322907 319565
rect 322982 319562 323042 319774
rect 323669 319698 323735 319701
rect 324270 319698 324330 320179
rect 326383 320106 326449 320109
rect 326935 320106 327001 320109
rect 338389 320106 338455 320109
rect 326383 320104 326722 320106
rect 326383 320048 326388 320104
rect 326444 320048 326722 320104
rect 326383 320046 326722 320048
rect 326383 320043 326449 320046
rect 326662 319970 326722 320046
rect 326935 320104 338455 320106
rect 326935 320048 326940 320104
rect 326996 320048 338394 320104
rect 338450 320048 338455 320104
rect 326935 320046 338455 320048
rect 326935 320043 327001 320046
rect 338389 320043 338455 320046
rect 328637 319970 328703 319973
rect 326662 319968 328703 319970
rect 325187 319934 325253 319939
rect 325187 319878 325192 319934
rect 325248 319878 325253 319934
rect 326662 319912 328642 319968
rect 328698 319912 328703 319968
rect 326662 319910 328703 319912
rect 328637 319907 328703 319910
rect 325187 319873 325253 319878
rect 323669 319696 324330 319698
rect 323669 319640 323674 319696
rect 323730 319640 324330 319696
rect 323669 319638 324330 319640
rect 324497 319698 324563 319701
rect 325190 319698 325250 319873
rect 326981 319834 327047 319837
rect 324497 319696 325250 319698
rect 324497 319640 324502 319696
rect 324558 319640 325250 319696
rect 324497 319638 325250 319640
rect 326846 319832 327047 319834
rect 326846 319776 326986 319832
rect 327042 319776 327047 319832
rect 326846 319774 327047 319776
rect 323669 319635 323735 319638
rect 324497 319635 324563 319638
rect 322841 319560 323042 319562
rect 322841 319504 322846 319560
rect 322902 319504 323042 319560
rect 322841 319502 323042 319504
rect 322841 319499 322907 319502
rect 323158 319500 323164 319564
rect 323228 319562 323234 319564
rect 323393 319562 323459 319565
rect 323228 319560 323459 319562
rect 323228 319504 323398 319560
rect 323454 319504 323459 319560
rect 323228 319502 323459 319504
rect 323228 319500 323234 319502
rect 323393 319499 323459 319502
rect 326705 319562 326771 319565
rect 326846 319562 326906 319774
rect 326981 319771 327047 319774
rect 326705 319560 326906 319562
rect 326705 319504 326710 319560
rect 326766 319504 326906 319560
rect 326705 319502 326906 319504
rect 326705 319499 326771 319502
rect 318057 319426 318123 319429
rect 317462 319424 318123 319426
rect 317462 319368 318062 319424
rect 318118 319368 318123 319424
rect 317462 319366 318123 319368
rect 318057 319363 318123 319366
rect 318374 319364 318380 319428
rect 318444 319426 318450 319428
rect 318517 319426 318583 319429
rect 319621 319428 319687 319429
rect 323945 319428 324011 319429
rect 319621 319426 319668 319428
rect 318444 319424 318583 319426
rect 318444 319368 318522 319424
rect 318578 319368 318583 319424
rect 318444 319366 318583 319368
rect 319576 319424 319668 319426
rect 319576 319368 319626 319424
rect 319576 319366 319668 319368
rect 318444 319364 318450 319366
rect 318517 319363 318583 319366
rect 319621 319364 319668 319366
rect 319732 319364 319738 319428
rect 323342 319426 323348 319428
rect 321510 319366 323348 319426
rect 319621 319363 319687 319364
rect 305494 319290 305500 319292
rect 292530 319230 305500 319290
rect 305494 319228 305500 319230
rect 305564 319228 305570 319292
rect 306741 319290 306807 319293
rect 307150 319290 307156 319292
rect 306741 319288 307156 319290
rect 306741 319232 306746 319288
rect 306802 319232 307156 319288
rect 306741 319230 307156 319232
rect 306741 319227 306807 319230
rect 307150 319228 307156 319230
rect 307220 319228 307226 319292
rect 309225 319290 309291 319293
rect 309726 319290 309732 319292
rect 309225 319288 309732 319290
rect 309225 319232 309230 319288
rect 309286 319232 309732 319288
rect 309225 319230 309732 319232
rect 309225 319227 309291 319230
rect 309726 319228 309732 319230
rect 309796 319228 309802 319292
rect 309910 319228 309916 319292
rect 309980 319290 309986 319292
rect 310145 319290 310211 319293
rect 309980 319288 310211 319290
rect 309980 319232 310150 319288
rect 310206 319232 310211 319288
rect 309980 319230 310211 319232
rect 309980 319228 309986 319230
rect 310145 319227 310211 319230
rect 310605 319290 310671 319293
rect 311341 319292 311407 319293
rect 310830 319290 310836 319292
rect 310605 319288 310836 319290
rect 310605 319232 310610 319288
rect 310666 319232 310836 319288
rect 310605 319230 310836 319232
rect 310605 319227 310671 319230
rect 310830 319228 310836 319230
rect 310900 319228 310906 319292
rect 311341 319290 311388 319292
rect 311296 319288 311388 319290
rect 311296 319232 311346 319288
rect 311296 319230 311388 319232
rect 311341 319228 311388 319230
rect 311452 319228 311458 319292
rect 314653 319290 314719 319293
rect 320214 319290 320220 319292
rect 314653 319288 320220 319290
rect 314653 319232 314658 319288
rect 314714 319232 320220 319288
rect 314653 319230 320220 319232
rect 311341 319227 311407 319228
rect 314653 319227 314719 319230
rect 320214 319228 320220 319230
rect 320284 319228 320290 319292
rect 284201 319154 284267 319157
rect 321510 319154 321570 319366
rect 323342 319364 323348 319366
rect 323412 319364 323418 319428
rect 323894 319364 323900 319428
rect 323964 319426 324011 319428
rect 325233 319426 325299 319429
rect 331489 319426 331555 319429
rect 323964 319424 324056 319426
rect 324006 319368 324056 319424
rect 323964 319366 324056 319368
rect 325233 319424 331555 319426
rect 325233 319368 325238 319424
rect 325294 319368 331494 319424
rect 331550 319368 331555 319424
rect 325233 319366 331555 319368
rect 323964 319364 324011 319366
rect 323945 319363 324011 319364
rect 325233 319363 325299 319366
rect 331489 319363 331555 319366
rect 324221 319290 324287 319293
rect 334249 319290 334315 319293
rect 324221 319288 334315 319290
rect 324221 319232 324226 319288
rect 324282 319232 334254 319288
rect 334310 319232 334315 319288
rect 324221 319230 334315 319232
rect 324221 319227 324287 319230
rect 334249 319227 334315 319230
rect 284201 319152 321570 319154
rect 284201 319096 284206 319152
rect 284262 319096 321570 319152
rect 284201 319094 321570 319096
rect 284201 319091 284267 319094
rect 324078 319092 324084 319156
rect 324148 319154 324154 319156
rect 335629 319154 335695 319157
rect 324148 319152 335695 319154
rect 324148 319096 335634 319152
rect 335690 319096 335695 319152
rect 324148 319094 335695 319096
rect 324148 319092 324154 319094
rect 335629 319091 335695 319094
rect 246798 318956 246804 319020
rect 246868 319018 246874 319020
rect 306097 319018 306163 319021
rect 246868 319016 306163 319018
rect 246868 318960 306102 319016
rect 306158 318960 306163 319016
rect 246868 318958 306163 318960
rect 246868 318956 246874 318958
rect 306097 318955 306163 318958
rect 309777 319018 309843 319021
rect 310278 319018 310284 319020
rect 309777 319016 310284 319018
rect 309777 318960 309782 319016
rect 309838 318960 310284 319016
rect 309777 318958 310284 318960
rect 309777 318955 309843 318958
rect 310278 318956 310284 318958
rect 310348 318956 310354 319020
rect 310789 319018 310855 319021
rect 311198 319018 311204 319020
rect 310789 319016 311204 319018
rect 310789 318960 310794 319016
rect 310850 318960 311204 319016
rect 310789 318958 311204 318960
rect 310789 318955 310855 318958
rect 311198 318956 311204 318958
rect 311268 318956 311274 319020
rect 312629 319018 312695 319021
rect 313222 319018 313228 319020
rect 312629 319016 313228 319018
rect 312629 318960 312634 319016
rect 312690 318960 313228 319016
rect 312629 318958 313228 318960
rect 312629 318955 312695 318958
rect 313222 318956 313228 318958
rect 313292 318956 313298 319020
rect 316309 319018 316375 319021
rect 319069 319020 319135 319021
rect 316534 319018 316540 319020
rect 316309 319016 316540 319018
rect 316309 318960 316314 319016
rect 316370 318960 316540 319016
rect 316309 318958 316540 318960
rect 316309 318955 316375 318958
rect 316534 318956 316540 318958
rect 316604 318956 316610 319020
rect 319069 319018 319116 319020
rect 319024 319016 319116 319018
rect 319024 318960 319074 319016
rect 319024 318958 319116 318960
rect 319069 318956 319116 318958
rect 319180 318956 319186 319020
rect 324681 319018 324747 319021
rect 334157 319018 334223 319021
rect 324681 319016 334223 319018
rect 324681 318960 324686 319016
rect 324742 318960 334162 319016
rect 334218 318960 334223 319016
rect 324681 318958 334223 318960
rect 319069 318955 319135 318956
rect 324681 318955 324747 318958
rect 334157 318955 334223 318958
rect 232262 318820 232268 318884
rect 232332 318882 232338 318884
rect 291929 318882 291995 318885
rect 232332 318880 291995 318882
rect 232332 318824 291934 318880
rect 291990 318824 291995 318880
rect 232332 318822 291995 318824
rect 232332 318820 232338 318822
rect 291929 318819 291995 318822
rect 292062 318820 292068 318884
rect 292132 318882 292138 318884
rect 292205 318882 292271 318885
rect 292132 318880 292271 318882
rect 292132 318824 292210 318880
rect 292266 318824 292271 318880
rect 292132 318822 292271 318824
rect 292132 318820 292138 318822
rect 292205 318819 292271 318822
rect 293217 318882 293283 318885
rect 293350 318882 293356 318884
rect 293217 318880 293356 318882
rect 293217 318824 293222 318880
rect 293278 318824 293356 318880
rect 293217 318822 293356 318824
rect 293217 318819 293283 318822
rect 293350 318820 293356 318822
rect 293420 318820 293426 318884
rect 294229 318882 294295 318885
rect 294454 318882 294460 318884
rect 294229 318880 294460 318882
rect 294229 318824 294234 318880
rect 294290 318824 294460 318880
rect 294229 318822 294460 318824
rect 294229 318819 294295 318822
rect 294454 318820 294460 318822
rect 294524 318820 294530 318884
rect 294597 318882 294663 318885
rect 295006 318882 295012 318884
rect 294597 318880 295012 318882
rect 294597 318824 294602 318880
rect 294658 318824 295012 318880
rect 294597 318822 295012 318824
rect 294597 318819 294663 318822
rect 295006 318820 295012 318822
rect 295076 318820 295082 318884
rect 295926 318820 295932 318884
rect 295996 318882 296002 318884
rect 296437 318882 296503 318885
rect 296713 318884 296779 318885
rect 296662 318882 296668 318884
rect 295996 318880 296503 318882
rect 295996 318824 296442 318880
rect 296498 318824 296503 318880
rect 295996 318822 296503 318824
rect 296622 318822 296668 318882
rect 296732 318880 296779 318884
rect 296774 318824 296779 318880
rect 295996 318820 296002 318822
rect 296437 318819 296503 318822
rect 296662 318820 296668 318822
rect 296732 318820 296779 318824
rect 296846 318820 296852 318884
rect 296916 318882 296922 318884
rect 297173 318882 297239 318885
rect 296916 318880 297239 318882
rect 296916 318824 297178 318880
rect 297234 318824 297239 318880
rect 296916 318822 297239 318824
rect 296916 318820 296922 318822
rect 296713 318819 296779 318820
rect 297173 318819 297239 318822
rect 299013 318882 299079 318885
rect 299238 318882 299244 318884
rect 299013 318880 299244 318882
rect 299013 318824 299018 318880
rect 299074 318824 299244 318880
rect 299013 318822 299244 318824
rect 299013 318819 299079 318822
rect 299238 318820 299244 318822
rect 299308 318820 299314 318884
rect 299657 318882 299723 318885
rect 299790 318882 299796 318884
rect 299657 318880 299796 318882
rect 299657 318824 299662 318880
rect 299718 318824 299796 318880
rect 299657 318822 299796 318824
rect 299657 318819 299723 318822
rect 299790 318820 299796 318822
rect 299860 318820 299866 318884
rect 300526 318820 300532 318884
rect 300596 318882 300602 318884
rect 301037 318882 301103 318885
rect 300596 318880 301103 318882
rect 300596 318824 301042 318880
rect 301098 318824 301103 318880
rect 300596 318822 301103 318824
rect 300596 318820 300602 318822
rect 301037 318819 301103 318822
rect 304993 318882 305059 318885
rect 305678 318882 305684 318884
rect 304993 318880 305684 318882
rect 304993 318824 304998 318880
rect 305054 318824 305684 318880
rect 304993 318822 305684 318824
rect 304993 318819 305059 318822
rect 305678 318820 305684 318822
rect 305748 318820 305754 318884
rect 311985 318882 312051 318885
rect 312854 318882 312860 318884
rect 311985 318880 312860 318882
rect 311985 318824 311990 318880
rect 312046 318824 312860 318880
rect 311985 318822 312860 318824
rect 311985 318819 312051 318822
rect 312854 318820 312860 318822
rect 312924 318820 312930 318884
rect 321686 318820 321692 318884
rect 321756 318882 321762 318884
rect 332685 318882 332751 318885
rect 321756 318880 332751 318882
rect 321756 318824 332690 318880
rect 332746 318824 332751 318880
rect 321756 318822 332751 318824
rect 321756 318820 321762 318822
rect 332685 318819 332751 318822
rect 221917 318746 221983 318749
rect 282453 318746 282519 318749
rect 286685 318748 286751 318749
rect 286685 318746 286732 318748
rect 221917 318744 282519 318746
rect 221917 318688 221922 318744
rect 221978 318688 282458 318744
rect 282514 318688 282519 318744
rect 221917 318686 282519 318688
rect 286640 318744 286732 318746
rect 286640 318688 286690 318744
rect 286640 318686 286732 318688
rect 221917 318683 221983 318686
rect 282453 318683 282519 318686
rect 286685 318684 286732 318686
rect 286796 318684 286802 318748
rect 287094 318684 287100 318748
rect 287164 318746 287170 318748
rect 287789 318746 287855 318749
rect 287164 318744 287855 318746
rect 287164 318688 287794 318744
rect 287850 318688 287855 318744
rect 287164 318686 287855 318688
rect 287164 318684 287170 318686
rect 286685 318683 286751 318684
rect 287789 318683 287855 318686
rect 287973 318748 288039 318749
rect 287973 318744 288020 318748
rect 288084 318746 288090 318748
rect 287973 318688 287978 318744
rect 287973 318684 288020 318688
rect 288084 318686 288130 318746
rect 288084 318684 288090 318686
rect 288198 318684 288204 318748
rect 288268 318746 288274 318748
rect 288341 318746 288407 318749
rect 288268 318744 288407 318746
rect 288268 318688 288346 318744
rect 288402 318688 288407 318744
rect 288268 318686 288407 318688
rect 288268 318684 288274 318686
rect 287973 318683 288039 318684
rect 288341 318683 288407 318686
rect 288750 318684 288756 318748
rect 288820 318746 288826 318748
rect 288893 318746 288959 318749
rect 288820 318744 288959 318746
rect 288820 318688 288898 318744
rect 288954 318688 288959 318744
rect 288820 318686 288959 318688
rect 288820 318684 288826 318686
rect 288893 318683 288959 318686
rect 289486 318684 289492 318748
rect 289556 318746 289562 318748
rect 290089 318746 290155 318749
rect 289556 318744 290155 318746
rect 289556 318688 290094 318744
rect 290150 318688 290155 318744
rect 289556 318686 290155 318688
rect 289556 318684 289562 318686
rect 290089 318683 290155 318686
rect 290917 318746 290983 318749
rect 291142 318746 291148 318748
rect 290917 318744 291148 318746
rect 290917 318688 290922 318744
rect 290978 318688 291148 318744
rect 290917 318686 291148 318688
rect 290917 318683 290983 318686
rect 291142 318684 291148 318686
rect 291212 318684 291218 318748
rect 297909 318746 297975 318749
rect 292530 318744 297975 318746
rect 292530 318688 297914 318744
rect 297970 318688 297975 318744
rect 292530 318686 297975 318688
rect 220670 318548 220676 318612
rect 220740 318610 220746 318612
rect 277577 318610 277643 318613
rect 220740 318608 277643 318610
rect 220740 318552 277582 318608
rect 277638 318552 277643 318608
rect 220740 318550 277643 318552
rect 220740 318548 220746 318550
rect 277577 318547 277643 318550
rect 278405 318610 278471 318613
rect 282545 318610 282611 318613
rect 278405 318608 282611 318610
rect 278405 318552 278410 318608
rect 278466 318552 282550 318608
rect 282606 318552 282611 318608
rect 278405 318550 282611 318552
rect 278405 318547 278471 318550
rect 282545 318547 282611 318550
rect 282862 318548 282868 318612
rect 282932 318610 282938 318612
rect 292530 318610 292590 318686
rect 297909 318683 297975 318686
rect 298134 318684 298140 318748
rect 298204 318746 298210 318748
rect 298921 318746 298987 318749
rect 298204 318744 298987 318746
rect 298204 318688 298926 318744
rect 298982 318688 298987 318744
rect 298204 318686 298987 318688
rect 298204 318684 298210 318686
rect 298921 318683 298987 318686
rect 299054 318684 299060 318748
rect 299124 318746 299130 318748
rect 299197 318746 299263 318749
rect 299124 318744 299263 318746
rect 299124 318688 299202 318744
rect 299258 318688 299263 318744
rect 299124 318686 299263 318688
rect 299124 318684 299130 318686
rect 299197 318683 299263 318686
rect 301998 318684 302004 318748
rect 302068 318746 302074 318748
rect 302969 318746 303035 318749
rect 302068 318744 303035 318746
rect 302068 318688 302974 318744
rect 303030 318688 303035 318744
rect 302068 318686 303035 318688
rect 302068 318684 302074 318686
rect 302969 318683 303035 318686
rect 304390 318684 304396 318748
rect 304460 318746 304466 318748
rect 307334 318746 307340 318748
rect 304460 318686 307340 318746
rect 304460 318684 304466 318686
rect 307334 318684 307340 318686
rect 307404 318684 307410 318748
rect 310094 318684 310100 318748
rect 310164 318746 310170 318748
rect 314510 318746 314516 318748
rect 310164 318686 314516 318746
rect 310164 318684 310170 318686
rect 314510 318684 314516 318686
rect 314580 318684 314586 318748
rect 282932 318550 292590 318610
rect 282932 318548 282938 318550
rect 295926 318548 295932 318612
rect 295996 318610 296002 318612
rect 307845 318610 307911 318613
rect 295996 318608 307911 318610
rect 295996 318552 307850 318608
rect 307906 318552 307911 318608
rect 295996 318550 307911 318552
rect 295996 318548 296002 318550
rect 307845 318547 307911 318550
rect 317086 318548 317092 318612
rect 317156 318610 317162 318612
rect 317321 318610 317387 318613
rect 317156 318608 317387 318610
rect 317156 318552 317326 318608
rect 317382 318552 317387 318608
rect 317156 318550 317387 318552
rect 317156 318548 317162 318550
rect 317321 318547 317387 318550
rect 326521 318610 326587 318613
rect 327257 318610 327323 318613
rect 326521 318608 327323 318610
rect 326521 318552 326526 318608
rect 326582 318552 327262 318608
rect 327318 318552 327323 318608
rect 326521 318550 327323 318552
rect 326521 318547 326587 318550
rect 327257 318547 327323 318550
rect 212165 318474 212231 318477
rect 278405 318474 278471 318477
rect 289537 318474 289603 318477
rect 212165 318472 278330 318474
rect 212165 318416 212170 318472
rect 212226 318416 278330 318472
rect 212165 318414 278330 318416
rect 212165 318411 212231 318414
rect 212349 318338 212415 318341
rect 278270 318338 278330 318414
rect 278405 318472 289603 318474
rect 278405 318416 278410 318472
rect 278466 318416 289542 318472
rect 289598 318416 289603 318472
rect 278405 318414 289603 318416
rect 278405 318411 278471 318414
rect 289537 318411 289603 318414
rect 292614 318412 292620 318476
rect 292684 318474 292690 318476
rect 293585 318474 293651 318477
rect 292684 318472 293651 318474
rect 292684 318416 293590 318472
rect 293646 318416 293651 318472
rect 292684 318414 293651 318416
rect 292684 318412 292690 318414
rect 293585 318411 293651 318414
rect 296897 318474 296963 318477
rect 297950 318474 297956 318476
rect 296897 318472 297956 318474
rect 296897 318416 296902 318472
rect 296958 318416 297956 318472
rect 296897 318414 297956 318416
rect 296897 318411 296963 318414
rect 297950 318412 297956 318414
rect 298020 318412 298026 318476
rect 302969 318474 303035 318477
rect 307886 318474 307892 318476
rect 302969 318472 307892 318474
rect 302969 318416 302974 318472
rect 303030 318416 307892 318472
rect 302969 318414 307892 318416
rect 302969 318411 303035 318414
rect 307886 318412 307892 318414
rect 307956 318412 307962 318476
rect 319253 318474 319319 318477
rect 326613 318474 326679 318477
rect 334709 318474 334775 318477
rect 319253 318472 326354 318474
rect 319253 318416 319258 318472
rect 319314 318416 326354 318472
rect 319253 318414 326354 318416
rect 319253 318411 319319 318414
rect 283598 318338 283604 318340
rect 212349 318336 278146 318338
rect 212349 318280 212354 318336
rect 212410 318280 278146 318336
rect 212349 318278 278146 318280
rect 278270 318278 283604 318338
rect 212349 318275 212415 318278
rect 212073 318202 212139 318205
rect 277761 318202 277827 318205
rect 212073 318200 277827 318202
rect 212073 318144 212078 318200
rect 212134 318144 277766 318200
rect 277822 318144 277827 318200
rect 212073 318142 277827 318144
rect 278086 318202 278146 318278
rect 283598 318276 283604 318278
rect 283668 318276 283674 318340
rect 284017 318338 284083 318341
rect 292798 318338 292804 318340
rect 284017 318336 292804 318338
rect 284017 318280 284022 318336
rect 284078 318280 292804 318336
rect 284017 318278 292804 318280
rect 284017 318275 284083 318278
rect 292798 318276 292804 318278
rect 292868 318276 292874 318340
rect 299974 318276 299980 318340
rect 300044 318338 300050 318340
rect 302325 318338 302391 318341
rect 300044 318336 302391 318338
rect 300044 318280 302330 318336
rect 302386 318280 302391 318336
rect 300044 318278 302391 318280
rect 300044 318276 300050 318278
rect 302325 318275 302391 318278
rect 303470 318276 303476 318340
rect 303540 318338 303546 318340
rect 312997 318338 313063 318341
rect 303540 318336 313063 318338
rect 303540 318280 313002 318336
rect 313058 318280 313063 318336
rect 303540 318278 313063 318280
rect 303540 318276 303546 318278
rect 312997 318275 313063 318278
rect 318609 318338 318675 318341
rect 325417 318338 325483 318341
rect 318609 318336 325483 318338
rect 318609 318280 318614 318336
rect 318670 318280 325422 318336
rect 325478 318280 325483 318336
rect 318609 318278 325483 318280
rect 326294 318338 326354 318414
rect 326613 318472 334775 318474
rect 326613 318416 326618 318472
rect 326674 318416 334714 318472
rect 334770 318416 334775 318472
rect 326613 318414 334775 318416
rect 326613 318411 326679 318414
rect 334709 318411 334775 318414
rect 326294 318278 340890 318338
rect 318609 318275 318675 318278
rect 325417 318275 325483 318278
rect 281901 318202 281967 318205
rect 278086 318200 281967 318202
rect 278086 318144 281906 318200
rect 281962 318144 281967 318200
rect 278086 318142 281967 318144
rect 212073 318139 212139 318142
rect 277761 318139 277827 318142
rect 281901 318139 281967 318142
rect 282545 318202 282611 318205
rect 282862 318202 282868 318204
rect 282545 318200 282868 318202
rect 282545 318144 282550 318200
rect 282606 318144 282868 318200
rect 282545 318142 282868 318144
rect 282545 318139 282611 318142
rect 282862 318140 282868 318142
rect 282932 318140 282938 318204
rect 284201 318202 284267 318205
rect 287145 318202 287211 318205
rect 284201 318200 287211 318202
rect 284201 318144 284206 318200
rect 284262 318144 287150 318200
rect 287206 318144 287211 318200
rect 284201 318142 287211 318144
rect 284201 318139 284267 318142
rect 287145 318139 287211 318142
rect 288617 318202 288683 318205
rect 291142 318202 291148 318204
rect 288617 318200 291148 318202
rect 288617 318144 288622 318200
rect 288678 318144 291148 318200
rect 288617 318142 291148 318144
rect 288617 318139 288683 318142
rect 291142 318140 291148 318142
rect 291212 318140 291218 318204
rect 292430 318140 292436 318204
rect 292500 318202 292506 318204
rect 293493 318202 293559 318205
rect 292500 318200 293559 318202
rect 292500 318144 293498 318200
rect 293554 318144 293559 318200
rect 292500 318142 293559 318144
rect 292500 318140 292506 318142
rect 293493 318139 293559 318142
rect 303705 318202 303771 318205
rect 303838 318202 303844 318204
rect 303705 318200 303844 318202
rect 303705 318144 303710 318200
rect 303766 318144 303844 318200
rect 303705 318142 303844 318144
rect 303705 318139 303771 318142
rect 303838 318140 303844 318142
rect 303908 318140 303914 318204
rect 319161 318202 319227 318205
rect 331673 318202 331739 318205
rect 319161 318200 331739 318202
rect 319161 318144 319166 318200
rect 319222 318144 331678 318200
rect 331734 318144 331739 318200
rect 319161 318142 331739 318144
rect 319161 318139 319227 318142
rect 331673 318139 331739 318142
rect 212441 318066 212507 318069
rect 278405 318066 278471 318069
rect 212441 318064 278471 318066
rect 212441 318008 212446 318064
rect 212502 318008 278410 318064
rect 278466 318008 278471 318064
rect 212441 318006 278471 318008
rect 212441 318003 212507 318006
rect 278405 318003 278471 318006
rect 287145 318066 287211 318069
rect 291694 318066 291700 318068
rect 287145 318064 291700 318066
rect 287145 318008 287150 318064
rect 287206 318008 291700 318064
rect 287145 318006 291700 318008
rect 287145 318003 287211 318006
rect 291694 318004 291700 318006
rect 291764 318004 291770 318068
rect 325417 318066 325483 318069
rect 329189 318066 329255 318069
rect 325417 318064 329255 318066
rect 325417 318008 325422 318064
rect 325478 318008 329194 318064
rect 329250 318008 329255 318064
rect 325417 318006 329255 318008
rect 325417 318003 325483 318006
rect 329189 318003 329255 318006
rect 282361 317930 282427 317933
rect 283782 317930 283788 317932
rect 282361 317928 283788 317930
rect 282361 317872 282366 317928
rect 282422 317872 283788 317928
rect 282361 317870 283788 317872
rect 282361 317867 282427 317870
rect 283782 317868 283788 317870
rect 283852 317868 283858 317932
rect 284937 317930 285003 317933
rect 285622 317930 285628 317932
rect 284937 317928 285628 317930
rect 284937 317872 284942 317928
rect 284998 317872 285628 317928
rect 284937 317870 285628 317872
rect 284937 317867 285003 317870
rect 285622 317868 285628 317870
rect 285692 317868 285698 317932
rect 289537 317930 289603 317933
rect 294781 317932 294847 317933
rect 291878 317930 291884 317932
rect 289537 317928 291884 317930
rect 289537 317872 289542 317928
rect 289598 317872 291884 317928
rect 289537 317870 291884 317872
rect 289537 317867 289603 317870
rect 291878 317868 291884 317870
rect 291948 317868 291954 317932
rect 294781 317928 294828 317932
rect 294892 317930 294898 317932
rect 294781 317872 294786 317928
rect 294781 317868 294828 317872
rect 294892 317870 294938 317930
rect 294892 317868 294898 317870
rect 298502 317868 298508 317932
rect 298572 317930 298578 317932
rect 299473 317930 299539 317933
rect 298572 317928 299539 317930
rect 298572 317872 299478 317928
rect 299534 317872 299539 317928
rect 298572 317870 299539 317872
rect 298572 317868 298578 317870
rect 294781 317867 294847 317868
rect 299473 317867 299539 317870
rect 302734 317868 302740 317932
rect 302804 317930 302810 317932
rect 305913 317930 305979 317933
rect 302804 317928 305979 317930
rect 302804 317872 305918 317928
rect 305974 317872 305979 317928
rect 302804 317870 305979 317872
rect 302804 317868 302810 317870
rect 305913 317867 305979 317870
rect 306230 317868 306236 317932
rect 306300 317930 306306 317932
rect 308673 317930 308739 317933
rect 306300 317928 308739 317930
rect 306300 317872 308678 317928
rect 308734 317872 308739 317928
rect 306300 317870 308739 317872
rect 306300 317868 306306 317870
rect 308673 317867 308739 317870
rect 319294 317868 319300 317932
rect 319364 317930 319370 317932
rect 322473 317930 322539 317933
rect 319364 317928 322539 317930
rect 319364 317872 322478 317928
rect 322534 317872 322539 317928
rect 319364 317870 322539 317872
rect 319364 317868 319370 317870
rect 322473 317867 322539 317870
rect 277761 317794 277827 317797
rect 285765 317794 285831 317797
rect 277761 317792 285831 317794
rect 277761 317736 277766 317792
rect 277822 317736 285770 317792
rect 285826 317736 285831 317792
rect 277761 317734 285831 317736
rect 277761 317731 277827 317734
rect 285765 317731 285831 317734
rect 287789 317794 287855 317797
rect 290181 317794 290247 317797
rect 287789 317792 290247 317794
rect 287789 317736 287794 317792
rect 287850 317736 290186 317792
rect 290242 317736 290247 317792
rect 287789 317734 290247 317736
rect 287789 317731 287855 317734
rect 290181 317731 290247 317734
rect 302918 317732 302924 317796
rect 302988 317794 302994 317796
rect 305269 317794 305335 317797
rect 302988 317792 305335 317794
rect 302988 317736 305274 317792
rect 305330 317736 305335 317792
rect 302988 317734 305335 317736
rect 302988 317732 302994 317734
rect 305269 317731 305335 317734
rect 306046 317732 306052 317796
rect 306116 317794 306122 317796
rect 308489 317794 308555 317797
rect 306116 317792 308555 317794
rect 306116 317736 308494 317792
rect 308550 317736 308555 317792
rect 306116 317734 308555 317736
rect 306116 317732 306122 317734
rect 308489 317731 308555 317734
rect 314142 317732 314148 317796
rect 314212 317794 314218 317796
rect 314561 317794 314627 317797
rect 314212 317792 314627 317794
rect 314212 317736 314566 317792
rect 314622 317736 314627 317792
rect 314212 317734 314627 317736
rect 314212 317732 314218 317734
rect 314561 317731 314627 317734
rect 318006 317732 318012 317796
rect 318076 317794 318082 317796
rect 318742 317794 318748 317796
rect 318076 317734 318748 317794
rect 318076 317732 318082 317734
rect 318742 317732 318748 317734
rect 318812 317794 318818 317796
rect 325969 317794 326035 317797
rect 327717 317794 327783 317797
rect 318812 317734 321570 317794
rect 318812 317732 318818 317734
rect 284518 317596 284524 317660
rect 284588 317658 284594 317660
rect 285213 317658 285279 317661
rect 284588 317656 285279 317658
rect 284588 317600 285218 317656
rect 285274 317600 285279 317656
rect 284588 317598 285279 317600
rect 284588 317596 284594 317598
rect 285213 317595 285279 317598
rect 285990 317596 285996 317660
rect 286060 317658 286066 317660
rect 286961 317658 287027 317661
rect 286060 317656 287027 317658
rect 286060 317600 286966 317656
rect 287022 317600 287027 317656
rect 286060 317598 287027 317600
rect 286060 317596 286066 317598
rect 286961 317595 287027 317598
rect 289077 317658 289143 317661
rect 291326 317658 291332 317660
rect 289077 317656 291332 317658
rect 289077 317600 289082 317656
rect 289138 317600 291332 317656
rect 289077 317598 291332 317600
rect 289077 317595 289143 317598
rect 291326 317596 291332 317598
rect 291396 317596 291402 317660
rect 292849 317658 292915 317661
rect 294454 317658 294460 317660
rect 292849 317656 294460 317658
rect 292849 317600 292854 317656
rect 292910 317600 294460 317656
rect 292849 317598 294460 317600
rect 292849 317595 292915 317598
rect 294454 317596 294460 317598
rect 294524 317596 294530 317660
rect 303838 317596 303844 317660
rect 303908 317658 303914 317660
rect 304717 317658 304783 317661
rect 303908 317656 304783 317658
rect 303908 317600 304722 317656
rect 304778 317600 304783 317656
rect 303908 317598 304783 317600
rect 303908 317596 303914 317598
rect 304717 317595 304783 317598
rect 305085 317658 305151 317661
rect 305678 317658 305684 317660
rect 305085 317656 305684 317658
rect 305085 317600 305090 317656
rect 305146 317600 305684 317656
rect 305085 317598 305684 317600
rect 305085 317595 305151 317598
rect 305678 317596 305684 317598
rect 305748 317596 305754 317660
rect 306598 317596 306604 317660
rect 306668 317658 306674 317660
rect 307569 317658 307635 317661
rect 306668 317656 307635 317658
rect 306668 317600 307574 317656
rect 307630 317600 307635 317656
rect 306668 317598 307635 317600
rect 321510 317658 321570 317734
rect 325969 317792 327783 317794
rect 325969 317736 325974 317792
rect 326030 317736 327722 317792
rect 327778 317736 327783 317792
rect 325969 317734 327783 317736
rect 325969 317731 326035 317734
rect 327717 317731 327783 317734
rect 326613 317658 326679 317661
rect 321510 317656 326679 317658
rect 321510 317600 326618 317656
rect 326674 317600 326679 317656
rect 321510 317598 326679 317600
rect 306668 317596 306674 317598
rect 307569 317595 307635 317598
rect 326613 317595 326679 317598
rect 326797 317658 326863 317661
rect 326797 317656 328562 317658
rect 326797 317600 326802 317656
rect 326858 317600 328562 317656
rect 326797 317598 328562 317600
rect 326797 317595 326863 317598
rect 285622 317460 285628 317524
rect 285692 317522 285698 317524
rect 286133 317522 286199 317525
rect 285692 317520 286199 317522
rect 285692 317464 286138 317520
rect 286194 317464 286199 317520
rect 285692 317462 286199 317464
rect 285692 317460 285698 317462
rect 286133 317459 286199 317462
rect 287053 317522 287119 317525
rect 287278 317522 287284 317524
rect 287053 317520 287284 317522
rect 287053 317464 287058 317520
rect 287114 317464 287284 317520
rect 287053 317462 287284 317464
rect 287053 317459 287119 317462
rect 287278 317460 287284 317462
rect 287348 317460 287354 317524
rect 287462 317460 287468 317524
rect 287532 317522 287538 317524
rect 287697 317522 287763 317525
rect 287532 317520 287763 317522
rect 287532 317464 287702 317520
rect 287758 317464 287763 317520
rect 287532 317462 287763 317464
rect 287532 317460 287538 317462
rect 287697 317459 287763 317462
rect 288382 317460 288388 317524
rect 288452 317522 288458 317524
rect 288525 317522 288591 317525
rect 288452 317520 288591 317522
rect 288452 317464 288530 317520
rect 288586 317464 288591 317520
rect 288452 317462 288591 317464
rect 288452 317460 288458 317462
rect 288525 317459 288591 317462
rect 291285 317524 291351 317525
rect 291561 317524 291627 317525
rect 292665 317524 292731 317525
rect 291285 317520 291332 317524
rect 291396 317522 291402 317524
rect 291285 317464 291290 317520
rect 291285 317460 291332 317464
rect 291396 317462 291442 317522
rect 291396 317460 291402 317462
rect 291510 317460 291516 317524
rect 291580 317522 291627 317524
rect 292614 317522 292620 317524
rect 291580 317520 291672 317522
rect 291622 317464 291672 317520
rect 291580 317462 291672 317464
rect 292574 317462 292620 317522
rect 292684 317520 292731 317524
rect 295558 317522 295564 317524
rect 292726 317464 292731 317520
rect 291580 317460 291627 317462
rect 292614 317460 292620 317462
rect 292684 317460 292731 317464
rect 291285 317459 291351 317460
rect 291561 317459 291627 317460
rect 292665 317459 292731 317460
rect 294830 317462 295564 317522
rect 278313 317386 278379 317389
rect 294830 317386 294890 317462
rect 295558 317460 295564 317462
rect 295628 317460 295634 317524
rect 296161 317522 296227 317525
rect 297081 317522 297147 317525
rect 296161 317520 297147 317522
rect 296161 317464 296166 317520
rect 296222 317464 297086 317520
rect 297142 317464 297147 317520
rect 296161 317462 297147 317464
rect 296161 317459 296227 317462
rect 297081 317459 297147 317462
rect 299606 317460 299612 317524
rect 299676 317522 299682 317524
rect 300577 317522 300643 317525
rect 299676 317520 300643 317522
rect 299676 317464 300582 317520
rect 300638 317464 300643 317520
rect 299676 317462 300643 317464
rect 299676 317460 299682 317462
rect 300577 317459 300643 317462
rect 300945 317522 301011 317525
rect 301814 317522 301820 317524
rect 300945 317520 301820 317522
rect 300945 317464 300950 317520
rect 301006 317464 301820 317520
rect 300945 317462 301820 317464
rect 300945 317459 301011 317462
rect 301814 317460 301820 317462
rect 301884 317460 301890 317524
rect 304206 317460 304212 317524
rect 304276 317522 304282 317524
rect 305177 317522 305243 317525
rect 305545 317524 305611 317525
rect 305494 317522 305500 317524
rect 304276 317520 305243 317522
rect 304276 317464 305182 317520
rect 305238 317464 305243 317520
rect 304276 317462 305243 317464
rect 305454 317462 305500 317522
rect 305564 317520 305611 317524
rect 305606 317464 305611 317520
rect 304276 317460 304282 317462
rect 305177 317459 305243 317462
rect 305494 317460 305500 317462
rect 305564 317460 305611 317464
rect 306414 317460 306420 317524
rect 306484 317522 306490 317524
rect 307017 317522 307083 317525
rect 306484 317520 307083 317522
rect 306484 317464 307022 317520
rect 307078 317464 307083 317520
rect 306484 317462 307083 317464
rect 306484 317460 306490 317462
rect 305545 317459 305611 317460
rect 307017 317459 307083 317462
rect 311709 317524 311775 317525
rect 311709 317520 311756 317524
rect 311820 317522 311826 317524
rect 311709 317464 311714 317520
rect 311709 317460 311756 317464
rect 311820 317462 311866 317522
rect 311820 317460 311826 317462
rect 313774 317460 313780 317524
rect 313844 317522 313850 317524
rect 314377 317522 314443 317525
rect 313844 317520 314443 317522
rect 313844 317464 314382 317520
rect 314438 317464 314443 317520
rect 313844 317462 314443 317464
rect 313844 317460 313850 317462
rect 311709 317459 311775 317460
rect 314377 317459 314443 317462
rect 317454 317460 317460 317524
rect 317524 317522 317530 317524
rect 318333 317522 318399 317525
rect 317524 317520 318399 317522
rect 317524 317464 318338 317520
rect 318394 317464 318399 317520
rect 317524 317462 318399 317464
rect 317524 317460 317530 317462
rect 318333 317459 318399 317462
rect 327349 317522 327415 317525
rect 328310 317522 328316 317524
rect 327349 317520 328316 317522
rect 327349 317464 327354 317520
rect 327410 317464 328316 317520
rect 327349 317462 328316 317464
rect 327349 317459 327415 317462
rect 328310 317460 328316 317462
rect 328380 317460 328386 317524
rect 328502 317522 328562 317598
rect 332041 317522 332107 317525
rect 328502 317520 332107 317522
rect 328502 317464 332046 317520
rect 332102 317464 332107 317520
rect 328502 317462 332107 317464
rect 340830 317522 340890 318278
rect 475377 317522 475443 317525
rect 340830 317520 475443 317522
rect 340830 317464 475382 317520
rect 475438 317464 475443 317520
rect 340830 317462 475443 317464
rect 332041 317459 332107 317462
rect 475377 317459 475443 317462
rect 278313 317384 294890 317386
rect 278313 317328 278318 317384
rect 278374 317328 294890 317384
rect 278313 317326 294890 317328
rect 294965 317386 295031 317389
rect 298093 317386 298159 317389
rect 294965 317384 298159 317386
rect 294965 317328 294970 317384
rect 295026 317328 298098 317384
rect 298154 317328 298159 317384
rect 294965 317326 298159 317328
rect 278313 317323 278379 317326
rect 294965 317323 295031 317326
rect 298093 317323 298159 317326
rect 271137 317250 271203 317253
rect 326889 317250 326955 317253
rect 271137 317248 326955 317250
rect 271137 317192 271142 317248
rect 271198 317192 326894 317248
rect 326950 317192 326955 317248
rect 271137 317190 326955 317192
rect 271137 317187 271203 317190
rect 326889 317187 326955 317190
rect 226742 317052 226748 317116
rect 226812 317114 226818 317116
rect 286593 317114 286659 317117
rect 226812 317112 286659 317114
rect 226812 317056 286598 317112
rect 286654 317056 286659 317112
rect 226812 317054 286659 317056
rect 226812 317052 226818 317054
rect 286593 317051 286659 317054
rect 219249 316978 219315 316981
rect 284753 316978 284819 316981
rect 219249 316976 284819 316978
rect 219249 316920 219254 316976
rect 219310 316920 284758 316976
rect 284814 316920 284819 316976
rect 219249 316918 284819 316920
rect 219249 316915 219315 316918
rect 284753 316915 284819 316918
rect 273897 316842 273963 316845
rect 320633 316842 320699 316845
rect 488533 316842 488599 316845
rect 273897 316840 488599 316842
rect 273897 316784 273902 316840
rect 273958 316784 320638 316840
rect 320694 316784 488538 316840
rect 488594 316784 488599 316840
rect 273897 316782 488599 316784
rect 273897 316779 273963 316782
rect 320633 316779 320699 316782
rect 488533 316779 488599 316782
rect 215109 316706 215175 316709
rect 289813 316706 289879 316709
rect 215109 316704 289879 316706
rect 215109 316648 215114 316704
rect 215170 316648 289818 316704
rect 289874 316648 289879 316704
rect 215109 316646 289879 316648
rect 215109 316643 215175 316646
rect 289813 316643 289879 316646
rect 326889 316706 326955 316709
rect 569953 316706 570019 316709
rect 326889 316704 570019 316706
rect 326889 316648 326894 316704
rect 326950 316648 569958 316704
rect 570014 316648 570019 316704
rect 326889 316646 570019 316648
rect 326889 316643 326955 316646
rect 569953 316643 570019 316646
rect 217777 316570 217843 316573
rect 284201 316570 284267 316573
rect 217777 316568 284267 316570
rect 217777 316512 217782 316568
rect 217838 316512 284206 316568
rect 284262 316512 284267 316568
rect 217777 316510 284267 316512
rect 217777 316507 217843 316510
rect 284201 316507 284267 316510
rect 323669 316162 323735 316165
rect 538213 316162 538279 316165
rect 323669 316160 538279 316162
rect 323669 316104 323674 316160
rect 323730 316104 538218 316160
rect 538274 316104 538279 316160
rect 323669 316102 538279 316104
rect 323669 316099 323735 316102
rect 538213 316099 538279 316102
rect 271597 315890 271663 315893
rect 299422 315890 299428 315892
rect 271597 315888 299428 315890
rect 271597 315832 271602 315888
rect 271658 315832 299428 315888
rect 271597 315830 299428 315832
rect 271597 315827 271663 315830
rect 299422 315828 299428 315830
rect 299492 315828 299498 315892
rect 232078 315692 232084 315756
rect 232148 315754 232154 315756
rect 291009 315754 291075 315757
rect 232148 315752 291075 315754
rect 232148 315696 291014 315752
rect 291070 315696 291075 315752
rect 232148 315694 291075 315696
rect 232148 315692 232154 315694
rect 291009 315691 291075 315694
rect 292389 315754 292455 315757
rect 293033 315754 293099 315757
rect 292389 315752 293099 315754
rect 292389 315696 292394 315752
rect 292450 315696 293038 315752
rect 293094 315696 293099 315752
rect 292389 315694 293099 315696
rect 292389 315691 292455 315694
rect 293033 315691 293099 315694
rect 253422 315556 253428 315620
rect 253492 315618 253498 315620
rect 312905 315618 312971 315621
rect 253492 315616 312971 315618
rect 253492 315560 312910 315616
rect 312966 315560 312971 315616
rect 253492 315558 312971 315560
rect 253492 315556 253498 315558
rect 312905 315555 312971 315558
rect 223430 315420 223436 315484
rect 223500 315482 223506 315484
rect 238845 315482 238911 315485
rect 223500 315480 238911 315482
rect 223500 315424 238850 315480
rect 238906 315424 238911 315480
rect 223500 315422 238911 315424
rect 223500 315420 223506 315422
rect 238845 315419 238911 315422
rect 243486 315420 243492 315484
rect 243556 315482 243562 315484
rect 303337 315482 303403 315485
rect 243556 315480 303403 315482
rect 243556 315424 303342 315480
rect 303398 315424 303403 315480
rect 243556 315422 303403 315424
rect 243556 315420 243562 315422
rect 303337 315419 303403 315422
rect 217593 315346 217659 315349
rect 294270 315346 294276 315348
rect 217593 315344 294276 315346
rect 217593 315288 217598 315344
rect 217654 315288 294276 315344
rect 217593 315286 294276 315288
rect 217593 315283 217659 315286
rect 294270 315284 294276 315286
rect 294340 315284 294346 315348
rect 281993 315210 282059 315213
rect 299606 315210 299612 315212
rect 281993 315208 299612 315210
rect 281993 315152 281998 315208
rect 282054 315152 299612 315208
rect 281993 315150 299612 315152
rect 281993 315147 282059 315150
rect 299606 315148 299612 315150
rect 299676 315148 299682 315212
rect 275461 315074 275527 315077
rect 314101 315076 314167 315077
rect 294822 315074 294828 315076
rect 275461 315072 294828 315074
rect 275461 315016 275466 315072
rect 275522 315016 294828 315072
rect 275461 315014 294828 315016
rect 275461 315011 275527 315014
rect 294822 315012 294828 315014
rect 294892 315012 294898 315076
rect 314101 315074 314148 315076
rect 314056 315072 314148 315074
rect 314056 315016 314106 315072
rect 314056 315014 314148 315016
rect 314101 315012 314148 315014
rect 314212 315012 314218 315076
rect 314101 315011 314167 315012
rect 310462 314938 310468 314940
rect 309182 314878 310468 314938
rect 222694 314604 222700 314668
rect 222764 314666 222770 314668
rect 247217 314666 247283 314669
rect 222764 314664 247283 314666
rect 222764 314608 247222 314664
rect 247278 314608 247283 314664
rect 222764 314606 247283 314608
rect 222764 314604 222770 314606
rect 247217 314603 247283 314606
rect 268469 314666 268535 314669
rect 309182 314666 309242 314878
rect 310462 314876 310468 314878
rect 310532 314938 310538 314940
rect 358077 314938 358143 314941
rect 310532 314936 358143 314938
rect 310532 314880 358082 314936
rect 358138 314880 358143 314936
rect 310532 314878 358143 314880
rect 310532 314876 310538 314878
rect 358077 314875 358143 314878
rect 311014 314740 311020 314804
rect 311084 314802 311090 314804
rect 311709 314802 311775 314805
rect 373993 314802 374059 314805
rect 311084 314800 374059 314802
rect 311084 314744 311714 314800
rect 311770 314744 373998 314800
rect 374054 314744 374059 314800
rect 311084 314742 374059 314744
rect 311084 314740 311090 314742
rect 311709 314739 311775 314742
rect 373993 314739 374059 314742
rect 268469 314664 309242 314666
rect 268469 314608 268474 314664
rect 268530 314608 309242 314664
rect 268469 314606 309242 314608
rect 268469 314603 268535 314606
rect 217869 314530 217935 314533
rect 285806 314530 285812 314532
rect 217869 314528 285812 314530
rect 217869 314472 217874 314528
rect 217930 314472 285812 314528
rect 217869 314470 285812 314472
rect 217869 314467 217935 314470
rect 285806 314468 285812 314470
rect 285876 314468 285882 314532
rect 213545 314394 213611 314397
rect 289118 314394 289124 314396
rect 213545 314392 289124 314394
rect 213545 314336 213550 314392
rect 213606 314336 289124 314392
rect 213545 314334 289124 314336
rect 213545 314331 213611 314334
rect 289118 314332 289124 314334
rect 289188 314332 289194 314396
rect 216213 314258 216279 314261
rect 295374 314258 295380 314260
rect 216213 314256 295380 314258
rect 216213 314200 216218 314256
rect 216274 314200 295380 314256
rect 216213 314198 295380 314200
rect 216213 314195 216279 314198
rect 295374 314196 295380 314198
rect 295444 314196 295450 314260
rect 216489 314122 216555 314125
rect 296662 314122 296668 314124
rect 216489 314120 296668 314122
rect 216489 314064 216494 314120
rect 216550 314064 296668 314120
rect 216489 314062 296668 314064
rect 216489 314059 216555 314062
rect 296662 314060 296668 314062
rect 296732 314060 296738 314124
rect 216581 313986 216647 313989
rect 297030 313986 297036 313988
rect 216581 313984 297036 313986
rect 216581 313928 216586 313984
rect 216642 313928 297036 313984
rect 216581 313926 297036 313928
rect 216581 313923 216647 313926
rect 297030 313924 297036 313926
rect 297100 313924 297106 313988
rect 241278 312972 241284 313036
rect 241348 313034 241354 313036
rect 301497 313034 301563 313037
rect 241348 313032 301563 313034
rect 241348 312976 301502 313032
rect 301558 312976 301563 313032
rect 241348 312974 301563 312976
rect 241348 312972 241354 312974
rect 301497 312971 301563 312974
rect 238150 312836 238156 312900
rect 238220 312898 238226 312900
rect 298093 312898 298159 312901
rect 238220 312896 298159 312898
rect 238220 312840 298098 312896
rect 298154 312840 298159 312896
rect 238220 312838 298159 312840
rect 238220 312836 238226 312838
rect 298093 312835 298159 312838
rect 238334 312700 238340 312764
rect 238404 312762 238410 312764
rect 298553 312762 298619 312765
rect 238404 312760 298619 312762
rect 238404 312704 298558 312760
rect 298614 312704 298619 312760
rect 238404 312702 298619 312704
rect 238404 312700 238410 312702
rect 298553 312699 298619 312702
rect 238702 312564 238708 312628
rect 238772 312626 238778 312628
rect 300761 312626 300827 312629
rect 238772 312624 300827 312626
rect 238772 312568 300766 312624
rect 300822 312568 300827 312624
rect 238772 312566 300827 312568
rect 238772 312564 238778 312566
rect 300761 312563 300827 312566
rect 220445 312490 220511 312493
rect 298502 312490 298508 312492
rect 220445 312488 298508 312490
rect 220445 312432 220450 312488
rect 220506 312432 298508 312488
rect 220445 312430 298508 312432
rect 220445 312427 220511 312430
rect 298502 312428 298508 312430
rect 298572 312428 298578 312492
rect 242198 312292 242204 312356
rect 242268 312354 242274 312356
rect 301405 312354 301471 312357
rect 242268 312352 301471 312354
rect 242268 312296 301410 312352
rect 301466 312296 301471 312352
rect 242268 312294 301471 312296
rect 242268 312292 242274 312294
rect 301405 312291 301471 312294
rect 243302 312156 243308 312220
rect 243372 312218 243378 312220
rect 302969 312218 303035 312221
rect 243372 312216 303035 312218
rect 243372 312160 302974 312216
rect 303030 312160 303035 312216
rect 243372 312158 303035 312160
rect 243372 312156 243378 312158
rect 302969 312155 303035 312158
rect 288433 312082 288499 312085
rect 288566 312082 288572 312084
rect 288433 312080 288572 312082
rect 288433 312024 288438 312080
rect 288494 312024 288572 312080
rect 288433 312022 288572 312024
rect 288433 312019 288499 312022
rect 288566 312020 288572 312022
rect 288636 312020 288642 312084
rect 292573 312082 292639 312085
rect 292982 312082 292988 312084
rect 292573 312080 292988 312082
rect 292573 312024 292578 312080
rect 292634 312024 292988 312080
rect 292573 312022 292988 312024
rect 292573 312019 292639 312022
rect 292982 312020 292988 312022
rect 293052 312020 293058 312084
rect 311157 312082 311223 312085
rect 311750 312082 311756 312084
rect 311157 312080 311756 312082
rect 311157 312024 311162 312080
rect 311218 312024 311756 312080
rect 311157 312022 311756 312024
rect 311157 312019 311223 312022
rect 311750 312020 311756 312022
rect 311820 312082 311826 312084
rect 378133 312082 378199 312085
rect 311820 312080 378199 312082
rect 311820 312024 378138 312080
rect 378194 312024 378199 312080
rect 311820 312022 378199 312024
rect 311820 312020 311826 312022
rect 378133 312019 378199 312022
rect 580441 312082 580507 312085
rect 583520 312082 584960 312172
rect 580441 312080 584960 312082
rect 580441 312024 580446 312080
rect 580502 312024 584960 312080
rect 580441 312022 584960 312024
rect 580441 312019 580507 312022
rect 322054 311884 322060 311948
rect 322124 311946 322130 311948
rect 508497 311946 508563 311949
rect 322124 311944 508563 311946
rect 322124 311888 508502 311944
rect 508558 311888 508563 311944
rect 583520 311932 584960 312022
rect 322124 311886 508563 311888
rect 322124 311884 322130 311886
rect 508497 311883 508563 311886
rect 249374 311748 249380 311812
rect 249444 311810 249450 311812
rect 308673 311810 308739 311813
rect 249444 311808 308739 311810
rect 249444 311752 308678 311808
rect 308734 311752 308739 311808
rect 249444 311750 308739 311752
rect 249444 311748 249450 311750
rect 308673 311747 308739 311750
rect 247718 311612 247724 311676
rect 247788 311674 247794 311676
rect 308765 311674 308831 311677
rect 247788 311672 308831 311674
rect 247788 311616 308770 311672
rect 308826 311616 308831 311672
rect 247788 311614 308831 311616
rect 247788 311612 247794 311614
rect 308765 311611 308831 311614
rect 249558 311476 249564 311540
rect 249628 311538 249634 311540
rect 309961 311538 310027 311541
rect 249628 311536 310027 311538
rect 249628 311480 309966 311536
rect 310022 311480 310027 311536
rect 249628 311478 310027 311480
rect 249628 311476 249634 311478
rect 309961 311475 310027 311478
rect 246430 311340 246436 311404
rect 246500 311402 246506 311404
rect 307109 311402 307175 311405
rect 246500 311400 307175 311402
rect 246500 311344 307114 311400
rect 307170 311344 307175 311400
rect 246500 311342 307175 311344
rect 246500 311340 246506 311342
rect 307109 311339 307175 311342
rect 248086 311204 248092 311268
rect 248156 311266 248162 311268
rect 308029 311266 308095 311269
rect 248156 311264 308095 311266
rect 248156 311208 308034 311264
rect 308090 311208 308095 311264
rect 248156 311206 308095 311208
rect 248156 311204 248162 311206
rect 308029 311203 308095 311206
rect 249190 311068 249196 311132
rect 249260 311130 249266 311132
rect 310237 311130 310303 311133
rect 249260 311128 310303 311130
rect 249260 311072 310242 311128
rect 310298 311072 310303 311128
rect 249260 311070 310303 311072
rect 249260 311068 249266 311070
rect 310237 311067 310303 311070
rect 234470 310932 234476 310996
rect 234540 310994 234546 310996
rect 293493 310994 293559 310997
rect 234540 310992 293559 310994
rect 234540 310936 293498 310992
rect 293554 310936 293559 310992
rect 234540 310934 293559 310936
rect 234540 310932 234546 310934
rect 293493 310931 293559 310934
rect 282269 310450 282335 310453
rect 288934 310450 288940 310452
rect 282269 310448 288940 310450
rect 282269 310392 282274 310448
rect 282330 310392 288940 310448
rect 282269 310390 288940 310392
rect 282269 310387 282335 310390
rect 288934 310388 288940 310390
rect 289004 310388 289010 310452
rect 254710 310252 254716 310316
rect 254780 310314 254786 310316
rect 315573 310314 315639 310317
rect 254780 310312 315639 310314
rect 254780 310256 315578 310312
rect 315634 310256 315639 310312
rect 254780 310254 315639 310256
rect 254780 310252 254786 310254
rect 315573 310251 315639 310254
rect 253238 310116 253244 310180
rect 253308 310178 253314 310180
rect 314193 310178 314259 310181
rect 253308 310176 314259 310178
rect 253308 310120 314198 310176
rect 314254 310120 314259 310176
rect 253308 310118 314259 310120
rect 253308 310116 253314 310118
rect 314193 310115 314259 310118
rect 253054 309980 253060 310044
rect 253124 310042 253130 310044
rect 314285 310042 314351 310045
rect 253124 310040 314351 310042
rect 253124 309984 314290 310040
rect 314346 309984 314351 310040
rect 253124 309982 314351 309984
rect 253124 309980 253130 309982
rect 314285 309979 314351 309982
rect 215201 309906 215267 309909
rect 282269 309906 282335 309909
rect 215201 309904 282335 309906
rect 215201 309848 215206 309904
rect 215262 309848 282274 309904
rect 282330 309848 282335 309904
rect 215201 309846 282335 309848
rect 215201 309843 215267 309846
rect 282269 309843 282335 309846
rect 285673 309906 285739 309909
rect 285990 309906 285996 309908
rect 285673 309904 285996 309906
rect 285673 309848 285678 309904
rect 285734 309848 285996 309904
rect 285673 309846 285996 309848
rect 285673 309843 285739 309846
rect 285990 309844 285996 309846
rect 286060 309844 286066 309908
rect 214833 309770 214899 309773
rect 290590 309770 290596 309772
rect 214833 309768 290596 309770
rect 214833 309712 214838 309768
rect 214894 309712 290596 309768
rect 214833 309710 290596 309712
rect 214833 309707 214899 309710
rect 290590 309708 290596 309710
rect 290660 309708 290666 309772
rect 283649 309634 283715 309637
rect 291510 309634 291516 309636
rect 283649 309632 291516 309634
rect 283649 309576 283654 309632
rect 283710 309576 291516 309632
rect 283649 309574 291516 309576
rect 283649 309571 283715 309574
rect 291510 309572 291516 309574
rect 291580 309572 291586 309636
rect 252134 309436 252140 309500
rect 252204 309498 252210 309500
rect 312721 309498 312787 309501
rect 252204 309496 312787 309498
rect 252204 309440 312726 309496
rect 312782 309440 312787 309496
rect 252204 309438 312787 309440
rect 252204 309436 252210 309438
rect 312721 309435 312787 309438
rect 287145 309362 287211 309365
rect 287462 309362 287468 309364
rect 287145 309360 287468 309362
rect 287145 309304 287150 309360
rect 287206 309304 287468 309360
rect 287145 309302 287468 309304
rect 287145 309299 287211 309302
rect 287462 309300 287468 309302
rect 287532 309300 287538 309364
rect 230974 308620 230980 308684
rect 231044 308682 231050 308684
rect 289353 308682 289419 308685
rect 231044 308680 289419 308682
rect 231044 308624 289358 308680
rect 289414 308624 289419 308680
rect 231044 308622 289419 308624
rect 231044 308620 231050 308622
rect 289353 308619 289419 308622
rect 259310 308484 259316 308548
rect 259380 308546 259386 308548
rect 317689 308546 317755 308549
rect 259380 308544 317755 308546
rect 259380 308488 317694 308544
rect 317750 308488 317755 308544
rect 259380 308486 317755 308488
rect 259380 308484 259386 308486
rect 317689 308483 317755 308486
rect 259126 308348 259132 308412
rect 259196 308410 259202 308412
rect 319897 308410 319963 308413
rect 259196 308408 319963 308410
rect 259196 308352 319902 308408
rect 319958 308352 319963 308408
rect 259196 308350 319963 308352
rect 259196 308348 259202 308350
rect 319897 308347 319963 308350
rect 245510 307668 245516 307732
rect 245580 307730 245586 307732
rect 302918 307730 302924 307732
rect 245580 307670 302924 307730
rect 245580 307668 245586 307670
rect 302918 307668 302924 307670
rect 302988 307668 302994 307732
rect 230238 307532 230244 307596
rect 230308 307594 230314 307596
rect 290365 307594 290431 307597
rect 230308 307592 290431 307594
rect 230308 307536 290370 307592
rect 290426 307536 290431 307592
rect 230308 307534 290431 307536
rect 230308 307532 230314 307534
rect 290365 307531 290431 307534
rect 223062 307396 223068 307460
rect 223132 307458 223138 307460
rect 283281 307458 283347 307461
rect 223132 307456 283347 307458
rect 223132 307400 283286 307456
rect 283342 307400 283347 307456
rect 223132 307398 283347 307400
rect 223132 307396 223138 307398
rect 283281 307395 283347 307398
rect 230054 307260 230060 307324
rect 230124 307322 230130 307324
rect 290089 307322 290155 307325
rect 230124 307320 290155 307322
rect 230124 307264 290094 307320
rect 290150 307264 290155 307320
rect 230124 307262 290155 307264
rect 230124 307260 230130 307262
rect 290089 307259 290155 307262
rect 211981 307186 212047 307189
rect 284518 307186 284524 307188
rect 211981 307184 284524 307186
rect 211981 307128 211986 307184
rect 212042 307128 284524 307184
rect 211981 307126 284524 307128
rect 211981 307123 212047 307126
rect 284518 307124 284524 307126
rect 284588 307124 284594 307188
rect 286593 307186 286659 307189
rect 295742 307186 295748 307188
rect 286593 307184 295748 307186
rect 286593 307128 286598 307184
rect 286654 307128 295748 307184
rect 286593 307126 295748 307128
rect 286593 307123 286659 307126
rect 295742 307124 295748 307126
rect 295812 307124 295818 307188
rect 214465 307050 214531 307053
rect 298318 307050 298324 307052
rect 214465 307048 298324 307050
rect 214465 306992 214470 307048
rect 214526 306992 298324 307048
rect 214465 306990 298324 306992
rect 214465 306987 214531 306990
rect 298318 306988 298324 306990
rect 298388 306988 298394 307052
rect 238150 306852 238156 306916
rect 238220 306914 238226 306916
rect 238518 306914 238524 306916
rect 238220 306854 238524 306914
rect 238220 306852 238226 306854
rect 238518 306852 238524 306854
rect 238588 306852 238594 306916
rect 238661 306370 238727 306373
rect 238886 306370 238892 306372
rect 238616 306368 238892 306370
rect -960 306234 480 306324
rect 238616 306312 238666 306368
rect 238722 306312 238892 306368
rect 238616 306310 238892 306312
rect 238661 306307 238727 306310
rect 238886 306308 238892 306310
rect 238956 306308 238962 306372
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 240910 305628 240916 305692
rect 240980 305690 240986 305692
rect 299749 305690 299815 305693
rect 240980 305688 299815 305690
rect 240980 305632 299754 305688
rect 299810 305632 299815 305688
rect 240980 305630 299815 305632
rect 240980 305628 240986 305630
rect 299749 305627 299815 305630
rect 228214 304268 228220 304332
rect 228284 304330 228290 304332
rect 287278 304330 287284 304332
rect 228284 304270 287284 304330
rect 228284 304268 228290 304270
rect 287278 304268 287284 304270
rect 287348 304268 287354 304332
rect 227846 304132 227852 304196
rect 227916 304194 227922 304196
rect 289537 304194 289603 304197
rect 227916 304192 289603 304194
rect 227916 304136 289542 304192
rect 289598 304136 289603 304192
rect 227916 304134 289603 304136
rect 227916 304132 227922 304134
rect 289537 304131 289603 304134
rect 318609 304060 318675 304061
rect 318558 304058 318564 304060
rect 318518 303998 318564 304058
rect 318628 304056 318675 304060
rect 318670 304000 318675 304056
rect 318558 303996 318564 303998
rect 318628 303996 318675 304000
rect 318609 303995 318675 303996
rect 228030 302772 228036 302836
rect 228100 302834 228106 302836
rect 288065 302834 288131 302837
rect 228100 302832 288131 302834
rect 228100 302776 288070 302832
rect 288126 302776 288131 302832
rect 228100 302774 288131 302776
rect 228100 302772 228106 302774
rect 288065 302771 288131 302774
rect 327574 302228 327580 302292
rect 327644 302290 327650 302292
rect 574737 302290 574803 302293
rect 327644 302288 574803 302290
rect 327644 302232 574742 302288
rect 574798 302232 574803 302288
rect 327644 302230 574803 302232
rect 327644 302228 327650 302230
rect 574737 302227 574803 302230
rect 242014 300324 242020 300388
rect 242084 300386 242090 300388
rect 301313 300386 301379 300389
rect 242084 300384 301379 300386
rect 242084 300328 301318 300384
rect 301374 300328 301379 300384
rect 242084 300326 301379 300328
rect 242084 300324 242090 300326
rect 301313 300323 301379 300326
rect 251582 300188 251588 300252
rect 251652 300250 251658 300252
rect 313181 300250 313247 300253
rect 251652 300248 313247 300250
rect 251652 300192 313186 300248
rect 313242 300192 313247 300248
rect 251652 300190 313247 300192
rect 251652 300188 251658 300190
rect 313181 300187 313247 300190
rect 239254 300052 239260 300116
rect 239324 300114 239330 300116
rect 300485 300114 300551 300117
rect 239324 300112 300551 300114
rect 239324 300056 300490 300112
rect 300546 300056 300551 300112
rect 239324 300054 300551 300056
rect 239324 300052 239330 300054
rect 300485 300051 300551 300054
rect 227294 298692 227300 298756
rect 227364 298754 227370 298756
rect 287421 298754 287487 298757
rect 227364 298752 287487 298754
rect 227364 298696 287426 298752
rect 287482 298696 287487 298752
rect 227364 298694 287487 298696
rect 227364 298692 227370 298694
rect 287421 298691 287487 298694
rect 580441 298754 580507 298757
rect 583520 298754 584960 298844
rect 580441 298752 584960 298754
rect 580441 298696 580446 298752
rect 580502 298696 584960 298752
rect 580441 298694 584960 298696
rect 580441 298691 580507 298694
rect 583520 298604 584960 298694
rect 231526 297740 231532 297804
rect 231596 297802 231602 297804
rect 283925 297802 283991 297805
rect 231596 297800 283991 297802
rect 231596 297744 283930 297800
rect 283986 297744 283991 297800
rect 231596 297742 283991 297744
rect 231596 297740 231602 297742
rect 283925 297739 283991 297742
rect 224718 297604 224724 297668
rect 224788 297666 224794 297668
rect 283097 297666 283163 297669
rect 224788 297664 283163 297666
rect 224788 297608 283102 297664
rect 283158 297608 283163 297664
rect 224788 297606 283163 297608
rect 224788 297604 224794 297606
rect 283097 297603 283163 297606
rect 247902 297468 247908 297532
rect 247972 297530 247978 297532
rect 306598 297530 306604 297532
rect 247972 297470 306604 297530
rect 247972 297468 247978 297470
rect 306598 297468 306604 297470
rect 306668 297468 306674 297532
rect 231710 297332 231716 297396
rect 231780 297394 231786 297396
rect 291326 297394 291332 297396
rect 231780 297334 291332 297394
rect 231780 297332 231786 297334
rect 291326 297332 291332 297334
rect 291396 297332 291402 297396
rect 238661 296850 238727 296853
rect 238886 296850 238892 296852
rect 238616 296848 238892 296850
rect 238616 296792 238666 296848
rect 238722 296792 238892 296848
rect 238616 296790 238892 296792
rect 238661 296787 238727 296790
rect 238886 296788 238892 296790
rect 238956 296788 238962 296852
rect 238661 296714 238727 296717
rect 238616 296712 238770 296714
rect 238616 296656 238666 296712
rect 238722 296656 238770 296712
rect 238616 296654 238770 296656
rect 238661 296651 238770 296654
rect 238710 296580 238770 296651
rect 238702 296516 238708 296580
rect 238772 296516 238778 296580
rect 226558 296108 226564 296172
rect 226628 296170 226634 296172
rect 286225 296170 286291 296173
rect 226628 296168 286291 296170
rect 226628 296112 286230 296168
rect 286286 296112 286291 296168
rect 226628 296110 286291 296112
rect 226628 296108 226634 296110
rect 286225 296107 286291 296110
rect 228398 295972 228404 296036
rect 228468 296034 228474 296036
rect 287329 296034 287395 296037
rect 228468 296032 287395 296034
rect 228468 295976 287334 296032
rect 287390 295976 287395 296032
rect 228468 295974 287395 295976
rect 228468 295972 228474 295974
rect 287329 295971 287395 295974
rect 242709 294810 242775 294813
rect 275318 294810 275324 294812
rect 242709 294808 275324 294810
rect 242709 294752 242714 294808
rect 242770 294752 275324 294808
rect 242709 294750 275324 294752
rect 242709 294747 242775 294750
rect 275318 294748 275324 294750
rect 275388 294748 275394 294812
rect 229870 294612 229876 294676
rect 229940 294674 229946 294676
rect 283833 294674 283899 294677
rect 229940 294672 283899 294674
rect 229940 294616 283838 294672
rect 283894 294616 283899 294672
rect 229940 294614 283899 294616
rect 229940 294612 229946 294614
rect 283833 294611 283899 294614
rect 252870 294476 252876 294540
rect 252940 294538 252946 294540
rect 313549 294538 313615 294541
rect 252940 294536 313615 294538
rect 252940 294480 313554 294536
rect 313610 294480 313615 294536
rect 252940 294478 313615 294480
rect 252940 294476 252946 294478
rect 313549 294475 313615 294478
rect 241605 293314 241671 293317
rect 277894 293314 277900 293316
rect 241605 293312 277900 293314
rect -960 293178 480 293268
rect 241605 293256 241610 293312
rect 241666 293256 277900 293312
rect 241605 293254 277900 293256
rect 241605 293251 241671 293254
rect 277894 293252 277900 293254
rect 277964 293252 277970 293316
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 239029 293178 239095 293181
rect 278078 293178 278084 293180
rect 239029 293176 278084 293178
rect 239029 293120 239034 293176
rect 239090 293120 278084 293176
rect 239029 293118 278084 293120
rect 239029 293115 239095 293118
rect 278078 293116 278084 293118
rect 278148 293116 278154 293180
rect 252645 292090 252711 292093
rect 275134 292090 275140 292092
rect 252645 292088 275140 292090
rect 252645 292032 252650 292088
rect 252706 292032 275140 292088
rect 252645 292030 275140 292032
rect 252645 292027 252711 292030
rect 275134 292028 275140 292030
rect 275204 292028 275210 292092
rect 231158 291892 231164 291956
rect 231228 291954 231234 291956
rect 287237 291954 287303 291957
rect 231228 291952 287303 291954
rect 231228 291896 287242 291952
rect 287298 291896 287303 291952
rect 231228 291894 287303 291896
rect 231228 291892 231234 291894
rect 287237 291891 287303 291894
rect 242382 291756 242388 291820
rect 242452 291818 242458 291820
rect 300853 291818 300919 291821
rect 242452 291816 300919 291818
rect 242452 291760 300858 291816
rect 300914 291760 300919 291816
rect 242452 291758 300919 291760
rect 242452 291756 242458 291758
rect 300853 291755 300919 291758
rect 228725 291546 228791 291549
rect 263542 291546 263548 291548
rect 228725 291544 263548 291546
rect 228725 291488 228730 291544
rect 228786 291488 263548 291544
rect 228725 291486 263548 291488
rect 228725 291483 228791 291486
rect 263542 291484 263548 291486
rect 263612 291484 263618 291548
rect 206277 291410 206343 291413
rect 264329 291410 264395 291413
rect 206277 291408 264395 291410
rect 206277 291352 206282 291408
rect 206338 291352 264334 291408
rect 264390 291352 264395 291408
rect 206277 291350 264395 291352
rect 206277 291347 206343 291350
rect 264329 291347 264395 291350
rect 43437 291274 43503 291277
rect 265893 291274 265959 291277
rect 43437 291272 265959 291274
rect 43437 291216 43442 291272
rect 43498 291216 265898 291272
rect 265954 291216 265959 291272
rect 43437 291214 265959 291216
rect 43437 291211 43503 291214
rect 265893 291211 265959 291214
rect 226425 291138 226491 291141
rect 227621 291138 227687 291141
rect 226425 291136 227687 291138
rect 226425 291080 226430 291136
rect 226486 291080 227626 291136
rect 227682 291080 227687 291136
rect 226425 291078 227687 291080
rect 226425 291075 226491 291078
rect 227621 291075 227687 291078
rect 260598 290804 260604 290868
rect 260668 290866 260674 290868
rect 320633 290866 320699 290869
rect 260668 290864 320699 290866
rect 260668 290808 320638 290864
rect 320694 290808 320699 290864
rect 260668 290806 320699 290808
rect 260668 290804 260674 290806
rect 320633 290803 320699 290806
rect 226926 290668 226932 290732
rect 226996 290730 227002 290732
rect 287973 290730 288039 290733
rect 226996 290728 288039 290730
rect 226996 290672 287978 290728
rect 288034 290672 288039 290728
rect 226996 290670 288039 290672
rect 226996 290668 227002 290670
rect 287973 290667 288039 290670
rect 245326 290532 245332 290596
rect 245396 290594 245402 290596
rect 305678 290594 305684 290596
rect 245396 290534 305684 290594
rect 245396 290532 245402 290534
rect 305678 290532 305684 290534
rect 305748 290532 305754 290596
rect 257102 290396 257108 290460
rect 257172 290458 257178 290460
rect 317597 290458 317663 290461
rect 257172 290456 317663 290458
rect 257172 290400 317602 290456
rect 317658 290400 317663 290456
rect 257172 290398 317663 290400
rect 257172 290396 257178 290398
rect 317597 290395 317663 290398
rect 238661 290322 238727 290325
rect 238886 290322 238892 290324
rect 238616 290320 238892 290322
rect 238616 290264 238666 290320
rect 238722 290264 238892 290320
rect 238616 290262 238892 290264
rect 238661 290259 238727 290262
rect 238886 290260 238892 290262
rect 238956 290260 238962 290324
rect 224585 290050 224651 290053
rect 224542 290048 224651 290050
rect 224542 289992 224590 290048
rect 224646 289992 224651 290048
rect 224542 289987 224651 289992
rect 249006 289988 249012 290052
rect 249076 290050 249082 290052
rect 249609 290050 249675 290053
rect 249076 290048 249675 290050
rect 249076 289992 249614 290048
rect 249670 289992 249675 290048
rect 249076 289990 249675 289992
rect 249076 289988 249082 289990
rect 249609 289987 249675 289990
rect 250478 289988 250484 290052
rect 250548 290050 250554 290052
rect 250713 290050 250779 290053
rect 250548 290048 250779 290050
rect 250548 289992 250718 290048
rect 250774 289992 250779 290048
rect 250548 289990 250779 289992
rect 250548 289988 250554 289990
rect 250713 289987 250779 289990
rect 255446 289988 255452 290052
rect 255516 290050 255522 290052
rect 256509 290050 256575 290053
rect 255516 290048 256575 290050
rect 255516 289992 256514 290048
rect 256570 289992 256575 290048
rect 255516 289990 256575 289992
rect 255516 289988 255522 289990
rect 256509 289987 256575 289990
rect 223614 289716 223620 289780
rect 223684 289778 223690 289780
rect 224542 289778 224602 289987
rect 227621 289914 227687 289917
rect 269614 289914 269620 289916
rect 227621 289912 269620 289914
rect 227621 289856 227626 289912
rect 227682 289856 269620 289912
rect 227621 289854 269620 289856
rect 227621 289851 227687 289854
rect 269614 289852 269620 289854
rect 269684 289852 269690 289916
rect 223684 289718 224602 289778
rect 223684 289716 223690 289718
rect 231894 289716 231900 289780
rect 231964 289778 231970 289780
rect 233049 289778 233115 289781
rect 231964 289776 233115 289778
rect 231964 289720 233054 289776
rect 233110 289720 233115 289776
rect 231964 289718 233115 289720
rect 231964 289716 231970 289718
rect 233049 289715 233115 289718
rect 235206 289716 235212 289780
rect 235276 289778 235282 289780
rect 235625 289778 235691 289781
rect 235276 289776 235691 289778
rect 235276 289720 235630 289776
rect 235686 289720 235691 289776
rect 235276 289718 235691 289720
rect 235276 289716 235282 289718
rect 235625 289715 235691 289718
rect 250662 289716 250668 289780
rect 250732 289778 250738 289780
rect 251081 289778 251147 289781
rect 250732 289776 251147 289778
rect 250732 289720 251086 289776
rect 251142 289720 251147 289776
rect 250732 289718 251147 289720
rect 250732 289716 250738 289718
rect 251081 289715 251147 289718
rect 255630 289716 255636 289780
rect 255700 289778 255706 289780
rect 256233 289778 256299 289781
rect 255700 289776 256299 289778
rect 255700 289720 256238 289776
rect 256294 289720 256299 289776
rect 255700 289718 256299 289720
rect 255700 289716 255706 289718
rect 256233 289715 256299 289718
rect 256509 289778 256575 289781
rect 256509 289776 277410 289778
rect 256509 289720 256514 289776
rect 256570 289720 277410 289776
rect 256509 289718 277410 289720
rect 256509 289715 256575 289718
rect 223982 289580 223988 289644
rect 224052 289642 224058 289644
rect 224953 289642 225019 289645
rect 224052 289640 225019 289642
rect 224052 289584 224958 289640
rect 225014 289584 225019 289640
rect 224052 289582 225019 289584
rect 224052 289580 224058 289582
rect 224953 289579 225019 289582
rect 235390 289580 235396 289644
rect 235460 289642 235466 289644
rect 235901 289642 235967 289645
rect 250989 289642 251055 289645
rect 235460 289640 235967 289642
rect 235460 289584 235906 289640
rect 235962 289584 235967 289640
rect 235460 289582 235967 289584
rect 235460 289580 235466 289582
rect 235901 289579 235967 289582
rect 250854 289640 251055 289642
rect 250854 289584 250994 289640
rect 251050 289584 251055 289640
rect 250854 289582 251055 289584
rect 250294 289444 250300 289508
rect 250364 289506 250370 289508
rect 250854 289506 250914 289582
rect 250989 289579 251055 289582
rect 251766 289580 251772 289644
rect 251836 289642 251842 289644
rect 252553 289642 252619 289645
rect 251836 289640 252619 289642
rect 251836 289584 252558 289640
rect 252614 289584 252619 289640
rect 251836 289582 252619 289584
rect 251836 289580 251842 289582
rect 252553 289579 252619 289582
rect 255814 289580 255820 289644
rect 255884 289642 255890 289644
rect 256601 289642 256667 289645
rect 263869 289642 263935 289645
rect 255884 289640 256667 289642
rect 255884 289584 256606 289640
rect 256662 289584 256667 289640
rect 255884 289582 256667 289584
rect 255884 289580 255890 289582
rect 256601 289579 256667 289582
rect 258030 289640 263935 289642
rect 258030 289584 263874 289640
rect 263930 289584 263935 289640
rect 258030 289582 263935 289584
rect 250364 289446 250914 289506
rect 250364 289444 250370 289446
rect 186957 289234 187023 289237
rect 258030 289234 258090 289582
rect 263869 289579 263935 289582
rect 264973 289642 265039 289645
rect 264973 289640 265082 289642
rect 264973 289584 264978 289640
rect 265034 289584 265082 289640
rect 264973 289579 265082 289584
rect 265022 289370 265082 289579
rect 265157 289370 265223 289373
rect 186957 289232 258090 289234
rect 186957 289176 186962 289232
rect 187018 289176 258090 289232
rect 186957 289174 258090 289176
rect 262814 289368 265223 289370
rect 262814 289312 265162 289368
rect 265218 289312 265223 289368
rect 262814 289310 265223 289312
rect 186957 289171 187023 289174
rect 7557 289098 7623 289101
rect 262814 289098 262874 289310
rect 265157 289307 265223 289310
rect 7557 289096 262874 289098
rect 7557 289040 7562 289096
rect 7618 289040 262874 289096
rect 7557 289038 262874 289040
rect 277350 289098 277410 289718
rect 282678 289098 282684 289100
rect 277350 289038 282684 289098
rect 7557 289035 7623 289038
rect 282678 289036 282684 289038
rect 282748 289098 282754 289100
rect 580441 289098 580507 289101
rect 282748 289096 580507 289098
rect 282748 289040 580446 289096
rect 580502 289040 580507 289096
rect 282748 289038 580507 289040
rect 282748 289036 282754 289038
rect 580441 289035 580507 289038
rect 256182 287676 256188 287740
rect 256252 287738 256258 287740
rect 316401 287738 316467 287741
rect 256252 287736 316467 287738
rect 256252 287680 316406 287736
rect 316462 287680 316467 287736
rect 256252 287678 316467 287680
rect 256252 287676 256258 287678
rect 316401 287675 316467 287678
rect 263542 286996 263548 287060
rect 263612 287058 263618 287060
rect 281441 287058 281507 287061
rect 263612 287056 281507 287058
rect 263612 287000 281446 287056
rect 281502 287000 281507 287056
rect 263612 286998 281507 287000
rect 263612 286996 263618 286998
rect 281441 286995 281507 286998
rect 270125 286514 270191 286517
rect 318006 286514 318012 286516
rect 270125 286512 318012 286514
rect 270125 286456 270130 286512
rect 270186 286456 318012 286512
rect 270125 286454 318012 286456
rect 270125 286451 270191 286454
rect 318006 286452 318012 286454
rect 318076 286452 318082 286516
rect 281441 286378 281507 286381
rect 580625 286378 580691 286381
rect 281441 286376 580691 286378
rect 281441 286320 281446 286376
rect 281502 286320 580630 286376
rect 580686 286320 580691 286376
rect 281441 286318 580691 286320
rect 281441 286315 281507 286318
rect 580625 286315 580691 286318
rect 583520 285276 584960 285516
rect 284886 283460 284892 283524
rect 284956 283522 284962 283524
rect 418797 283522 418863 283525
rect 284956 283520 418863 283522
rect 284956 283464 418802 283520
rect 418858 283464 418863 283520
rect 284956 283462 418863 283464
rect 284956 283460 284962 283462
rect 418797 283459 418863 283462
rect -960 279972 480 280212
rect 267549 272506 267615 272509
rect 326981 272506 327047 272509
rect 267549 272504 327047 272506
rect 267549 272448 267554 272504
rect 267610 272448 326986 272504
rect 327042 272448 327047 272504
rect 267549 272446 327047 272448
rect 267549 272443 267615 272446
rect 326981 272443 327047 272446
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 266486 271084 266492 271148
rect 266556 271146 266562 271148
rect 326613 271146 326679 271149
rect 266556 271144 326679 271146
rect 266556 271088 326618 271144
rect 326674 271088 326679 271144
rect 266556 271086 326679 271088
rect 266556 271084 266562 271086
rect 326613 271083 326679 271086
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 267406 258844 267412 258908
rect 267476 258906 267482 258908
rect 327257 258906 327323 258909
rect 267476 258904 327323 258906
rect 267476 258848 327262 258904
rect 327318 258848 327323 258904
rect 267476 258846 327323 258848
rect 267476 258844 267482 258846
rect 327257 258843 327323 258846
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 263726 258708 263732 258772
rect 263796 258770 263802 258772
rect 324681 258770 324747 258773
rect 263796 258768 324747 258770
rect 263796 258712 324686 258768
rect 324742 258712 324747 258768
rect 583520 258756 584960 258846
rect 263796 258710 324747 258712
rect 263796 258708 263802 258710
rect 324681 258707 324747 258710
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 309869 254010 309935 254013
rect 310094 254010 310100 254012
rect 309869 254008 310100 254010
rect 309869 253952 309874 254008
rect 309930 253952 310100 254008
rect 309869 253950 310100 253952
rect 309869 253947 309935 253950
rect 310094 253948 310100 253950
rect 310164 254010 310170 254012
rect 434713 254010 434779 254013
rect 310164 254008 434779 254010
rect 310164 253952 434718 254008
rect 434774 253952 434779 254008
rect 310164 253950 434779 253952
rect 310164 253948 310170 253950
rect 434713 253947 434779 253950
rect 267641 250474 267707 250477
rect 325969 250474 326035 250477
rect 267641 250472 326035 250474
rect 267641 250416 267646 250472
rect 267702 250416 325974 250472
rect 326030 250416 326035 250472
rect 267641 250414 326035 250416
rect 267641 250411 267707 250414
rect 325969 250411 326035 250414
rect 264094 247692 264100 247756
rect 264164 247754 264170 247756
rect 288525 247754 288591 247757
rect 264164 247752 288591 247754
rect 264164 247696 288530 247752
rect 288586 247696 288591 247752
rect 264164 247694 288591 247696
rect 264164 247692 264170 247694
rect 288525 247691 288591 247694
rect 269297 247618 269363 247621
rect 327993 247618 328059 247621
rect 269297 247616 328059 247618
rect 269297 247560 269302 247616
rect 269358 247560 327998 247616
rect 328054 247560 328059 247616
rect 269297 247558 328059 247560
rect 269297 247555 269363 247558
rect 327993 247555 328059 247558
rect 267917 246258 267983 246261
rect 324589 246258 324655 246261
rect 267917 246256 324655 246258
rect 267917 246200 267922 246256
rect 267978 246200 324594 246256
rect 324650 246200 324655 246256
rect 267917 246198 324655 246200
rect 267917 246195 267983 246198
rect 324589 246195 324655 246198
rect 580717 245578 580783 245581
rect 583520 245578 584960 245668
rect 580717 245576 584960 245578
rect 580717 245520 580722 245576
rect 580778 245520 584960 245576
rect 580717 245518 584960 245520
rect 580717 245515 580783 245518
rect 583520 245428 584960 245518
rect 266118 244972 266124 245036
rect 266188 245034 266194 245036
rect 325877 245034 325943 245037
rect 266188 245032 325943 245034
rect 266188 244976 325882 245032
rect 325938 244976 325943 245032
rect 266188 244974 325943 244976
rect 266188 244972 266194 244974
rect 325877 244971 325943 244974
rect 263542 244836 263548 244900
rect 263612 244898 263618 244900
rect 323209 244898 323275 244901
rect 263612 244896 323275 244898
rect 263612 244840 323214 244896
rect 323270 244840 323275 244896
rect 263612 244838 323275 244840
rect 263612 244836 263618 244838
rect 323209 244835 323275 244838
rect 267549 244220 267615 244221
rect 267549 244216 267596 244220
rect 267660 244218 267666 244220
rect 267549 244160 267554 244216
rect 267549 244156 267596 244160
rect 267660 244158 267706 244218
rect 267660 244156 267666 244158
rect 267549 244155 267615 244156
rect 267549 244082 267615 244085
rect 319621 244082 319687 244085
rect 267549 244080 319687 244082
rect 267549 244024 267554 244080
rect 267610 244024 319626 244080
rect 319682 244024 319687 244080
rect 267549 244022 319687 244024
rect 267549 244019 267615 244022
rect 319621 244019 319687 244022
rect 264462 243884 264468 243948
rect 264532 243946 264538 243948
rect 324313 243946 324379 243949
rect 264532 243944 324379 243946
rect 264532 243888 324318 243944
rect 324374 243888 324379 243944
rect 264532 243886 324379 243888
rect 264532 243884 264538 243886
rect 324313 243883 324379 243886
rect 269481 243810 269547 243813
rect 325785 243810 325851 243813
rect 269481 243808 325851 243810
rect 269481 243752 269486 243808
rect 269542 243752 325790 243808
rect 325846 243752 325851 243808
rect 269481 243750 325851 243752
rect 269481 243747 269547 243750
rect 325785 243747 325851 243750
rect 268837 243674 268903 243677
rect 323117 243674 323183 243677
rect 268837 243672 323183 243674
rect 268837 243616 268842 243672
rect 268898 243616 323122 243672
rect 323178 243616 323183 243672
rect 268837 243614 323183 243616
rect 268837 243611 268903 243614
rect 323117 243611 323183 243614
rect 267825 243538 267891 243541
rect 327574 243538 327580 243540
rect 267825 243536 327580 243538
rect 267825 243480 267830 243536
rect 267886 243480 327580 243536
rect 267825 243478 327580 243480
rect 267825 243475 267891 243478
rect 327574 243476 327580 243478
rect 327644 243476 327650 243540
rect 264278 242252 264284 242316
rect 264348 242314 264354 242316
rect 269113 242314 269179 242317
rect 264348 242312 269179 242314
rect 264348 242256 269118 242312
rect 269174 242256 269179 242312
rect 264348 242254 269179 242256
rect 264348 242252 264354 242254
rect 269113 242251 269179 242254
rect 263726 242116 263732 242180
rect 263796 242178 263802 242180
rect 322054 242178 322060 242180
rect 263796 242118 322060 242178
rect 263796 242116 263802 242118
rect 322054 242116 322060 242118
rect 322124 242116 322130 242180
rect 260966 241980 260972 242044
rect 261036 242042 261042 242044
rect 321369 242042 321435 242045
rect 261036 242040 321435 242042
rect 261036 241984 321374 242040
rect 321430 241984 321435 242040
rect 261036 241982 321435 241984
rect 261036 241980 261042 241982
rect 321369 241979 321435 241982
rect 264646 241844 264652 241908
rect 264716 241906 264722 241908
rect 323945 241906 324011 241909
rect 264716 241904 324011 241906
rect 264716 241848 323950 241904
rect 324006 241848 324011 241904
rect 264716 241846 324011 241848
rect 264716 241844 264722 241846
rect 323945 241843 324011 241846
rect 239070 241708 239076 241772
rect 239140 241770 239146 241772
rect 298277 241770 298343 241773
rect 239140 241768 298343 241770
rect 239140 241712 298282 241768
rect 298338 241712 298343 241768
rect 239140 241710 298343 241712
rect 239140 241708 239146 241710
rect 298277 241707 298343 241710
rect 258758 241572 258764 241636
rect 258828 241634 258834 241636
rect 267549 241634 267615 241637
rect 258828 241632 267615 241634
rect 258828 241576 267554 241632
rect 267610 241576 267615 241632
rect 258828 241574 267615 241576
rect 258828 241572 258834 241574
rect 267549 241571 267615 241574
rect 246614 241436 246620 241500
rect 246684 241498 246690 241500
rect 302734 241498 302740 241500
rect 246684 241438 302740 241498
rect 246684 241436 246690 241438
rect 302734 241436 302740 241438
rect 302804 241436 302810 241500
rect 222285 241362 222351 241365
rect 223246 241362 223252 241364
rect 222285 241360 223252 241362
rect 222285 241304 222290 241360
rect 222346 241304 223252 241360
rect 222285 241302 223252 241304
rect 222285 241299 222351 241302
rect 223246 241300 223252 241302
rect 223316 241300 223322 241364
rect 226190 241300 226196 241364
rect 226260 241362 226266 241364
rect 284845 241362 284911 241365
rect 226260 241360 284911 241362
rect 226260 241304 284850 241360
rect 284906 241304 284911 241360
rect 226260 241302 284911 241304
rect 226260 241300 226266 241302
rect 284845 241299 284911 241302
rect 220077 241226 220143 241229
rect 227662 241226 227668 241228
rect 220077 241224 227668 241226
rect -960 241090 480 241180
rect 220077 241168 220082 241224
rect 220138 241168 227668 241224
rect 220077 241166 227668 241168
rect 220077 241163 220143 241166
rect 227662 241164 227668 241166
rect 227732 241164 227738 241228
rect 267457 241226 267523 241229
rect 269113 241226 269179 241229
rect 323577 241226 323643 241229
rect 267457 241224 267704 241226
rect 267457 241168 267462 241224
rect 267518 241168 267704 241224
rect 267457 241166 267704 241168
rect 267457 241163 267523 241166
rect 267644 241093 267704 241166
rect 269113 241224 323643 241226
rect 269113 241168 269118 241224
rect 269174 241168 323582 241224
rect 323638 241168 323643 241224
rect 269113 241166 323643 241168
rect 269113 241163 269179 241166
rect 323577 241163 323643 241166
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 213269 241090 213335 241093
rect 215937 241090 216003 241093
rect 223798 241090 223804 241092
rect 213269 241088 215310 241090
rect 213269 241032 213274 241088
rect 213330 241032 215310 241088
rect 213269 241030 215310 241032
rect 213269 241027 213335 241030
rect 215250 240818 215310 241030
rect 215937 241088 223804 241090
rect 215937 241032 215942 241088
rect 215998 241032 223804 241088
rect 215937 241030 223804 241032
rect 215937 241027 216003 241030
rect 223798 241028 223804 241030
rect 223868 241028 223874 241092
rect 226006 241028 226012 241092
rect 226076 241090 226082 241092
rect 234286 241090 234292 241092
rect 226076 241030 234292 241090
rect 226076 241028 226082 241030
rect 234286 241028 234292 241030
rect 234356 241028 234362 241092
rect 267641 241088 267707 241093
rect 267641 241032 267646 241088
rect 267702 241032 267707 241088
rect 267641 241027 267707 241032
rect 268009 241090 268075 241093
rect 325141 241090 325207 241093
rect 268009 241088 325207 241090
rect 268009 241032 268014 241088
rect 268070 241032 325146 241088
rect 325202 241032 325207 241088
rect 268009 241030 325207 241032
rect 268009 241027 268075 241030
rect 325141 241027 325207 241030
rect 217501 240954 217567 240957
rect 232446 240954 232452 240956
rect 217501 240952 232452 240954
rect 217501 240896 217506 240952
rect 217562 240896 232452 240952
rect 217501 240894 232452 240896
rect 217501 240891 217567 240894
rect 232446 240892 232452 240894
rect 232516 240892 232522 240956
rect 265934 240892 265940 240956
rect 266004 240954 266010 240956
rect 327717 240954 327783 240957
rect 266004 240952 327783 240954
rect 266004 240896 327722 240952
rect 327778 240896 327783 240952
rect 266004 240894 327783 240896
rect 266004 240892 266010 240894
rect 327717 240891 327783 240894
rect 226926 240818 226932 240820
rect 215250 240758 226932 240818
rect 226926 240756 226932 240758
rect 226996 240756 227002 240820
rect 228582 240756 228588 240820
rect 228652 240818 228658 240820
rect 231158 240818 231164 240820
rect 228652 240758 231164 240818
rect 228652 240756 228658 240758
rect 231158 240756 231164 240758
rect 231228 240756 231234 240820
rect 268745 240818 268811 240821
rect 327901 240818 327967 240821
rect 268745 240816 327967 240818
rect 268745 240760 268750 240816
rect 268806 240760 327906 240816
rect 327962 240760 327967 240816
rect 268745 240758 327967 240760
rect 268745 240755 268811 240758
rect 327901 240755 327967 240758
rect 217133 240682 217199 240685
rect 217501 240682 217567 240685
rect 217133 240680 217567 240682
rect 217133 240624 217138 240680
rect 217194 240624 217506 240680
rect 217562 240624 217567 240680
rect 217133 240622 217567 240624
rect 217133 240619 217199 240622
rect 217501 240619 217567 240622
rect 218697 240682 218763 240685
rect 229686 240682 229692 240684
rect 218697 240680 229692 240682
rect 218697 240624 218702 240680
rect 218758 240624 229692 240680
rect 218697 240622 229692 240624
rect 218697 240619 218763 240622
rect 229686 240620 229692 240622
rect 229756 240620 229762 240684
rect 248270 240620 248276 240684
rect 248340 240682 248346 240684
rect 295926 240682 295932 240684
rect 248340 240622 295932 240682
rect 248340 240620 248346 240622
rect 295926 240620 295932 240622
rect 295996 240620 296002 240684
rect 213637 240546 213703 240549
rect 220077 240546 220143 240549
rect 213637 240544 220143 240546
rect 213637 240488 213642 240544
rect 213698 240488 220082 240544
rect 220138 240488 220143 240544
rect 213637 240486 220143 240488
rect 213637 240483 213703 240486
rect 220077 240483 220143 240486
rect 220353 240546 220419 240549
rect 227478 240546 227484 240548
rect 220353 240544 227484 240546
rect 220353 240488 220358 240544
rect 220414 240488 227484 240544
rect 220353 240486 227484 240488
rect 220353 240483 220419 240486
rect 227478 240484 227484 240486
rect 227548 240484 227554 240548
rect 217593 240410 217659 240413
rect 217593 240408 223498 240410
rect 217593 240352 217598 240408
rect 217654 240352 223498 240408
rect 217593 240350 223498 240352
rect 217593 240347 217659 240350
rect 215661 240274 215727 240277
rect 215937 240274 216003 240277
rect 215661 240272 216003 240274
rect 215661 240216 215666 240272
rect 215722 240216 215942 240272
rect 215998 240216 216003 240272
rect 215661 240214 216003 240216
rect 215661 240211 215727 240214
rect 215937 240211 216003 240214
rect 217409 240274 217475 240277
rect 220353 240274 220419 240277
rect 217409 240272 220419 240274
rect 217409 240216 217414 240272
rect 217470 240216 220358 240272
rect 220414 240216 220419 240272
rect 217409 240214 220419 240216
rect 217409 240211 217475 240214
rect 220353 240211 220419 240214
rect 220905 240274 220971 240277
rect 222285 240274 222351 240277
rect 220905 240272 222351 240274
rect 220905 240216 220910 240272
rect 220966 240216 222290 240272
rect 222346 240216 222351 240272
rect 220905 240214 222351 240216
rect 223438 240274 223498 240350
rect 223798 240348 223804 240412
rect 223868 240410 223874 240412
rect 223868 240350 226258 240410
rect 223868 240348 223874 240350
rect 226006 240274 226012 240276
rect 223438 240214 226012 240274
rect 220905 240211 220971 240214
rect 222285 240211 222351 240214
rect 226006 240212 226012 240214
rect 226076 240212 226082 240276
rect 222285 240138 222351 240141
rect 223430 240138 223436 240140
rect 222285 240136 223436 240138
rect 222285 240080 222290 240136
rect 222346 240080 223436 240136
rect 222285 240078 223436 240080
rect 222285 240075 222351 240078
rect 223430 240076 223436 240078
rect 223500 240076 223506 240140
rect 215753 240002 215819 240005
rect 216305 240002 216371 240005
rect 215753 240000 216371 240002
rect 215753 239944 215758 240000
rect 215814 239944 216310 240000
rect 216366 239944 216371 240000
rect 215753 239942 216371 239944
rect 215753 239939 215819 239942
rect 216305 239939 216371 239942
rect 223067 239898 223133 239903
rect 222510 239804 222516 239868
rect 222580 239866 222586 239868
rect 223067 239866 223072 239898
rect 222580 239842 223072 239866
rect 223128 239842 223133 239898
rect 224171 239898 224237 239903
rect 224171 239868 224176 239898
rect 224232 239868 224237 239898
rect 222580 239837 223133 239842
rect 222580 239806 223130 239837
rect 222580 239804 222586 239806
rect 224166 239804 224172 239868
rect 224236 239866 224242 239868
rect 224236 239806 224294 239866
rect 224236 239804 224242 239806
rect 224534 239804 224540 239868
rect 224604 239866 224610 239868
rect 225183 239866 225249 239869
rect 226011 239868 226077 239869
rect 226006 239866 226012 239868
rect 224604 239864 225249 239866
rect 224604 239808 225188 239864
rect 225244 239808 225249 239864
rect 224604 239806 225249 239808
rect 225920 239806 226012 239866
rect 224604 239804 224610 239806
rect 225183 239803 225249 239806
rect 226006 239804 226012 239806
rect 226076 239804 226082 239868
rect 226198 239866 226258 240350
rect 230054 240348 230060 240412
rect 230124 240410 230130 240412
rect 230422 240410 230428 240412
rect 230124 240350 230428 240410
rect 230124 240348 230130 240350
rect 230422 240348 230428 240350
rect 230492 240348 230498 240412
rect 230790 240348 230796 240412
rect 230860 240410 230866 240412
rect 238334 240410 238340 240412
rect 230860 240350 238340 240410
rect 230860 240348 230866 240350
rect 238334 240348 238340 240350
rect 238404 240348 238410 240412
rect 230974 240274 230980 240276
rect 228820 240214 230980 240274
rect 228214 240138 228220 240140
rect 227118 240078 228220 240138
rect 226374 239940 226380 240004
rect 226444 240002 226450 240004
rect 227118 240002 227178 240078
rect 228214 240076 228220 240078
rect 228284 240076 228290 240140
rect 226444 239942 227178 240002
rect 226444 239940 226450 239942
rect 227118 239869 227178 239942
rect 227846 239940 227852 240004
rect 227916 240002 227922 240004
rect 227916 239942 228558 240002
rect 227916 239940 227922 239942
rect 227299 239900 227365 239903
rect 227299 239898 227422 239900
rect 226379 239866 226445 239869
rect 226198 239864 226445 239866
rect 226198 239808 226384 239864
rect 226440 239808 226445 239864
rect 226198 239806 226445 239808
rect 226011 239803 226077 239804
rect 226379 239803 226445 239806
rect 226558 239804 226564 239868
rect 226628 239866 226634 239868
rect 226977 239866 227043 239869
rect 226628 239864 227043 239866
rect 226628 239808 226982 239864
rect 227038 239808 227043 239864
rect 226628 239806 227043 239808
rect 226628 239804 226634 239806
rect 226977 239803 227043 239806
rect 227115 239864 227181 239869
rect 227299 239868 227304 239898
rect 227360 239868 227422 239898
rect 227115 239808 227120 239864
rect 227176 239808 227181 239864
rect 227115 239803 227181 239808
rect 227294 239804 227300 239868
rect 227364 239840 227422 239868
rect 227667 239898 227733 239903
rect 227667 239842 227672 239898
rect 227728 239842 227733 239898
rect 228498 239869 228558 239942
rect 228820 239869 228880 240214
rect 230974 240212 230980 240214
rect 231044 240212 231050 240276
rect 268837 240274 268903 240277
rect 265022 240272 268903 240274
rect 265022 240216 268842 240272
rect 268898 240216 268903 240272
rect 265022 240214 268903 240216
rect 231894 240138 231900 240140
rect 230568 240078 231900 240138
rect 230568 240002 230628 240078
rect 231894 240076 231900 240078
rect 231964 240076 231970 240140
rect 237230 240138 237236 240140
rect 237100 240078 237236 240138
rect 229050 239942 230628 240002
rect 229050 239869 229110 239942
rect 231526 239940 231532 240004
rect 231596 240002 231602 240004
rect 231596 239942 232514 240002
rect 231596 239940 231602 239942
rect 227364 239804 227370 239840
rect 227667 239837 227733 239842
rect 227943 239866 228009 239869
rect 228214 239866 228220 239868
rect 227943 239864 228220 239866
rect 227670 239733 227730 239837
rect 227943 239808 227948 239864
rect 228004 239808 228220 239864
rect 227943 239806 228220 239808
rect 227943 239803 228009 239806
rect 228214 239804 228220 239806
rect 228284 239804 228290 239868
rect 228495 239864 228561 239869
rect 228495 239808 228500 239864
rect 228556 239808 228561 239864
rect 228495 239803 228561 239808
rect 228771 239866 228880 239869
rect 228771 239864 228972 239866
rect 228771 239808 228776 239864
rect 228832 239808 228972 239864
rect 228771 239806 228972 239808
rect 228771 239803 228837 239806
rect 228912 239733 228972 239806
rect 229047 239864 229113 239869
rect 229047 239808 229052 239864
rect 229108 239808 229113 239864
rect 229047 239803 229113 239808
rect 229323 239866 229389 239869
rect 230606 239866 230612 239868
rect 229323 239864 230612 239866
rect 229323 239808 229328 239864
rect 229384 239808 230612 239864
rect 229323 239806 230612 239808
rect 229323 239803 229389 239806
rect 230606 239804 230612 239806
rect 230676 239804 230682 239868
rect 231163 239864 231229 239869
rect 231163 239808 231168 239864
rect 231224 239808 231229 239864
rect 231163 239803 231229 239808
rect 231991 239866 232057 239869
rect 232262 239866 232268 239868
rect 231991 239864 232268 239866
rect 231991 239808 231996 239864
rect 232052 239808 232268 239864
rect 231991 239806 232268 239808
rect 231991 239803 232057 239806
rect 232262 239804 232268 239806
rect 232332 239804 232338 239868
rect 232454 239866 232514 239942
rect 232635 239898 232701 239903
rect 232911 239900 232977 239903
rect 232635 239866 232640 239898
rect 232454 239842 232640 239866
rect 232696 239842 232701 239898
rect 232454 239837 232701 239842
rect 232868 239898 232977 239900
rect 232868 239842 232916 239898
rect 232972 239866 232977 239898
rect 233923 239900 233989 239903
rect 236959 239900 237025 239903
rect 237100 239900 237160 240078
rect 237230 240076 237236 240078
rect 237300 240076 237306 240140
rect 265022 240138 265082 240214
rect 268837 240211 268903 240214
rect 268653 240138 268719 240141
rect 262998 240078 265082 240138
rect 265206 240136 268719 240138
rect 265206 240080 268658 240136
rect 268714 240080 268719 240136
rect 265206 240078 268719 240080
rect 237414 239940 237420 240004
rect 237484 240002 237490 240004
rect 238150 240002 238156 240004
rect 237484 239942 238156 240002
rect 237484 239940 237490 239942
rect 238150 239940 238156 239942
rect 238220 240002 238226 240004
rect 238220 239942 238770 240002
rect 238220 239940 238226 239942
rect 233923 239898 234046 239900
rect 233647 239866 233713 239869
rect 233923 239868 233928 239898
rect 233984 239868 234046 239898
rect 236959 239898 237160 239900
rect 234291 239868 234357 239869
rect 234659 239868 234725 239869
rect 232972 239842 233388 239866
rect 232454 239806 232698 239837
rect 232868 239806 233388 239842
rect 231166 239733 231226 239803
rect 222745 239732 222811 239733
rect 223113 239732 223179 239733
rect 222694 239668 222700 239732
rect 222764 239730 222811 239732
rect 223062 239730 223068 239732
rect 222764 239728 222856 239730
rect 222806 239672 222856 239728
rect 222764 239670 222856 239672
rect 223022 239670 223068 239730
rect 223132 239728 223179 239732
rect 223174 239672 223179 239728
rect 222764 239668 222811 239670
rect 223062 239668 223068 239670
rect 223132 239668 223179 239672
rect 223246 239668 223252 239732
rect 223316 239730 223322 239732
rect 223389 239730 223455 239733
rect 223849 239732 223915 239733
rect 223316 239728 223455 239730
rect 223316 239672 223394 239728
rect 223450 239672 223455 239728
rect 223316 239670 223455 239672
rect 223316 239668 223322 239670
rect 222745 239667 222811 239668
rect 223113 239667 223179 239668
rect 223389 239667 223455 239670
rect 223798 239668 223804 239732
rect 223868 239730 223915 239732
rect 224309 239730 224375 239733
rect 224718 239730 224724 239732
rect 223868 239728 223960 239730
rect 223910 239672 223960 239728
rect 223868 239670 223960 239672
rect 224309 239728 224724 239730
rect 224309 239672 224314 239728
rect 224370 239672 224724 239728
rect 224309 239670 224724 239672
rect 223868 239668 223915 239670
rect 223806 239667 223915 239668
rect 224309 239667 224375 239670
rect 224718 239668 224724 239670
rect 224788 239668 224794 239732
rect 224902 239668 224908 239732
rect 224972 239730 224978 239732
rect 226057 239730 226123 239733
rect 226701 239732 226767 239733
rect 226885 239732 226951 239733
rect 226701 239730 226748 239732
rect 224972 239728 226123 239730
rect 224972 239672 226062 239728
rect 226118 239672 226123 239728
rect 224972 239670 226123 239672
rect 226656 239728 226748 239730
rect 226656 239672 226706 239728
rect 226656 239670 226748 239672
rect 224972 239668 224978 239670
rect 226057 239667 226123 239670
rect 226701 239668 226748 239670
rect 226812 239668 226818 239732
rect 226885 239728 226932 239732
rect 226996 239730 227002 239732
rect 227621 239730 227730 239733
rect 228030 239730 228036 239732
rect 226885 239672 226890 239728
rect 226885 239668 226932 239672
rect 226996 239670 227042 239730
rect 227540 239728 228036 239730
rect 227540 239672 227626 239728
rect 227682 239672 228036 239728
rect 227540 239670 228036 239672
rect 226996 239668 227002 239670
rect 226701 239667 226767 239668
rect 226885 239667 226951 239668
rect 227621 239667 227687 239670
rect 228030 239668 228036 239670
rect 228100 239668 228106 239732
rect 228909 239728 228975 239733
rect 228909 239672 228914 239728
rect 228970 239672 228975 239728
rect 228909 239667 228975 239672
rect 229870 239668 229876 239732
rect 229940 239730 229946 239732
rect 230197 239730 230263 239733
rect 229940 239728 230263 239730
rect 229940 239672 230202 239728
rect 230258 239672 230263 239728
rect 229940 239670 230263 239672
rect 229940 239668 229946 239670
rect 230197 239667 230263 239670
rect 230381 239732 230447 239733
rect 230381 239728 230428 239732
rect 230492 239730 230498 239732
rect 230749 239730 230815 239733
rect 230974 239730 230980 239732
rect 230381 239672 230386 239728
rect 230381 239668 230428 239672
rect 230492 239670 230538 239730
rect 230749 239728 230980 239730
rect 230749 239672 230754 239728
rect 230810 239672 230980 239728
rect 230749 239670 230980 239672
rect 230492 239668 230498 239670
rect 230381 239667 230447 239668
rect 230749 239667 230815 239670
rect 230974 239668 230980 239670
rect 231044 239668 231050 239732
rect 231166 239730 231275 239733
rect 232078 239730 232084 239732
rect 231166 239728 232084 239730
rect 231166 239672 231214 239728
rect 231270 239672 232084 239728
rect 231166 239670 232084 239672
rect 231209 239667 231275 239670
rect 232078 239668 232084 239670
rect 232148 239668 232154 239732
rect 232446 239668 232452 239732
rect 232516 239730 232522 239732
rect 233141 239730 233207 239733
rect 232516 239728 233207 239730
rect 232516 239672 233146 239728
rect 233202 239672 233207 239728
rect 232516 239670 233207 239672
rect 232516 239668 232522 239670
rect 233141 239667 233207 239670
rect 220721 239594 220787 239597
rect 223573 239594 223639 239597
rect 220721 239592 223639 239594
rect 220721 239536 220726 239592
rect 220782 239536 223578 239592
rect 223634 239536 223639 239592
rect 220721 239534 223639 239536
rect 220721 239531 220787 239534
rect 223573 239531 223639 239534
rect 220670 239396 220676 239460
rect 220740 239458 220746 239460
rect 222607 239458 222673 239461
rect 222929 239458 222995 239461
rect 220740 239456 222995 239458
rect 220740 239400 222612 239456
rect 222668 239400 222934 239456
rect 222990 239400 222995 239456
rect 220740 239398 222995 239400
rect 220740 239396 220746 239398
rect 222607 239395 222673 239398
rect 222929 239395 222995 239398
rect 223297 239458 223363 239461
rect 223806 239458 223866 239667
rect 223941 239596 224007 239597
rect 223941 239592 223988 239596
rect 224052 239594 224058 239596
rect 224585 239594 224651 239597
rect 224052 239592 224651 239594
rect 223941 239536 223946 239592
rect 224052 239536 224590 239592
rect 224646 239536 224651 239592
rect 223941 239532 223988 239536
rect 224052 239534 224651 239536
rect 224052 239532 224058 239534
rect 223941 239531 224007 239532
rect 224585 239531 224651 239534
rect 225321 239594 225387 239597
rect 226190 239594 226196 239596
rect 225321 239592 226196 239594
rect 225321 239536 225326 239592
rect 225382 239536 226196 239592
rect 225321 239534 226196 239536
rect 225321 239531 225387 239534
rect 226190 239532 226196 239534
rect 226260 239532 226266 239596
rect 227110 239532 227116 239596
rect 227180 239594 227186 239596
rect 227253 239594 227319 239597
rect 227180 239592 227319 239594
rect 227180 239536 227258 239592
rect 227314 239536 227319 239592
rect 227180 239534 227319 239536
rect 227180 239532 227186 239534
rect 227253 239531 227319 239534
rect 227478 239532 227484 239596
rect 227548 239594 227554 239596
rect 227713 239594 227779 239597
rect 227548 239592 227779 239594
rect 227548 239536 227718 239592
rect 227774 239536 227779 239592
rect 227548 239534 227779 239536
rect 227548 239532 227554 239534
rect 227713 239531 227779 239534
rect 230381 239594 230447 239597
rect 230790 239594 230796 239596
rect 230381 239592 230796 239594
rect 230381 239536 230386 239592
rect 230442 239536 230796 239592
rect 230381 239534 230796 239536
rect 230381 239531 230447 239534
rect 230790 239532 230796 239534
rect 230860 239532 230866 239596
rect 231301 239594 231367 239597
rect 231710 239594 231716 239596
rect 231301 239592 231716 239594
rect 231301 239536 231306 239592
rect 231362 239536 231716 239592
rect 231301 239534 231716 239536
rect 231301 239531 231367 239534
rect 231710 239532 231716 239534
rect 231780 239532 231786 239596
rect 231894 239532 231900 239596
rect 231964 239594 231970 239596
rect 232589 239594 232655 239597
rect 231964 239592 232655 239594
rect 231964 239536 232594 239592
rect 232650 239536 232655 239592
rect 231964 239534 232655 239536
rect 231964 239532 231970 239534
rect 232589 239531 232655 239534
rect 232865 239594 232931 239597
rect 233328 239594 233388 239806
rect 233647 239864 233756 239866
rect 233647 239808 233652 239864
rect 233708 239808 233756 239864
rect 233647 239803 233756 239808
rect 233918 239804 233924 239868
rect 233988 239840 234046 239868
rect 234286 239866 234292 239868
rect 233988 239804 233994 239840
rect 234200 239806 234292 239866
rect 234286 239804 234292 239806
rect 234356 239804 234362 239868
rect 234654 239866 234660 239868
rect 234568 239806 234660 239866
rect 234654 239804 234660 239806
rect 234724 239804 234730 239868
rect 235206 239804 235212 239868
rect 235276 239866 235282 239868
rect 235947 239866 236013 239869
rect 235276 239864 236013 239866
rect 235276 239808 235952 239864
rect 236008 239808 236013 239864
rect 235276 239806 236013 239808
rect 235276 239804 235282 239806
rect 234291 239803 234357 239804
rect 234659 239803 234725 239804
rect 235947 239803 236013 239806
rect 236126 239804 236132 239868
rect 236196 239866 236202 239868
rect 236591 239866 236657 239869
rect 236196 239864 236657 239866
rect 236196 239808 236596 239864
rect 236652 239808 236657 239864
rect 236959 239842 236964 239898
rect 237020 239842 237160 239898
rect 238710 239869 238770 239942
rect 243118 239940 243124 240004
rect 243188 240002 243194 240004
rect 259310 240002 259316 240004
rect 243188 239940 243232 240002
rect 240639 239900 240705 239903
rect 240639 239898 240748 239900
rect 236959 239840 237160 239842
rect 238155 239866 238221 239869
rect 238518 239866 238524 239868
rect 238155 239864 238524 239866
rect 236959 239837 237025 239840
rect 236196 239806 236657 239808
rect 236196 239804 236202 239806
rect 236591 239803 236657 239806
rect 238155 239808 238160 239864
rect 238216 239808 238524 239864
rect 238155 239806 238524 239808
rect 238155 239803 238221 239806
rect 238518 239804 238524 239806
rect 238588 239804 238594 239868
rect 238707 239864 238773 239869
rect 238707 239808 238712 239864
rect 238768 239808 238773 239864
rect 238707 239803 238773 239808
rect 239070 239804 239076 239868
rect 239140 239866 239146 239868
rect 239259 239866 239325 239869
rect 239140 239864 239325 239866
rect 239140 239808 239264 239864
rect 239320 239808 239325 239864
rect 240639 239842 240644 239898
rect 240700 239866 240748 239898
rect 240910 239866 240916 239868
rect 240700 239842 240916 239866
rect 240639 239837 240916 239842
rect 239140 239806 239325 239808
rect 240688 239806 240916 239837
rect 239140 239804 239146 239806
rect 239259 239803 239325 239806
rect 240910 239804 240916 239806
rect 240980 239804 240986 239868
rect 241743 239866 241809 239869
rect 242014 239866 242020 239868
rect 241743 239864 242020 239866
rect 241743 239808 241748 239864
rect 241804 239808 242020 239864
rect 241743 239806 242020 239808
rect 241743 239803 241809 239806
rect 242014 239804 242020 239806
rect 242084 239804 242090 239868
rect 242341 239866 242407 239869
rect 242479 239866 242545 239869
rect 242755 239868 242821 239869
rect 242750 239866 242756 239868
rect 242341 239864 242545 239866
rect 242341 239808 242346 239864
rect 242402 239808 242484 239864
rect 242540 239808 242545 239864
rect 242341 239806 242545 239808
rect 242664 239806 242756 239866
rect 242341 239803 242407 239806
rect 242479 239803 242545 239806
rect 242750 239804 242756 239806
rect 242820 239804 242826 239868
rect 243031 239866 243097 239869
rect 243172 239866 243232 239940
rect 258582 239942 259316 240002
rect 257475 239898 257541 239903
rect 257935 239900 258001 239903
rect 246205 239868 246271 239869
rect 246205 239866 246252 239868
rect 243031 239864 243232 239866
rect 243031 239808 243036 239864
rect 243092 239808 243232 239864
rect 243031 239806 243232 239808
rect 246124 239864 246252 239866
rect 246316 239866 246322 239868
rect 246798 239866 246804 239868
rect 246124 239808 246210 239864
rect 246124 239806 246252 239808
rect 242755 239803 242821 239804
rect 243031 239803 243097 239806
rect 246205 239804 246252 239806
rect 246316 239806 246804 239866
rect 246316 239804 246322 239806
rect 246798 239804 246804 239806
rect 246868 239804 246874 239868
rect 247534 239804 247540 239868
rect 247604 239866 247610 239868
rect 247815 239866 247881 239869
rect 248086 239866 248092 239868
rect 247604 239864 248092 239866
rect 247604 239808 247820 239864
rect 247876 239808 248092 239864
rect 247604 239806 248092 239808
rect 247604 239804 247610 239806
rect 246205 239803 246271 239804
rect 247815 239803 247881 239806
rect 248086 239804 248092 239806
rect 248156 239804 248162 239868
rect 249006 239804 249012 239868
rect 249076 239866 249082 239868
rect 249747 239866 249813 239869
rect 249076 239864 249813 239866
rect 249076 239808 249752 239864
rect 249808 239808 249813 239864
rect 249076 239806 249813 239808
rect 249076 239804 249082 239806
rect 249747 239803 249813 239806
rect 250294 239804 250300 239868
rect 250364 239866 250370 239868
rect 250851 239866 250917 239869
rect 251030 239866 251036 239868
rect 250364 239864 251036 239866
rect 250364 239808 250856 239864
rect 250912 239808 251036 239864
rect 250364 239806 251036 239808
rect 250364 239804 250370 239806
rect 250851 239803 250917 239806
rect 251030 239804 251036 239806
rect 251100 239804 251106 239868
rect 251403 239864 251469 239869
rect 251403 239808 251408 239864
rect 251464 239808 251469 239864
rect 251403 239803 251469 239808
rect 251582 239804 251588 239868
rect 251652 239866 251658 239868
rect 251955 239866 252021 239869
rect 251652 239864 252021 239866
rect 251652 239808 251960 239864
rect 252016 239808 252021 239864
rect 251652 239806 252021 239808
rect 251652 239804 251658 239806
rect 251955 239803 252021 239806
rect 252870 239804 252876 239868
rect 252940 239866 252946 239868
rect 253335 239866 253401 239869
rect 252940 239864 254042 239866
rect 252940 239808 253340 239864
rect 253396 239808 254042 239864
rect 252940 239806 254042 239808
rect 252940 239804 252946 239806
rect 253335 239803 253401 239806
rect 233696 239732 233756 239803
rect 233696 239670 233740 239732
rect 233734 239668 233740 239670
rect 233804 239668 233810 239732
rect 235390 239668 235396 239732
rect 235460 239730 235466 239732
rect 235717 239730 235783 239733
rect 235460 239728 235783 239730
rect 235460 239672 235722 239728
rect 235778 239672 235783 239728
rect 235460 239670 235783 239672
rect 235460 239668 235466 239670
rect 235717 239667 235783 239670
rect 235993 239730 236059 239733
rect 237281 239730 237347 239733
rect 235993 239728 237347 239730
rect 235993 239672 235998 239728
rect 236054 239672 237286 239728
rect 237342 239672 237347 239728
rect 235993 239670 237347 239672
rect 235993 239667 236059 239670
rect 237281 239667 237347 239670
rect 238385 239730 238451 239733
rect 238385 239728 238586 239730
rect 238385 239672 238390 239728
rect 238446 239672 238586 239728
rect 238385 239670 238586 239672
rect 238385 239667 238451 239670
rect 232865 239592 233388 239594
rect 232865 239536 232870 239592
rect 232926 239536 233388 239592
rect 232865 239534 233388 239536
rect 232865 239531 232931 239534
rect 233550 239532 233556 239596
rect 233620 239594 233626 239596
rect 233693 239594 233759 239597
rect 234470 239594 234476 239596
rect 233620 239592 234476 239594
rect 233620 239536 233698 239592
rect 233754 239536 234476 239592
rect 233620 239534 234476 239536
rect 233620 239532 233626 239534
rect 233693 239531 233759 239534
rect 234470 239532 234476 239534
rect 234540 239532 234546 239596
rect 234613 239594 234679 239597
rect 236453 239594 236519 239597
rect 234613 239592 236519 239594
rect 234613 239536 234618 239592
rect 234674 239536 236458 239592
rect 236514 239536 236519 239592
rect 234613 239534 236519 239536
rect 234613 239531 234679 239534
rect 236453 239531 236519 239534
rect 238526 239461 238586 239670
rect 238886 239668 238892 239732
rect 238956 239730 238962 239732
rect 239213 239730 239279 239733
rect 238956 239728 239279 239730
rect 238956 239672 239218 239728
rect 239274 239672 239279 239728
rect 238956 239670 239279 239672
rect 238956 239668 238962 239670
rect 239213 239667 239279 239670
rect 242382 239668 242388 239732
rect 242452 239730 242458 239732
rect 242525 239730 242591 239733
rect 242452 239728 242591 239730
rect 242452 239672 242530 239728
rect 242586 239672 242591 239728
rect 242452 239670 242591 239672
rect 242452 239668 242458 239670
rect 242525 239667 242591 239670
rect 244958 239668 244964 239732
rect 245028 239730 245034 239732
rect 245193 239730 245259 239733
rect 245028 239728 245259 239730
rect 245028 239672 245198 239728
rect 245254 239672 245259 239728
rect 245028 239670 245259 239672
rect 245028 239668 245034 239670
rect 245193 239667 245259 239670
rect 246062 239668 246068 239732
rect 246132 239730 246138 239732
rect 246757 239730 246823 239733
rect 247861 239732 247927 239733
rect 247861 239730 247908 239732
rect 246132 239728 246823 239730
rect 246132 239672 246762 239728
rect 246818 239672 246823 239728
rect 246132 239670 246823 239672
rect 247816 239728 247908 239730
rect 247816 239672 247866 239728
rect 247816 239670 247908 239672
rect 246132 239668 246138 239670
rect 246757 239667 246823 239670
rect 247861 239668 247908 239670
rect 247972 239668 247978 239732
rect 248045 239730 248111 239733
rect 248270 239730 248276 239732
rect 248045 239728 248276 239730
rect 248045 239672 248050 239728
rect 248106 239672 248276 239728
rect 248045 239670 248276 239672
rect 247861 239667 247927 239668
rect 248045 239667 248154 239670
rect 248270 239668 248276 239670
rect 248340 239668 248346 239732
rect 249241 239730 249307 239733
rect 249558 239730 249564 239732
rect 249241 239728 249564 239730
rect 249241 239672 249246 239728
rect 249302 239672 249564 239728
rect 249241 239670 249564 239672
rect 249241 239667 249307 239670
rect 249558 239668 249564 239670
rect 249628 239668 249634 239732
rect 250345 239730 250411 239733
rect 250662 239730 250668 239732
rect 250345 239728 250668 239730
rect 250345 239672 250350 239728
rect 250406 239672 250668 239728
rect 250345 239670 250668 239672
rect 250345 239667 250411 239670
rect 250662 239668 250668 239670
rect 250732 239668 250738 239732
rect 251406 239730 251466 239803
rect 251950 239730 251956 239732
rect 251406 239670 251956 239730
rect 251950 239668 251956 239670
rect 252020 239668 252026 239732
rect 252134 239668 252140 239732
rect 252204 239730 252210 239732
rect 252645 239730 252711 239733
rect 253105 239730 253171 239733
rect 252204 239728 252711 239730
rect 252204 239672 252650 239728
rect 252706 239672 252711 239728
rect 252204 239670 252711 239672
rect 252204 239668 252210 239670
rect 252645 239667 252711 239670
rect 252878 239728 253171 239730
rect 252878 239672 253110 239728
rect 253166 239672 253171 239728
rect 252878 239670 253171 239672
rect 238702 239532 238708 239596
rect 238772 239594 238778 239596
rect 239438 239594 239444 239596
rect 238772 239534 239444 239594
rect 238772 239532 238778 239534
rect 239438 239532 239444 239534
rect 239508 239594 239514 239596
rect 240041 239594 240107 239597
rect 241329 239596 241395 239597
rect 239508 239592 240107 239594
rect 239508 239536 240046 239592
rect 240102 239536 240107 239592
rect 239508 239534 240107 239536
rect 239508 239532 239514 239534
rect 240041 239531 240107 239534
rect 241278 239532 241284 239596
rect 241348 239594 241395 239596
rect 241348 239592 241440 239594
rect 241390 239536 241440 239592
rect 241348 239534 241440 239536
rect 241348 239532 241395 239534
rect 242198 239532 242204 239596
rect 242268 239594 242274 239596
rect 242893 239594 242959 239597
rect 242268 239592 242959 239594
rect 242268 239536 242898 239592
rect 242954 239536 242959 239592
rect 242268 239534 242959 239536
rect 242268 239532 242274 239534
rect 241329 239531 241395 239532
rect 242893 239531 242959 239534
rect 243169 239594 243235 239597
rect 243302 239594 243308 239596
rect 243169 239592 243308 239594
rect 243169 239536 243174 239592
rect 243230 239536 243308 239592
rect 243169 239534 243308 239536
rect 243169 239531 243235 239534
rect 243302 239532 243308 239534
rect 243372 239532 243378 239596
rect 245193 239594 245259 239597
rect 245510 239594 245516 239596
rect 245193 239592 245516 239594
rect 245193 239536 245198 239592
rect 245254 239536 245516 239592
rect 245193 239534 245516 239536
rect 245193 239531 245259 239534
rect 245510 239532 245516 239534
rect 245580 239532 245586 239596
rect 246021 239594 246087 239597
rect 246614 239594 246620 239596
rect 246021 239592 246620 239594
rect 246021 239536 246026 239592
rect 246082 239536 246620 239592
rect 246021 239534 246620 239536
rect 246021 239531 246087 239534
rect 246614 239532 246620 239534
rect 246684 239532 246690 239596
rect 247718 239532 247724 239596
rect 247788 239594 247794 239596
rect 248094 239594 248154 239667
rect 252878 239597 252938 239670
rect 253105 239667 253171 239670
rect 253238 239668 253244 239732
rect 253308 239730 253314 239732
rect 253749 239730 253815 239733
rect 253308 239728 253815 239730
rect 253308 239672 253754 239728
rect 253810 239672 253815 239728
rect 253308 239670 253815 239672
rect 253308 239668 253314 239670
rect 253749 239667 253815 239670
rect 247788 239534 248154 239594
rect 248873 239594 248939 239597
rect 249374 239594 249380 239596
rect 248873 239592 249380 239594
rect 248873 239536 248878 239592
rect 248934 239536 249380 239592
rect 248873 239534 249380 239536
rect 247788 239532 247794 239534
rect 248873 239531 248939 239534
rect 249374 239532 249380 239534
rect 249444 239594 249450 239596
rect 249517 239594 249583 239597
rect 249444 239592 249583 239594
rect 249444 239536 249522 239592
rect 249578 239536 249583 239592
rect 249444 239534 249583 239536
rect 249444 239532 249450 239534
rect 249517 239531 249583 239534
rect 251633 239594 251699 239597
rect 251766 239594 251772 239596
rect 251633 239592 251772 239594
rect 251633 239536 251638 239592
rect 251694 239536 251772 239592
rect 251633 239534 251772 239536
rect 251633 239531 251699 239534
rect 251766 239532 251772 239534
rect 251836 239594 251842 239596
rect 252461 239594 252527 239597
rect 251836 239592 252527 239594
rect 251836 239536 252466 239592
rect 252522 239536 252527 239592
rect 251836 239534 252527 239536
rect 252878 239592 252987 239597
rect 252878 239536 252926 239592
rect 252982 239536 252987 239592
rect 252878 239534 252987 239536
rect 251836 239532 251842 239534
rect 252461 239531 252527 239534
rect 252921 239531 252987 239534
rect 253054 239532 253060 239596
rect 253124 239594 253130 239596
rect 253381 239594 253447 239597
rect 253124 239592 253447 239594
rect 253124 239536 253386 239592
rect 253442 239536 253447 239592
rect 253124 239534 253447 239536
rect 253124 239532 253130 239534
rect 253381 239531 253447 239534
rect 253749 239594 253815 239597
rect 253982 239594 254042 239806
rect 254163 239864 254229 239869
rect 254163 239808 254168 239864
rect 254224 239808 254229 239864
rect 254163 239803 254229 239808
rect 254531 239864 254597 239869
rect 255175 239866 255241 239869
rect 254531 239808 254536 239864
rect 254592 239808 254597 239864
rect 254531 239803 254597 239808
rect 255040 239864 255241 239866
rect 255040 239808 255180 239864
rect 255236 239808 255241 239864
rect 255040 239806 255241 239808
rect 253749 239592 254042 239594
rect 253749 239536 253754 239592
rect 253810 239536 254042 239592
rect 253749 239534 254042 239536
rect 253749 239531 253815 239534
rect 223297 239456 223866 239458
rect 223297 239400 223302 239456
rect 223358 239400 223866 239456
rect 223297 239398 223866 239400
rect 223297 239395 223363 239398
rect 227662 239396 227668 239460
rect 227732 239458 227738 239460
rect 228173 239458 228239 239461
rect 227732 239456 228239 239458
rect 227732 239400 228178 239456
rect 228234 239400 228239 239456
rect 227732 239398 228239 239400
rect 227732 239396 227738 239398
rect 228173 239395 228239 239398
rect 228357 239458 228423 239461
rect 228582 239458 228588 239460
rect 228357 239456 228588 239458
rect 228357 239400 228362 239456
rect 228418 239400 228588 239456
rect 228357 239398 228588 239400
rect 228357 239395 228423 239398
rect 228582 239396 228588 239398
rect 228652 239396 228658 239460
rect 229461 239458 229527 239461
rect 236126 239458 236132 239460
rect 229461 239456 236132 239458
rect 229461 239400 229466 239456
rect 229522 239400 236132 239456
rect 229461 239398 236132 239400
rect 229461 239395 229527 239398
rect 236126 239396 236132 239398
rect 236196 239396 236202 239460
rect 238526 239456 238635 239461
rect 238526 239400 238574 239456
rect 238630 239400 238635 239456
rect 238526 239398 238635 239400
rect 238569 239395 238635 239398
rect 243353 239458 243419 239461
rect 243486 239458 243492 239460
rect 243353 239456 243492 239458
rect 243353 239400 243358 239456
rect 243414 239400 243492 239456
rect 243353 239398 243492 239400
rect 243353 239395 243419 239398
rect 243486 239396 243492 239398
rect 243556 239396 243562 239460
rect 247350 239396 247356 239460
rect 247420 239458 247426 239460
rect 248045 239458 248111 239461
rect 247420 239456 248111 239458
rect 247420 239400 248050 239456
rect 248106 239400 248111 239456
rect 247420 239398 248111 239400
rect 247420 239396 247426 239398
rect 248045 239395 248111 239398
rect 249190 239396 249196 239460
rect 249260 239458 249266 239460
rect 249333 239458 249399 239461
rect 249260 239456 249399 239458
rect 249260 239400 249338 239456
rect 249394 239400 249399 239456
rect 249260 239398 249399 239400
rect 249260 239396 249266 239398
rect 249333 239395 249399 239398
rect 250069 239458 250135 239461
rect 250846 239458 250852 239460
rect 250069 239456 250852 239458
rect 250069 239400 250074 239456
rect 250130 239400 250852 239456
rect 250069 239398 250852 239400
rect 250069 239395 250135 239398
rect 250846 239396 250852 239398
rect 250916 239396 250922 239460
rect 254166 239458 254226 239803
rect 254534 239597 254594 239803
rect 255040 239730 255100 239806
rect 255175 239803 255241 239806
rect 255630 239804 255636 239868
rect 255700 239866 255706 239868
rect 255700 239806 256112 239866
rect 255700 239804 255706 239806
rect 255221 239730 255287 239733
rect 255040 239728 255287 239730
rect 255040 239672 255226 239728
rect 255282 239672 255287 239728
rect 255040 239670 255287 239672
rect 256052 239730 256112 239806
rect 256182 239804 256188 239868
rect 256252 239866 256258 239868
rect 256647 239866 256713 239869
rect 256252 239864 256713 239866
rect 256252 239808 256652 239864
rect 256708 239808 256713 239864
rect 256252 239806 256713 239808
rect 256252 239804 256258 239806
rect 256647 239803 256713 239806
rect 256918 239804 256924 239868
rect 256988 239866 256994 239868
rect 257475 239866 257480 239898
rect 256988 239842 257480 239866
rect 257536 239842 257541 239898
rect 256988 239837 257541 239842
rect 257892 239898 258001 239900
rect 257892 239842 257940 239898
rect 257996 239842 258001 239898
rect 257892 239837 258001 239842
rect 258211 239898 258277 239903
rect 258211 239842 258216 239898
rect 258272 239842 258277 239898
rect 258582 239869 258642 239942
rect 259310 239940 259316 239942
rect 259380 239940 259386 240004
rect 262998 239903 263058 240078
rect 263910 239940 263916 240004
rect 263980 240002 263986 240004
rect 263980 239942 264944 240002
rect 263980 239940 263986 239942
rect 264884 239903 264944 239942
rect 261891 239898 261957 239903
rect 258211 239837 258277 239842
rect 258579 239864 258645 239869
rect 256988 239806 257538 239837
rect 256988 239804 256994 239806
rect 256509 239730 256575 239733
rect 256052 239728 256575 239730
rect 256052 239672 256514 239728
rect 256570 239672 256575 239728
rect 256052 239670 256575 239672
rect 255221 239667 255287 239670
rect 256509 239667 256575 239670
rect 256734 239668 256740 239732
rect 256804 239730 256810 239732
rect 256969 239730 257035 239733
rect 256804 239728 257035 239730
rect 256804 239672 256974 239728
rect 257030 239672 257035 239728
rect 256804 239670 257035 239672
rect 257892 239730 257952 239837
rect 258214 239733 258274 239837
rect 258579 239808 258584 239864
rect 258640 239808 258645 239864
rect 258579 239803 258645 239808
rect 258942 239804 258948 239868
rect 259012 239866 259018 239868
rect 259131 239866 259197 239869
rect 259012 239864 259197 239866
rect 259012 239808 259136 239864
rect 259192 239808 259197 239864
rect 259012 239806 259197 239808
rect 259012 239804 259018 239806
rect 259131 239803 259197 239806
rect 259591 239866 259657 239869
rect 259591 239864 259700 239866
rect 259591 239808 259596 239864
rect 259652 239808 259700 239864
rect 259591 239803 259700 239808
rect 260419 239864 260485 239869
rect 260419 239808 260424 239864
rect 260480 239808 260485 239864
rect 260419 239803 260485 239808
rect 260782 239804 260788 239868
rect 260852 239866 260858 239868
rect 261891 239866 261896 239898
rect 260852 239842 261896 239866
rect 261952 239842 261957 239898
rect 262075 239898 262141 239903
rect 262075 239868 262080 239898
rect 262136 239868 262141 239898
rect 262995 239898 263061 239903
rect 260852 239837 261957 239842
rect 260852 239806 261954 239837
rect 260852 239804 260858 239806
rect 262070 239804 262076 239868
rect 262140 239866 262146 239868
rect 262581 239866 262647 239869
rect 262140 239806 262198 239866
rect 262581 239864 262874 239866
rect 262581 239808 262586 239864
rect 262642 239808 262874 239864
rect 262995 239842 263000 239898
rect 263056 239842 263061 239898
rect 264884 239898 264993 239903
rect 262995 239837 263061 239842
rect 263823 239866 263889 239869
rect 264278 239866 264284 239868
rect 263823 239864 264284 239866
rect 262581 239806 262874 239808
rect 262140 239804 262146 239806
rect 262581 239803 262647 239806
rect 259640 239733 259700 239803
rect 258073 239730 258139 239733
rect 257892 239728 258139 239730
rect 257892 239672 258078 239728
rect 258134 239672 258139 239728
rect 257892 239670 258139 239672
rect 258214 239728 258323 239733
rect 258214 239672 258262 239728
rect 258318 239672 258323 239728
rect 258214 239670 258323 239672
rect 256804 239668 256810 239670
rect 256969 239667 257035 239670
rect 258073 239667 258139 239670
rect 258257 239667 258323 239670
rect 258441 239730 258507 239733
rect 258441 239728 258642 239730
rect 258441 239672 258446 239728
rect 258502 239672 258642 239728
rect 258441 239670 258642 239672
rect 258441 239667 258507 239670
rect 254534 239592 254643 239597
rect 254534 239536 254582 239592
rect 254638 239536 254643 239592
rect 254534 239534 254643 239536
rect 254577 239531 254643 239534
rect 254710 239532 254716 239596
rect 254780 239594 254786 239596
rect 255037 239594 255103 239597
rect 254780 239592 255103 239594
rect 254780 239536 255042 239592
rect 255098 239536 255103 239592
rect 254780 239534 255103 239536
rect 254780 239532 254786 239534
rect 255037 239531 255103 239534
rect 255446 239532 255452 239596
rect 255516 239594 255522 239596
rect 255589 239594 255655 239597
rect 256325 239596 256391 239597
rect 255516 239592 255655 239594
rect 255516 239536 255594 239592
rect 255650 239536 255655 239592
rect 255516 239534 255655 239536
rect 255516 239532 255522 239534
rect 255589 239531 255655 239534
rect 255814 239532 255820 239596
rect 255884 239594 255890 239596
rect 256325 239594 256372 239596
rect 255884 239592 256372 239594
rect 256436 239594 256442 239596
rect 255884 239536 256330 239592
rect 255884 239534 256372 239536
rect 255884 239532 255890 239534
rect 256325 239532 256372 239534
rect 256436 239534 256518 239594
rect 256436 239532 256442 239534
rect 257102 239532 257108 239596
rect 257172 239594 257178 239596
rect 257889 239594 257955 239597
rect 257172 239592 257955 239594
rect 257172 239536 257894 239592
rect 257950 239536 257955 239592
rect 257172 239534 257955 239536
rect 257172 239532 257178 239534
rect 256325 239531 256391 239532
rect 257889 239531 257955 239534
rect 255037 239458 255103 239461
rect 254166 239456 255103 239458
rect 254166 239400 255042 239456
rect 255098 239400 255103 239456
rect 254166 239398 255103 239400
rect 255037 239395 255103 239398
rect 256141 239458 256207 239461
rect 256734 239458 256740 239460
rect 256141 239456 256740 239458
rect 256141 239400 256146 239456
rect 256202 239400 256740 239456
rect 256141 239398 256740 239400
rect 256141 239395 256207 239398
rect 256734 239396 256740 239398
rect 256804 239396 256810 239460
rect 258582 239458 258642 239670
rect 259637 239728 259703 239733
rect 259637 239672 259642 239728
rect 259698 239672 259703 239728
rect 259637 239667 259703 239672
rect 260422 239730 260482 239803
rect 262489 239730 262555 239733
rect 262622 239730 262628 239732
rect 260422 239670 262092 239730
rect 258758 239532 258764 239596
rect 258828 239594 258834 239596
rect 259085 239594 259151 239597
rect 258828 239592 259151 239594
rect 258828 239536 259090 239592
rect 259146 239536 259151 239592
rect 258828 239534 259151 239536
rect 258828 239532 258834 239534
rect 259085 239531 259151 239534
rect 260097 239594 260163 239597
rect 260925 239596 260991 239597
rect 260598 239594 260604 239596
rect 260097 239592 260604 239594
rect 260097 239536 260102 239592
rect 260158 239536 260604 239592
rect 260097 239534 260604 239536
rect 260097 239531 260163 239534
rect 260598 239532 260604 239534
rect 260668 239532 260674 239596
rect 260925 239594 260972 239596
rect 260880 239592 260972 239594
rect 260880 239536 260930 239592
rect 260880 239534 260972 239536
rect 260925 239532 260972 239534
rect 261036 239532 261042 239596
rect 260925 239531 260991 239532
rect 259177 239460 259243 239461
rect 258582 239398 259056 239458
rect 222837 239322 222903 239325
rect 237925 239322 237991 239325
rect 222837 239320 237991 239322
rect 222837 239264 222842 239320
rect 222898 239264 237930 239320
rect 237986 239264 237991 239320
rect 222837 239262 237991 239264
rect 222837 239259 222903 239262
rect 237925 239259 237991 239262
rect 238334 239260 238340 239324
rect 238404 239322 238410 239324
rect 238845 239322 238911 239325
rect 238404 239320 238911 239322
rect 238404 239264 238850 239320
rect 238906 239264 238911 239320
rect 238404 239262 238911 239264
rect 238404 239260 238410 239262
rect 238845 239259 238911 239262
rect 239213 239322 239279 239325
rect 258809 239322 258875 239325
rect 239213 239320 258875 239322
rect 239213 239264 239218 239320
rect 239274 239264 258814 239320
rect 258870 239264 258875 239320
rect 239213 239262 258875 239264
rect 258996 239322 259056 239398
rect 259126 239396 259132 239460
rect 259196 239458 259243 239460
rect 262032 239458 262092 239670
rect 262489 239728 262628 239730
rect 262489 239672 262494 239728
rect 262550 239672 262628 239728
rect 262489 239670 262628 239672
rect 262489 239667 262555 239670
rect 262622 239668 262628 239670
rect 262692 239668 262698 239732
rect 262814 239730 262874 239806
rect 263823 239808 263828 239864
rect 263884 239808 264284 239864
rect 263823 239806 264284 239808
rect 263823 239803 263889 239806
rect 264278 239804 264284 239806
rect 264348 239804 264354 239868
rect 264467 239866 264533 239869
rect 264467 239864 264668 239866
rect 264467 239808 264472 239864
rect 264528 239808 264668 239864
rect 264467 239806 264668 239808
rect 264884 239842 264932 239898
rect 264988 239866 264993 239898
rect 264988 239842 265040 239866
rect 264884 239806 265040 239842
rect 264467 239803 264533 239806
rect 264608 239733 264668 239806
rect 262949 239730 263015 239733
rect 263501 239732 263567 239733
rect 263501 239730 263548 239732
rect 262814 239728 263015 239730
rect 262814 239672 262954 239728
rect 263010 239672 263015 239728
rect 262814 239670 263015 239672
rect 263456 239728 263548 239730
rect 263456 239672 263506 239728
rect 263456 239670 263548 239672
rect 262949 239667 263015 239670
rect 263501 239668 263548 239670
rect 263612 239668 263618 239732
rect 264329 239730 264395 239733
rect 264462 239730 264468 239732
rect 264329 239728 264468 239730
rect 264329 239672 264334 239728
rect 264390 239672 264468 239728
rect 264329 239670 264468 239672
rect 263501 239667 263567 239668
rect 264329 239667 264395 239670
rect 264462 239668 264468 239670
rect 264532 239668 264538 239732
rect 264605 239728 264671 239733
rect 264605 239672 264610 239728
rect 264666 239672 264671 239728
rect 264605 239667 264671 239672
rect 264973 239730 265039 239733
rect 265206 239730 265266 240078
rect 268653 240075 268719 240078
rect 267549 240004 267615 240005
rect 266486 239940 266492 240004
rect 266556 240002 266562 240004
rect 267549 240002 267596 240004
rect 266556 239942 267152 240002
rect 267504 240000 267596 240002
rect 267504 239944 267554 240000
rect 267504 239942 267596 239944
rect 266556 239940 266562 239942
rect 267092 239869 267152 239942
rect 267549 239940 267596 239942
rect 267660 239940 267666 240004
rect 267549 239939 267615 239940
rect 265939 239868 266005 239869
rect 265934 239866 265940 239868
rect 265848 239806 265940 239866
rect 265934 239804 265940 239806
rect 266004 239804 266010 239868
rect 266583 239866 266649 239869
rect 266540 239864 266649 239866
rect 266540 239808 266588 239864
rect 266644 239808 266649 239864
rect 265939 239803 266005 239804
rect 266540 239803 266649 239808
rect 267089 239864 267155 239869
rect 267089 239808 267094 239864
rect 267150 239808 267155 239864
rect 267089 239803 267155 239808
rect 267406 239804 267412 239868
rect 267476 239866 267482 239868
rect 267641 239866 267707 239869
rect 267476 239864 267707 239866
rect 267476 239808 267646 239864
rect 267702 239808 267707 239864
rect 267476 239806 267707 239808
rect 267476 239804 267482 239806
rect 267641 239803 267707 239806
rect 266540 239733 266600 239803
rect 264973 239728 265266 239730
rect 264973 239672 264978 239728
rect 265034 239672 265266 239728
rect 264973 239670 265266 239672
rect 265341 239730 265407 239733
rect 266077 239732 266143 239733
rect 265934 239730 265940 239732
rect 265341 239728 265940 239730
rect 265341 239672 265346 239728
rect 265402 239672 265940 239728
rect 265341 239670 265940 239672
rect 264973 239667 265039 239670
rect 265341 239667 265407 239670
rect 265934 239668 265940 239670
rect 266004 239668 266010 239732
rect 266077 239728 266124 239732
rect 266188 239730 266194 239732
rect 266077 239672 266082 239728
rect 266077 239668 266124 239672
rect 266188 239670 266234 239730
rect 266537 239728 266603 239733
rect 266537 239672 266542 239728
rect 266598 239672 266603 239728
rect 266188 239668 266194 239670
rect 266077 239667 266143 239668
rect 266537 239667 266603 239672
rect 266813 239730 266879 239733
rect 271137 239730 271203 239733
rect 266813 239728 271203 239730
rect 266813 239672 266818 239728
rect 266874 239672 271142 239728
rect 271198 239672 271203 239728
rect 266813 239670 271203 239672
rect 266813 239667 266879 239670
rect 271137 239667 271203 239670
rect 262622 239532 262628 239596
rect 262692 239594 262698 239596
rect 263504 239594 263564 239667
rect 262692 239534 263564 239594
rect 264237 239594 264303 239597
rect 269113 239594 269179 239597
rect 264237 239592 269179 239594
rect 264237 239536 264242 239592
rect 264298 239536 269118 239592
rect 269174 239536 269179 239592
rect 264237 239534 269179 239536
rect 262692 239532 262698 239534
rect 264237 239531 264303 239534
rect 269113 239531 269179 239534
rect 273897 239458 273963 239461
rect 259196 239456 259288 239458
rect 259238 239400 259288 239456
rect 259196 239398 259288 239400
rect 262032 239456 273963 239458
rect 262032 239400 273902 239456
rect 273958 239400 273963 239456
rect 262032 239398 273963 239400
rect 259196 239396 259243 239398
rect 259177 239395 259243 239396
rect 273897 239395 273963 239398
rect 260230 239322 260236 239324
rect 258996 239262 260236 239322
rect 239213 239259 239279 239262
rect 258809 239259 258875 239262
rect 260230 239260 260236 239262
rect 260300 239260 260306 239324
rect 260465 239322 260531 239325
rect 261661 239322 261727 239325
rect 260465 239320 261727 239322
rect 260465 239264 260470 239320
rect 260526 239264 261666 239320
rect 261722 239264 261727 239320
rect 260465 239262 261727 239264
rect 260465 239259 260531 239262
rect 261661 239259 261727 239262
rect 262070 239260 262076 239324
rect 262140 239322 262146 239324
rect 263542 239322 263548 239324
rect 262140 239262 263548 239322
rect 262140 239260 262146 239262
rect 263542 239260 263548 239262
rect 263612 239260 263618 239324
rect 263777 239322 263843 239325
rect 322197 239322 322263 239325
rect 263777 239320 322263 239322
rect 263777 239264 263782 239320
rect 263838 239264 322202 239320
rect 322258 239264 322263 239320
rect 263777 239262 322263 239264
rect 263777 239259 263843 239262
rect 322197 239259 322263 239262
rect 222193 239186 222259 239189
rect 223205 239186 223271 239189
rect 229461 239186 229527 239189
rect 229737 239188 229803 239189
rect 222193 239184 223271 239186
rect 222193 239128 222198 239184
rect 222254 239128 223210 239184
rect 223266 239128 223271 239184
rect 222193 239126 223271 239128
rect 222193 239123 222259 239126
rect 223205 239123 223271 239126
rect 224910 239184 229527 239186
rect 224910 239128 229466 239184
rect 229522 239128 229527 239184
rect 224910 239126 229527 239128
rect 215753 239050 215819 239053
rect 216121 239050 216187 239053
rect 219157 239050 219223 239053
rect 224910 239050 224970 239126
rect 229461 239123 229527 239126
rect 229686 239124 229692 239188
rect 229756 239186 229803 239188
rect 230381 239186 230447 239189
rect 236177 239186 236243 239189
rect 229756 239184 229848 239186
rect 229798 239128 229848 239184
rect 229756 239126 229848 239128
rect 230381 239184 236243 239186
rect 230381 239128 230386 239184
rect 230442 239128 236182 239184
rect 236238 239128 236243 239184
rect 230381 239126 236243 239128
rect 229756 239124 229803 239126
rect 229737 239123 229803 239124
rect 230381 239123 230447 239126
rect 236177 239123 236243 239126
rect 241646 239124 241652 239188
rect 241716 239186 241722 239188
rect 241973 239186 242039 239189
rect 241716 239184 242039 239186
rect 241716 239128 241978 239184
rect 242034 239128 242039 239184
rect 241716 239126 242039 239128
rect 241716 239124 241722 239126
rect 241973 239123 242039 239126
rect 252645 239186 252711 239189
rect 253473 239188 253539 239189
rect 253422 239186 253428 239188
rect 252645 239184 253428 239186
rect 253492 239186 253539 239188
rect 258993 239186 259059 239189
rect 262070 239186 262076 239188
rect 253492 239184 253584 239186
rect 252645 239128 252650 239184
rect 252706 239128 253428 239184
rect 253534 239128 253584 239184
rect 252645 239126 253428 239128
rect 252645 239123 252711 239126
rect 253422 239124 253428 239126
rect 253492 239126 253584 239128
rect 258993 239184 262076 239186
rect 258993 239128 258998 239184
rect 259054 239128 262076 239184
rect 258993 239126 262076 239128
rect 253492 239124 253539 239126
rect 253473 239123 253539 239124
rect 258993 239123 259059 239126
rect 262070 239124 262076 239126
rect 262140 239124 262146 239188
rect 263593 239186 263659 239189
rect 263869 239186 263935 239189
rect 264646 239186 264652 239188
rect 263593 239184 264652 239186
rect 263593 239128 263598 239184
rect 263654 239128 263874 239184
rect 263930 239128 264652 239184
rect 263593 239126 264652 239128
rect 263593 239123 263659 239126
rect 263869 239123 263935 239126
rect 264646 239124 264652 239126
rect 264716 239124 264722 239188
rect 265934 239124 265940 239188
rect 266004 239186 266010 239188
rect 325049 239186 325115 239189
rect 266004 239184 325115 239186
rect 266004 239128 325054 239184
rect 325110 239128 325115 239184
rect 266004 239126 325115 239128
rect 266004 239124 266010 239126
rect 325049 239123 325115 239126
rect 215753 239048 219082 239050
rect 215753 238992 215758 239048
rect 215814 238992 216126 239048
rect 216182 238992 219082 239048
rect 215753 238990 219082 238992
rect 215753 238987 215819 238990
rect 216121 238987 216187 238990
rect 219022 238914 219082 238990
rect 219157 239048 224970 239050
rect 219157 238992 219162 239048
rect 219218 238992 224970 239048
rect 219157 238990 224970 238992
rect 225505 239050 225571 239053
rect 284753 239050 284819 239053
rect 225505 239048 284819 239050
rect 225505 238992 225510 239048
rect 225566 238992 284758 239048
rect 284814 238992 284819 239048
rect 225505 238990 284819 238992
rect 219157 238987 219223 238990
rect 225505 238987 225571 238990
rect 284753 238987 284819 238990
rect 222837 238914 222903 238917
rect 219022 238912 222903 238914
rect 219022 238856 222842 238912
rect 222898 238856 222903 238912
rect 219022 238854 222903 238856
rect 222837 238851 222903 238854
rect 227897 238914 227963 238917
rect 229001 238914 229067 238917
rect 288985 238914 289051 238917
rect 227897 238912 289051 238914
rect 227897 238856 227902 238912
rect 227958 238856 229006 238912
rect 229062 238856 288990 238912
rect 289046 238856 289051 238912
rect 227897 238854 289051 238856
rect 227897 238851 227963 238854
rect 229001 238851 229067 238854
rect 288985 238851 289051 238854
rect 217317 238778 217383 238781
rect 226793 238778 226859 238781
rect 217317 238776 226859 238778
rect 217317 238720 217322 238776
rect 217378 238720 226798 238776
rect 226854 238720 226859 238776
rect 217317 238718 226859 238720
rect 217317 238715 217383 238718
rect 226793 238715 226859 238718
rect 227713 238778 227779 238781
rect 227846 238778 227852 238780
rect 227713 238776 227852 238778
rect 227713 238720 227718 238776
rect 227774 238720 227852 238776
rect 227713 238718 227852 238720
rect 227713 238715 227779 238718
rect 227846 238716 227852 238718
rect 227916 238716 227922 238780
rect 230105 238778 230171 238781
rect 230238 238778 230244 238780
rect 230105 238776 230244 238778
rect 230105 238720 230110 238776
rect 230166 238720 230244 238776
rect 230105 238718 230244 238720
rect 230105 238715 230171 238718
rect 230238 238716 230244 238718
rect 230308 238716 230314 238780
rect 231485 238778 231551 238781
rect 291377 238778 291443 238781
rect 231485 238776 291443 238778
rect 231485 238720 231490 238776
rect 231546 238720 291382 238776
rect 291438 238720 291443 238776
rect 231485 238718 291443 238720
rect 231485 238715 231551 238718
rect 291377 238715 291443 238718
rect 221181 238642 221247 238645
rect 224585 238642 224651 238645
rect 229001 238642 229067 238645
rect 221181 238640 224651 238642
rect 221181 238584 221186 238640
rect 221242 238584 224590 238640
rect 224646 238584 224651 238640
rect 221181 238582 224651 238584
rect 221181 238579 221247 238582
rect 224585 238579 224651 238582
rect 224910 238640 229067 238642
rect 224910 238584 229006 238640
rect 229062 238584 229067 238640
rect 224910 238582 229067 238584
rect 209681 238506 209747 238509
rect 223481 238506 223547 238509
rect 224910 238506 224970 238582
rect 229001 238579 229067 238582
rect 229461 238642 229527 238645
rect 231894 238642 231900 238644
rect 229461 238640 231900 238642
rect 229461 238584 229466 238640
rect 229522 238584 231900 238640
rect 229461 238582 231900 238584
rect 229461 238579 229527 238582
rect 231894 238580 231900 238582
rect 231964 238580 231970 238644
rect 233325 238642 233391 238645
rect 233918 238642 233924 238644
rect 233325 238640 233924 238642
rect 233325 238584 233330 238640
rect 233386 238584 233924 238640
rect 233325 238582 233924 238584
rect 233325 238579 233391 238582
rect 233918 238580 233924 238582
rect 233988 238642 233994 238644
rect 234245 238642 234311 238645
rect 233988 238640 234311 238642
rect 233988 238584 234250 238640
rect 234306 238584 234311 238640
rect 233988 238582 234311 238584
rect 233988 238580 233994 238582
rect 234245 238579 234311 238582
rect 234613 238644 234679 238645
rect 234613 238640 234660 238644
rect 234724 238642 234730 238644
rect 242433 238642 242499 238645
rect 242750 238642 242756 238644
rect 234613 238584 234618 238640
rect 234613 238580 234660 238584
rect 234724 238582 234770 238642
rect 242433 238640 242756 238642
rect 242433 238584 242438 238640
rect 242494 238584 242756 238640
rect 242433 238582 242756 238584
rect 234724 238580 234730 238582
rect 234613 238579 234679 238580
rect 242433 238579 242499 238582
rect 242750 238580 242756 238582
rect 242820 238580 242826 238644
rect 243302 238580 243308 238644
rect 243372 238642 243378 238644
rect 244273 238642 244339 238645
rect 243372 238640 244339 238642
rect 243372 238584 244278 238640
rect 244334 238584 244339 238640
rect 243372 238582 244339 238584
rect 243372 238580 243378 238582
rect 244273 238579 244339 238582
rect 244825 238642 244891 238645
rect 245142 238642 245148 238644
rect 244825 238640 245148 238642
rect 244825 238584 244830 238640
rect 244886 238584 245148 238640
rect 244825 238582 245148 238584
rect 244825 238579 244891 238582
rect 245142 238580 245148 238582
rect 245212 238580 245218 238644
rect 245326 238580 245332 238644
rect 245396 238642 245402 238644
rect 245469 238642 245535 238645
rect 245396 238640 245535 238642
rect 245396 238584 245474 238640
rect 245530 238584 245535 238640
rect 245396 238582 245535 238584
rect 245396 238580 245402 238582
rect 245469 238579 245535 238582
rect 246798 238580 246804 238644
rect 246868 238642 246874 238644
rect 246941 238642 247007 238645
rect 246868 238640 247007 238642
rect 246868 238584 246946 238640
rect 247002 238584 247007 238640
rect 246868 238582 247007 238584
rect 246868 238580 246874 238582
rect 246941 238579 247007 238582
rect 248270 238580 248276 238644
rect 248340 238642 248346 238644
rect 248413 238642 248479 238645
rect 248340 238640 248479 238642
rect 248340 238584 248418 238640
rect 248474 238584 248479 238640
rect 248340 238582 248479 238584
rect 248340 238580 248346 238582
rect 248413 238579 248479 238582
rect 248597 238642 248663 238645
rect 249374 238642 249380 238644
rect 248597 238640 249380 238642
rect 248597 238584 248602 238640
rect 248658 238584 249380 238640
rect 248597 238582 249380 238584
rect 248597 238579 248663 238582
rect 249374 238580 249380 238582
rect 249444 238580 249450 238644
rect 250110 238580 250116 238644
rect 250180 238642 250186 238644
rect 251081 238642 251147 238645
rect 253105 238644 253171 238645
rect 253054 238642 253060 238644
rect 250180 238640 251147 238642
rect 250180 238584 251086 238640
rect 251142 238584 251147 238640
rect 250180 238582 251147 238584
rect 253014 238582 253060 238642
rect 253124 238640 253171 238644
rect 268929 238642 268995 238645
rect 253166 238584 253171 238640
rect 250180 238580 250186 238582
rect 251081 238579 251147 238582
rect 253054 238580 253060 238582
rect 253124 238580 253171 238584
rect 253105 238579 253171 238580
rect 256650 238640 268995 238642
rect 256650 238584 268934 238640
rect 268990 238584 268995 238640
rect 256650 238582 268995 238584
rect 209681 238504 223547 238506
rect 209681 238448 209686 238504
rect 209742 238448 223486 238504
rect 223542 238448 223547 238504
rect 209681 238446 223547 238448
rect 209681 238443 209790 238446
rect 223481 238443 223547 238446
rect 223990 238446 224970 238506
rect 188337 237962 188403 237965
rect 209730 237962 209790 238443
rect 219433 238234 219499 238237
rect 220445 238234 220511 238237
rect 223990 238234 224050 238446
rect 226006 238444 226012 238508
rect 226076 238506 226082 238508
rect 226149 238506 226215 238509
rect 226517 238508 226583 238509
rect 226517 238506 226564 238508
rect 226076 238504 226215 238506
rect 226076 238448 226154 238504
rect 226210 238448 226215 238504
rect 226076 238446 226215 238448
rect 226472 238504 226564 238506
rect 226472 238448 226522 238504
rect 226472 238446 226564 238448
rect 226076 238444 226082 238446
rect 226149 238443 226215 238446
rect 226517 238444 226564 238446
rect 226628 238444 226634 238508
rect 231526 238444 231532 238508
rect 231596 238506 231602 238508
rect 232446 238506 232452 238508
rect 231596 238446 232452 238506
rect 231596 238444 231602 238446
rect 232446 238444 232452 238446
rect 232516 238444 232522 238508
rect 226517 238443 226583 238444
rect 224493 238370 224559 238373
rect 256650 238370 256710 238582
rect 268929 238579 268995 238582
rect 264278 238444 264284 238508
rect 264348 238506 264354 238508
rect 264513 238506 264579 238509
rect 264348 238504 264579 238506
rect 264348 238448 264518 238504
rect 264574 238448 264579 238504
rect 264348 238446 264579 238448
rect 264348 238444 264354 238446
rect 264513 238443 264579 238446
rect 264881 238506 264947 238509
rect 289445 238506 289511 238509
rect 264881 238504 289511 238506
rect 264881 238448 264886 238504
rect 264942 238448 289450 238504
rect 289506 238448 289511 238504
rect 264881 238446 289511 238448
rect 264881 238443 264947 238446
rect 289445 238443 289511 238446
rect 224493 238368 256710 238370
rect 224493 238312 224498 238368
rect 224554 238312 256710 238368
rect 224493 238310 256710 238312
rect 267549 238372 267615 238373
rect 267549 238368 267596 238372
rect 267660 238370 267666 238372
rect 267549 238312 267554 238368
rect 224493 238307 224559 238310
rect 267549 238308 267596 238312
rect 267660 238310 267706 238370
rect 267660 238308 267666 238310
rect 267549 238307 267615 238308
rect 219433 238232 224050 238234
rect 219433 238176 219438 238232
rect 219494 238176 220450 238232
rect 220506 238176 224050 238232
rect 219433 238174 224050 238176
rect 219433 238171 219499 238174
rect 220445 238171 220511 238174
rect 226374 238172 226380 238236
rect 226444 238234 226450 238236
rect 226793 238234 226859 238237
rect 226444 238232 226859 238234
rect 226444 238176 226798 238232
rect 226854 238176 226859 238232
rect 226444 238174 226859 238176
rect 226444 238172 226450 238174
rect 226793 238171 226859 238174
rect 228582 238172 228588 238236
rect 228652 238234 228658 238236
rect 228909 238234 228975 238237
rect 228652 238232 228975 238234
rect 228652 238176 228914 238232
rect 228970 238176 228975 238232
rect 228652 238174 228975 238176
rect 228652 238172 228658 238174
rect 228909 238171 228975 238174
rect 230105 238234 230171 238237
rect 230606 238234 230612 238236
rect 230105 238232 230612 238234
rect 230105 238176 230110 238232
rect 230166 238176 230612 238232
rect 230105 238174 230612 238176
rect 230105 238171 230171 238174
rect 230606 238172 230612 238174
rect 230676 238234 230682 238236
rect 264094 238234 264100 238236
rect 230676 238174 264100 238234
rect 230676 238172 230682 238174
rect 264094 238172 264100 238174
rect 264164 238172 264170 238236
rect 269481 238234 269547 238237
rect 264930 238232 269547 238234
rect 264930 238176 269486 238232
rect 269542 238176 269547 238232
rect 264930 238174 269547 238176
rect 216581 238098 216647 238101
rect 224534 238098 224540 238100
rect 216581 238096 224540 238098
rect 216581 238040 216586 238096
rect 216642 238040 224540 238096
rect 216581 238038 224540 238040
rect 216581 238035 216647 238038
rect 224534 238036 224540 238038
rect 224604 238036 224610 238100
rect 226609 238098 226675 238101
rect 226742 238098 226748 238100
rect 226609 238096 226748 238098
rect 226609 238040 226614 238096
rect 226670 238040 226748 238096
rect 226609 238038 226748 238040
rect 226609 238035 226675 238038
rect 226742 238036 226748 238038
rect 226812 238036 226818 238100
rect 227989 238098 228055 238101
rect 231669 238100 231735 238101
rect 228582 238098 228588 238100
rect 227989 238096 228588 238098
rect 227989 238040 227994 238096
rect 228050 238040 228588 238096
rect 227989 238038 228588 238040
rect 227989 238035 228055 238038
rect 228582 238036 228588 238038
rect 228652 238036 228658 238100
rect 231669 238096 231716 238100
rect 231780 238098 231786 238100
rect 236637 238098 236703 238101
rect 237230 238098 237236 238100
rect 231669 238040 231674 238096
rect 231669 238036 231716 238040
rect 231780 238038 231826 238098
rect 236637 238096 237236 238098
rect 236637 238040 236642 238096
rect 236698 238040 237236 238096
rect 236637 238038 237236 238040
rect 231780 238036 231786 238038
rect 231669 238035 231735 238036
rect 236637 238035 236703 238038
rect 237230 238036 237236 238038
rect 237300 238036 237306 238100
rect 258717 238098 258783 238101
rect 264930 238098 264990 238174
rect 269481 238171 269547 238174
rect 258717 238096 264990 238098
rect 258717 238040 258722 238096
rect 258778 238040 264990 238096
rect 258717 238038 264990 238040
rect 266629 238098 266695 238101
rect 315573 238098 315639 238101
rect 266629 238096 315639 238098
rect 266629 238040 266634 238096
rect 266690 238040 315578 238096
rect 315634 238040 315639 238096
rect 266629 238038 315639 238040
rect 258717 238035 258783 238038
rect 266629 238035 266695 238038
rect 315573 238035 315639 238038
rect 188337 237960 209790 237962
rect 188337 237904 188342 237960
rect 188398 237904 209790 237960
rect 188337 237902 209790 237904
rect 219985 237962 220051 237965
rect 227253 237962 227319 237965
rect 219985 237960 227319 237962
rect 219985 237904 219990 237960
rect 220046 237904 227258 237960
rect 227314 237904 227319 237960
rect 219985 237902 227319 237904
rect 188337 237899 188403 237902
rect 219985 237899 220051 237902
rect 227253 237899 227319 237902
rect 227662 237900 227668 237964
rect 227732 237962 227738 237964
rect 228817 237962 228883 237965
rect 227732 237960 228883 237962
rect 227732 237904 228822 237960
rect 228878 237904 228883 237960
rect 227732 237902 228883 237904
rect 227732 237900 227738 237902
rect 228817 237899 228883 237902
rect 231342 237900 231348 237964
rect 231412 237962 231418 237964
rect 231945 237962 232011 237965
rect 231412 237960 232011 237962
rect 231412 237904 231950 237960
rect 232006 237904 232011 237960
rect 231412 237902 232011 237904
rect 231412 237900 231418 237902
rect 231945 237899 232011 237902
rect 239489 237962 239555 237965
rect 250529 237964 250595 237965
rect 240910 237962 240916 237964
rect 239489 237960 240916 237962
rect 239489 237904 239494 237960
rect 239550 237904 240916 237960
rect 239489 237902 240916 237904
rect 239489 237899 239555 237902
rect 240910 237900 240916 237902
rect 240980 237900 240986 237964
rect 250478 237900 250484 237964
rect 250548 237962 250595 237964
rect 250548 237960 250640 237962
rect 250590 237904 250640 237960
rect 250548 237902 250640 237904
rect 250548 237900 250595 237902
rect 254710 237900 254716 237964
rect 254780 237962 254786 237964
rect 255221 237962 255287 237965
rect 254780 237960 255287 237962
rect 254780 237904 255226 237960
rect 255282 237904 255287 237960
rect 254780 237902 255287 237904
rect 254780 237900 254786 237902
rect 250529 237899 250595 237900
rect 255221 237899 255287 237902
rect 255497 237962 255563 237965
rect 256182 237962 256188 237964
rect 255497 237960 256188 237962
rect 255497 237904 255502 237960
rect 255558 237904 256188 237960
rect 255497 237902 256188 237904
rect 255497 237899 255563 237902
rect 256182 237900 256188 237902
rect 256252 237900 256258 237964
rect 264053 237962 264119 237965
rect 264462 237962 264468 237964
rect 264053 237960 264468 237962
rect 264053 237904 264058 237960
rect 264114 237904 264468 237960
rect 264053 237902 264468 237904
rect 264053 237899 264119 237902
rect 264462 237900 264468 237902
rect 264532 237900 264538 237964
rect 265709 237962 265775 237965
rect 324957 237962 325023 237965
rect 265709 237960 325023 237962
rect 265709 237904 265714 237960
rect 265770 237904 324962 237960
rect 325018 237904 325023 237960
rect 265709 237902 325023 237904
rect 265709 237899 265775 237902
rect 324957 237899 325023 237902
rect 209037 237826 209103 237829
rect 212165 237826 212231 237829
rect 219249 237826 219315 237829
rect 209037 237824 219315 237826
rect 209037 237768 209042 237824
rect 209098 237768 212170 237824
rect 212226 237768 219254 237824
rect 219310 237768 219315 237824
rect 209037 237766 219315 237768
rect 209037 237763 209103 237766
rect 212165 237763 212231 237766
rect 219249 237763 219315 237766
rect 222837 237826 222903 237829
rect 223665 237826 223731 237829
rect 222837 237824 263610 237826
rect 222837 237768 222842 237824
rect 222898 237768 223670 237824
rect 223726 237768 263610 237824
rect 222837 237766 263610 237768
rect 222837 237763 222903 237766
rect 223665 237763 223731 237766
rect 224861 237690 224927 237693
rect 255405 237690 255471 237693
rect 256734 237690 256740 237692
rect 224861 237688 237390 237690
rect 224861 237632 224866 237688
rect 224922 237632 237390 237688
rect 224861 237630 237390 237632
rect 224861 237627 224927 237630
rect 4153 237554 4219 237557
rect 222694 237554 222700 237556
rect 4153 237552 222700 237554
rect 4153 237496 4158 237552
rect 4214 237496 222700 237552
rect 4153 237494 222700 237496
rect 4153 237491 4219 237494
rect 222694 237492 222700 237494
rect 222764 237492 222770 237556
rect 230657 237554 230723 237557
rect 231526 237554 231532 237556
rect 230657 237552 231532 237554
rect 230657 237496 230662 237552
rect 230718 237496 231532 237552
rect 230657 237494 231532 237496
rect 230657 237491 230723 237494
rect 231526 237492 231532 237494
rect 231596 237492 231602 237556
rect 229645 237418 229711 237421
rect 229870 237418 229876 237420
rect 229645 237416 229876 237418
rect 229645 237360 229650 237416
rect 229706 237360 229876 237416
rect 229645 237358 229876 237360
rect 229645 237355 229711 237358
rect 229870 237356 229876 237358
rect 229940 237356 229946 237420
rect 237330 237418 237390 237630
rect 255405 237688 256740 237690
rect 255405 237632 255410 237688
rect 255466 237632 256740 237688
rect 255405 237630 256740 237632
rect 255405 237627 255471 237630
rect 256734 237628 256740 237630
rect 256804 237628 256810 237692
rect 260373 237556 260439 237557
rect 260373 237552 260420 237556
rect 260484 237554 260490 237556
rect 263550 237554 263610 237766
rect 263869 237690 263935 237693
rect 271781 237690 271847 237693
rect 263869 237688 271847 237690
rect 263869 237632 263874 237688
rect 263930 237632 271786 237688
rect 271842 237632 271847 237688
rect 263869 237630 271847 237632
rect 263869 237627 263935 237630
rect 271781 237627 271847 237630
rect 270953 237554 271019 237557
rect 260373 237496 260378 237552
rect 260373 237492 260420 237496
rect 260484 237494 260530 237554
rect 263550 237552 271019 237554
rect 263550 237496 270958 237552
rect 271014 237496 271019 237552
rect 263550 237494 271019 237496
rect 260484 237492 260490 237494
rect 260373 237491 260439 237492
rect 270953 237491 271019 237494
rect 263869 237418 263935 237421
rect 237330 237416 263935 237418
rect 237330 237360 263874 237416
rect 263930 237360 263935 237416
rect 237330 237358 263935 237360
rect 263869 237355 263935 237358
rect 184933 237282 184999 237285
rect 216489 237282 216555 237285
rect 236545 237282 236611 237285
rect 184933 237280 236611 237282
rect 184933 237224 184938 237280
rect 184994 237224 216494 237280
rect 216550 237224 236550 237280
rect 236606 237224 236611 237280
rect 184933 237222 236611 237224
rect 184933 237219 184999 237222
rect 216489 237219 216555 237222
rect 236545 237219 236611 237222
rect 250621 237282 250687 237285
rect 268653 237282 268719 237285
rect 250621 237280 268719 237282
rect 250621 237224 250626 237280
rect 250682 237224 268658 237280
rect 268714 237224 268719 237280
rect 250621 237222 268719 237224
rect 250621 237219 250687 237222
rect 268653 237219 268719 237222
rect 201493 237146 201559 237149
rect 238201 237146 238267 237149
rect 201493 237144 238267 237146
rect 201493 237088 201498 237144
rect 201554 237088 238206 237144
rect 238262 237088 238267 237144
rect 201493 237086 238267 237088
rect 201493 237083 201559 237086
rect 238201 237083 238267 237086
rect 259637 237146 259703 237149
rect 270033 237146 270099 237149
rect 259637 237144 270099 237146
rect 259637 237088 259642 237144
rect 259698 237088 270038 237144
rect 270094 237088 270099 237144
rect 259637 237086 270099 237088
rect 259637 237083 259703 237086
rect 270033 237083 270099 237086
rect 176653 237010 176719 237013
rect 216213 237010 216279 237013
rect 176653 237008 216279 237010
rect 176653 236952 176658 237008
rect 176714 236952 216218 237008
rect 216274 236952 216279 237008
rect 176653 236950 216279 236952
rect 176653 236947 176719 236950
rect 216213 236947 216279 236950
rect 218881 237010 218947 237013
rect 234429 237010 234495 237013
rect 218881 237008 234495 237010
rect 218881 236952 218886 237008
rect 218942 236952 234434 237008
rect 234490 236952 234495 237008
rect 218881 236950 234495 236952
rect 218881 236947 218947 236950
rect 234429 236947 234495 236950
rect 255313 237010 255379 237013
rect 268561 237010 268627 237013
rect 255313 237008 268627 237010
rect 255313 236952 255318 237008
rect 255374 236952 268566 237008
rect 268622 236952 268627 237008
rect 255313 236950 268627 236952
rect 255313 236947 255379 236950
rect 268561 236947 268627 236950
rect 173893 236874 173959 236877
rect 235206 236874 235212 236876
rect 173893 236872 235212 236874
rect 173893 236816 173898 236872
rect 173954 236816 235212 236872
rect 173893 236814 235212 236816
rect 173893 236811 173959 236814
rect 235206 236812 235212 236814
rect 235276 236812 235282 236876
rect 259453 236874 259519 236877
rect 259453 236872 335370 236874
rect 259453 236816 259458 236872
rect 259514 236816 335370 236872
rect 259453 236814 335370 236816
rect 259453 236811 259519 236814
rect 169753 236738 169819 236741
rect 235625 236738 235691 236741
rect 169753 236736 235691 236738
rect 169753 236680 169758 236736
rect 169814 236680 235630 236736
rect 235686 236680 235691 236736
rect 169753 236678 235691 236680
rect 169753 236675 169819 236678
rect 235625 236675 235691 236678
rect 242341 236740 242407 236741
rect 242341 236736 242388 236740
rect 242452 236738 242458 236740
rect 242341 236680 242346 236736
rect 242341 236676 242388 236680
rect 242452 236678 242498 236738
rect 242452 236676 242458 236678
rect 257102 236676 257108 236740
rect 257172 236738 257178 236740
rect 257981 236738 258047 236741
rect 257172 236736 258047 236738
rect 257172 236680 257986 236736
rect 258042 236680 258047 236736
rect 257172 236678 258047 236680
rect 257172 236676 257178 236678
rect 242341 236675 242407 236676
rect 257981 236675 258047 236678
rect 260782 236676 260788 236740
rect 260852 236738 260858 236740
rect 261845 236738 261911 236741
rect 260852 236736 261911 236738
rect 260852 236680 261850 236736
rect 261906 236680 261911 236736
rect 260852 236678 261911 236680
rect 260852 236676 260858 236678
rect 261845 236675 261911 236678
rect 264973 236738 265039 236741
rect 320909 236738 320975 236741
rect 264973 236736 320975 236738
rect 264973 236680 264978 236736
rect 265034 236680 320914 236736
rect 320970 236680 320975 236736
rect 264973 236678 320975 236680
rect 335310 236738 335370 236814
rect 354673 236738 354739 236741
rect 355317 236738 355383 236741
rect 335310 236736 355383 236738
rect 335310 236680 354678 236736
rect 354734 236680 355322 236736
rect 355378 236680 355383 236736
rect 335310 236678 355383 236680
rect 264973 236675 265039 236678
rect 320909 236675 320975 236678
rect 354673 236675 354739 236678
rect 355317 236675 355383 236678
rect 34513 236602 34579 236605
rect 214833 236602 214899 236605
rect 228725 236602 228791 236605
rect 34513 236600 200130 236602
rect 34513 236544 34518 236600
rect 34574 236544 200130 236600
rect 34513 236542 200130 236544
rect 34513 236539 34579 236542
rect 200070 236466 200130 236542
rect 214833 236600 228791 236602
rect 214833 236544 214838 236600
rect 214894 236544 228730 236600
rect 228786 236544 228791 236600
rect 214833 236542 228791 236544
rect 214833 236539 214899 236542
rect 228725 236539 228791 236542
rect 255681 236602 255747 236605
rect 264329 236602 264395 236605
rect 255681 236600 264395 236602
rect 255681 236544 255686 236600
rect 255742 236544 264334 236600
rect 264390 236544 264395 236600
rect 255681 236542 264395 236544
rect 255681 236539 255747 236542
rect 264329 236539 264395 236542
rect 211981 236466 212047 236469
rect 225045 236466 225111 236469
rect 200070 236464 225111 236466
rect 200070 236408 211986 236464
rect 212042 236408 225050 236464
rect 225106 236408 225111 236464
rect 200070 236406 225111 236408
rect 211981 236403 212047 236406
rect 225045 236403 225111 236406
rect 222377 236330 222443 236333
rect 222510 236330 222516 236332
rect 222377 236328 222516 236330
rect 222377 236272 222382 236328
rect 222438 236272 222516 236328
rect 222377 236270 222516 236272
rect 222377 236267 222443 236270
rect 222510 236268 222516 236270
rect 222580 236268 222586 236332
rect 223757 236330 223823 236333
rect 224166 236330 224172 236332
rect 223757 236328 224172 236330
rect 223757 236272 223762 236328
rect 223818 236272 224172 236328
rect 223757 236270 224172 236272
rect 223757 236267 223823 236270
rect 224166 236268 224172 236270
rect 224236 236268 224242 236332
rect 224585 236194 224651 236197
rect 224953 236196 225019 236197
rect 249609 236196 249675 236197
rect 224902 236194 224908 236196
rect 224585 236192 224908 236194
rect 224972 236194 225019 236196
rect 224972 236192 225064 236194
rect 224585 236136 224590 236192
rect 224646 236136 224908 236192
rect 225014 236136 225064 236192
rect 224585 236134 224908 236136
rect 224585 236131 224651 236134
rect 224902 236132 224908 236134
rect 224972 236134 225064 236136
rect 224972 236132 225019 236134
rect 249558 236132 249564 236196
rect 249628 236194 249675 236196
rect 249628 236192 249720 236194
rect 249670 236136 249720 236192
rect 249628 236134 249720 236136
rect 249628 236132 249675 236134
rect 250662 236132 250668 236196
rect 250732 236194 250738 236196
rect 250805 236194 250871 236197
rect 250732 236192 250871 236194
rect 250732 236136 250810 236192
rect 250866 236136 250871 236192
rect 250732 236134 250871 236136
rect 250732 236132 250738 236134
rect 224953 236131 225019 236132
rect 249609 236131 249675 236132
rect 250805 236131 250871 236134
rect 227989 236058 228055 236061
rect 228398 236058 228404 236060
rect 227989 236056 228404 236058
rect 227989 236000 227994 236056
rect 228050 236000 228404 236056
rect 227989 235998 228404 236000
rect 227989 235995 228055 235998
rect 228398 235996 228404 235998
rect 228468 235996 228474 236060
rect 254945 236058 255011 236061
rect 255078 236058 255084 236060
rect 254945 236056 255084 236058
rect 254945 236000 254950 236056
rect 255006 236000 255084 236056
rect 254945 235998 255084 236000
rect 254945 235995 255011 235998
rect 255078 235996 255084 235998
rect 255148 235996 255154 236060
rect 210693 235922 210759 235925
rect 211061 235922 211127 235925
rect 225873 235922 225939 235925
rect 241605 235924 241671 235925
rect 241605 235922 241652 235924
rect 210693 235920 225939 235922
rect 210693 235864 210698 235920
rect 210754 235864 211066 235920
rect 211122 235864 225878 235920
rect 225934 235864 225939 235920
rect 210693 235862 225939 235864
rect 241560 235920 241652 235922
rect 241560 235864 241610 235920
rect 241560 235862 241652 235864
rect 210693 235859 210759 235862
rect 211061 235859 211127 235862
rect 225873 235859 225939 235862
rect 241605 235860 241652 235862
rect 241716 235860 241722 235924
rect 254669 235922 254735 235925
rect 254894 235922 254900 235924
rect 254669 235920 254900 235922
rect 254669 235864 254674 235920
rect 254730 235864 254900 235920
rect 254669 235862 254900 235864
rect 241605 235859 241671 235860
rect 254669 235859 254735 235862
rect 254894 235860 254900 235862
rect 254964 235860 254970 235924
rect 213729 235786 213795 235789
rect 224033 235786 224099 235789
rect 213729 235784 224099 235786
rect 213729 235728 213734 235784
rect 213790 235728 224038 235784
rect 224094 235728 224099 235784
rect 213729 235726 224099 235728
rect 213729 235723 213795 235726
rect 224033 235723 224099 235726
rect 258073 235786 258139 235789
rect 316677 235786 316743 235789
rect 258073 235784 316743 235786
rect 258073 235728 258078 235784
rect 258134 235728 316682 235784
rect 316738 235728 316743 235784
rect 258073 235726 316743 235728
rect 258073 235723 258139 235726
rect 316677 235723 316743 235726
rect 217317 235650 217383 235653
rect 223430 235650 223436 235652
rect 217317 235648 223436 235650
rect 217317 235592 217322 235648
rect 217378 235592 223436 235648
rect 217317 235590 223436 235592
rect 217317 235587 217383 235590
rect 223430 235588 223436 235590
rect 223500 235588 223506 235652
rect 269113 235650 269179 235653
rect 297449 235650 297515 235653
rect 269113 235648 297515 235650
rect 269113 235592 269118 235648
rect 269174 235592 297454 235648
rect 297510 235592 297515 235648
rect 269113 235590 297515 235592
rect 269113 235587 269179 235590
rect 297449 235587 297515 235590
rect 263869 235514 263935 235517
rect 278037 235514 278103 235517
rect 263869 235512 278103 235514
rect 263869 235456 263874 235512
rect 263930 235456 278042 235512
rect 278098 235456 278103 235512
rect 263869 235454 278103 235456
rect 263869 235451 263935 235454
rect 278037 235451 278103 235454
rect 233509 235378 233575 235381
rect 234286 235378 234292 235380
rect 233509 235376 234292 235378
rect 233509 235320 233514 235376
rect 233570 235320 234292 235376
rect 233509 235318 234292 235320
rect 233509 235315 233575 235318
rect 234286 235316 234292 235318
rect 234356 235316 234362 235380
rect 251817 235378 251883 235381
rect 311157 235378 311223 235381
rect 251817 235376 311223 235378
rect 251817 235320 251822 235376
rect 251878 235320 311162 235376
rect 311218 235320 311223 235376
rect 251817 235318 311223 235320
rect 251817 235315 251883 235318
rect 311157 235315 311223 235318
rect 152457 235242 152523 235245
rect 232262 235242 232268 235244
rect 152457 235240 232268 235242
rect 152457 235184 152462 235240
rect 152518 235184 232268 235240
rect 152457 235182 232268 235184
rect 152457 235179 152523 235182
rect 232262 235180 232268 235182
rect 232332 235180 232338 235244
rect 256734 235180 256740 235244
rect 256804 235242 256810 235244
rect 257153 235242 257219 235245
rect 256804 235240 257219 235242
rect 256804 235184 257158 235240
rect 257214 235184 257219 235240
rect 256804 235182 257219 235184
rect 256804 235180 256810 235182
rect 257153 235179 257219 235182
rect 258349 235242 258415 235245
rect 260046 235242 260052 235244
rect 258349 235240 260052 235242
rect 258349 235184 258354 235240
rect 258410 235184 260052 235240
rect 258349 235182 260052 235184
rect 258349 235179 258415 235182
rect 260046 235180 260052 235182
rect 260116 235180 260122 235244
rect 262581 235242 262647 235245
rect 263174 235242 263180 235244
rect 262581 235240 263180 235242
rect 262581 235184 262586 235240
rect 262642 235184 263180 235240
rect 262581 235182 263180 235184
rect 262581 235179 262647 235182
rect 263174 235180 263180 235182
rect 263244 235180 263250 235244
rect 234889 234834 234955 234837
rect 235758 234834 235764 234836
rect 234889 234832 235764 234834
rect 234889 234776 234894 234832
rect 234950 234776 235764 234832
rect 234889 234774 235764 234776
rect 234889 234771 234955 234774
rect 235758 234772 235764 234774
rect 235828 234772 235834 234836
rect 234797 234562 234863 234565
rect 235574 234562 235580 234564
rect 234797 234560 235580 234562
rect 234797 234504 234802 234560
rect 234858 234504 235580 234560
rect 234797 234502 235580 234504
rect 234797 234499 234863 234502
rect 235574 234500 235580 234502
rect 235644 234500 235650 234564
rect 243118 234500 243124 234564
rect 243188 234562 243194 234564
rect 246757 234562 246823 234565
rect 243188 234560 246823 234562
rect 243188 234504 246762 234560
rect 246818 234504 246823 234560
rect 243188 234502 246823 234504
rect 243188 234500 243194 234502
rect 246757 234499 246823 234502
rect 263961 234562 264027 234565
rect 335905 234562 335971 234565
rect 336641 234562 336707 234565
rect 263961 234560 336707 234562
rect 263961 234504 263966 234560
rect 264022 234504 335910 234560
rect 335966 234504 336646 234560
rect 336702 234504 336707 234560
rect 263961 234502 336707 234504
rect 263961 234499 264027 234502
rect 335905 234499 335971 234502
rect 336641 234499 336707 234502
rect 260097 234426 260163 234429
rect 330477 234426 330543 234429
rect 260097 234424 330543 234426
rect 260097 234368 260102 234424
rect 260158 234368 330482 234424
rect 330538 234368 330543 234424
rect 260097 234366 330543 234368
rect 260097 234363 260163 234366
rect 330477 234363 330543 234366
rect 260005 234290 260071 234293
rect 330109 234290 330175 234293
rect 260005 234288 335370 234290
rect 260005 234232 260010 234288
rect 260066 234232 330114 234288
rect 330170 234232 335370 234288
rect 260005 234230 335370 234232
rect 260005 234227 260071 234230
rect 330109 234227 330175 234230
rect 262673 234154 262739 234157
rect 327441 234154 327507 234157
rect 327717 234154 327783 234157
rect 262673 234152 327783 234154
rect 262673 234096 262678 234152
rect 262734 234096 327446 234152
rect 327502 234096 327722 234152
rect 327778 234096 327783 234152
rect 262673 234094 327783 234096
rect 335310 234154 335370 234230
rect 483013 234154 483079 234157
rect 335310 234152 483079 234154
rect 335310 234096 483018 234152
rect 483074 234096 483079 234152
rect 335310 234094 483079 234096
rect 262673 234091 262739 234094
rect 327441 234091 327507 234094
rect 327717 234091 327783 234094
rect 483013 234091 483079 234094
rect 97993 234018 98059 234021
rect 230238 234018 230244 234020
rect 97993 234016 230244 234018
rect 97993 233960 97998 234016
rect 98054 233960 230244 234016
rect 97993 233958 230244 233960
rect 97993 233955 98059 233958
rect 230238 233956 230244 233958
rect 230308 233956 230314 234020
rect 262489 234018 262555 234021
rect 331397 234018 331463 234021
rect 502977 234018 503043 234021
rect 262489 234016 503043 234018
rect 262489 233960 262494 234016
rect 262550 233960 331402 234016
rect 331458 233960 502982 234016
rect 503038 233960 503043 234016
rect 262489 233958 503043 233960
rect 262489 233955 262555 233958
rect 331397 233955 331463 233958
rect 502977 233955 503043 233958
rect 44173 233882 44239 233885
rect 210693 233882 210759 233885
rect 44173 233880 210759 233882
rect 44173 233824 44178 233880
rect 44234 233824 210698 233880
rect 210754 233824 210759 233880
rect 44173 233822 210759 233824
rect 44173 233819 44239 233822
rect 210693 233819 210759 233822
rect 256785 233882 256851 233885
rect 312629 233882 312695 233885
rect 256785 233880 312695 233882
rect 256785 233824 256790 233880
rect 256846 233824 312634 233880
rect 312690 233824 312695 233880
rect 256785 233822 312695 233824
rect 256785 233819 256851 233822
rect 312629 233819 312695 233822
rect 336641 233882 336707 233885
rect 532693 233882 532759 233885
rect 336641 233880 532759 233882
rect 336641 233824 336646 233880
rect 336702 233824 532698 233880
rect 532754 233824 532759 233880
rect 336641 233822 532759 233824
rect 336641 233819 336707 233822
rect 532693 233819 532759 233822
rect 252093 233746 252159 233749
rect 268469 233746 268535 233749
rect 252093 233744 268535 233746
rect 252093 233688 252098 233744
rect 252154 233688 268474 233744
rect 268530 233688 268535 233744
rect 252093 233686 268535 233688
rect 252093 233683 252159 233686
rect 268469 233683 268535 233686
rect 253841 233202 253907 233205
rect 277301 233202 277367 233205
rect 278129 233202 278195 233205
rect 253841 233200 278195 233202
rect 253841 233144 253846 233200
rect 253902 233144 277306 233200
rect 277362 233144 278134 233200
rect 278190 233144 278195 233200
rect 253841 233142 278195 233144
rect 253841 233139 253907 233142
rect 277301 233139 277367 233142
rect 278129 233139 278195 233142
rect 303705 233202 303771 233205
rect 304390 233202 304396 233204
rect 303705 233200 304396 233202
rect 303705 233144 303710 233200
rect 303766 233144 304396 233200
rect 303705 233142 304396 233144
rect 303705 233139 303771 233142
rect 304390 233140 304396 233142
rect 304460 233140 304466 233204
rect 261937 233066 262003 233069
rect 261937 233064 325710 233066
rect 261937 233008 261942 233064
rect 261998 233008 325710 233064
rect 261937 233006 325710 233008
rect 261937 233003 262003 233006
rect 256550 232868 256556 232932
rect 256620 232930 256626 232932
rect 315297 232930 315363 232933
rect 256620 232928 315363 232930
rect 256620 232872 315302 232928
rect 315358 232872 315363 232928
rect 256620 232870 315363 232872
rect 256620 232868 256626 232870
rect 315297 232867 315363 232870
rect 262397 232794 262463 232797
rect 320817 232794 320883 232797
rect 262397 232792 320883 232794
rect 262397 232736 262402 232792
rect 262458 232736 320822 232792
rect 320878 232736 320883 232792
rect 262397 232734 320883 232736
rect 262397 232731 262463 232734
rect 320817 232731 320883 232734
rect 242750 232596 242756 232660
rect 242820 232658 242826 232660
rect 299974 232658 299980 232660
rect 242820 232598 299980 232658
rect 242820 232596 242826 232598
rect 299974 232596 299980 232598
rect 300044 232596 300050 232660
rect 325650 232658 325710 233006
rect 330017 232658 330083 232661
rect 507853 232658 507919 232661
rect 325650 232656 507919 232658
rect 325650 232600 330022 232656
rect 330078 232600 507858 232656
rect 507914 232600 507919 232656
rect 325650 232598 507919 232600
rect 330017 232595 330083 232598
rect 507853 232595 507919 232598
rect 138013 232522 138079 232525
rect 217133 232522 217199 232525
rect 138013 232520 217199 232522
rect 138013 232464 138018 232520
rect 138074 232464 217138 232520
rect 217194 232464 217199 232520
rect 138013 232462 217199 232464
rect 138013 232459 138079 232462
rect 217133 232459 217199 232462
rect 266813 232522 266879 232525
rect 314101 232522 314167 232525
rect 555417 232522 555483 232525
rect 266813 232520 314167 232522
rect 266813 232464 266818 232520
rect 266874 232464 314106 232520
rect 314162 232464 314167 232520
rect 266813 232462 314167 232464
rect 266813 232459 266879 232462
rect 314101 232459 314167 232462
rect 335310 232520 555483 232522
rect 335310 232464 555422 232520
rect 555478 232464 555483 232520
rect 335310 232462 555483 232464
rect 266261 232386 266327 232389
rect 334341 232386 334407 232389
rect 335310 232386 335370 232462
rect 555417 232459 555483 232462
rect 266261 232384 335370 232386
rect 266261 232328 266266 232384
rect 266322 232328 334346 232384
rect 334402 232328 335370 232384
rect 266261 232326 335370 232328
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 266261 232323 266327 232326
rect 334341 232323 334407 232326
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 260649 231842 260715 231845
rect 328361 231842 328427 231845
rect 260649 231840 328427 231842
rect 260649 231784 260654 231840
rect 260710 231784 328366 231840
rect 328422 231784 328427 231840
rect 260649 231782 328427 231784
rect 260649 231779 260715 231782
rect 328361 231779 328427 231782
rect 328729 231842 328795 231845
rect 329281 231842 329347 231845
rect 328729 231840 329347 231842
rect 328729 231784 328734 231840
rect 328790 231784 329286 231840
rect 329342 231784 329347 231840
rect 328729 231782 329347 231784
rect 328729 231779 328795 231782
rect 329281 231779 329347 231782
rect 261017 231706 261083 231709
rect 328913 231706 328979 231709
rect 261017 231704 328979 231706
rect 261017 231648 261022 231704
rect 261078 231648 328918 231704
rect 328974 231648 328979 231704
rect 261017 231646 328979 231648
rect 261017 231643 261083 231646
rect 328913 231643 328979 231646
rect 264881 231570 264947 231573
rect 331489 231570 331555 231573
rect 264881 231568 331555 231570
rect 264881 231512 264886 231568
rect 264942 231512 331494 231568
rect 331550 231512 331555 231568
rect 264881 231510 331555 231512
rect 264881 231507 264947 231510
rect 331489 231507 331555 231510
rect 155217 231434 155283 231437
rect 217593 231434 217659 231437
rect 155217 231432 217659 231434
rect 155217 231376 155222 231432
rect 155278 231376 217598 231432
rect 217654 231376 217659 231432
rect 155217 231374 217659 231376
rect 155217 231371 155283 231374
rect 217593 231371 217659 231374
rect 262765 231434 262831 231437
rect 328729 231434 328795 231437
rect 262765 231432 328795 231434
rect 262765 231376 262770 231432
rect 262826 231376 328734 231432
rect 328790 231376 328795 231432
rect 262765 231374 328795 231376
rect 262765 231371 262831 231374
rect 328729 231371 328795 231374
rect 208393 231298 208459 231301
rect 237925 231298 237991 231301
rect 299790 231298 299796 231300
rect 208393 231296 299796 231298
rect 208393 231240 208398 231296
rect 208454 231240 237930 231296
rect 237986 231240 299796 231296
rect 208393 231238 299796 231240
rect 208393 231235 208459 231238
rect 237925 231235 237991 231238
rect 299790 231236 299796 231238
rect 299860 231236 299866 231300
rect 51073 231162 51139 231165
rect 215661 231162 215727 231165
rect 51073 231160 215727 231162
rect 51073 231104 51078 231160
rect 51134 231104 215666 231160
rect 215722 231104 215727 231160
rect 51073 231102 215727 231104
rect 51073 231099 51139 231102
rect 215661 231099 215727 231102
rect 246614 231100 246620 231164
rect 246684 231162 246690 231164
rect 302233 231162 302299 231165
rect 246684 231160 302299 231162
rect 246684 231104 302238 231160
rect 302294 231104 302299 231160
rect 246684 231102 302299 231104
rect 246684 231100 246690 231102
rect 302233 231099 302299 231102
rect 328361 231162 328427 231165
rect 333053 231162 333119 231165
rect 490005 231162 490071 231165
rect 328361 231160 490071 231162
rect 328361 231104 328366 231160
rect 328422 231104 333058 231160
rect 333114 231104 490010 231160
rect 490066 231104 490071 231160
rect 328361 231102 490071 231104
rect 328361 231099 328427 231102
rect 333053 231099 333119 231102
rect 490005 231099 490071 231102
rect 265709 231026 265775 231029
rect 266118 231026 266124 231028
rect 265709 231024 266124 231026
rect 265709 230968 265714 231024
rect 265770 230968 266124 231024
rect 265709 230966 266124 230968
rect 265709 230963 265775 230966
rect 266118 230964 266124 230966
rect 266188 230964 266194 231028
rect 263777 230346 263843 230349
rect 334249 230346 334315 230349
rect 334801 230346 334867 230349
rect 263777 230344 334867 230346
rect 263777 230288 263782 230344
rect 263838 230288 334254 230344
rect 334310 230288 334806 230344
rect 334862 230288 334867 230344
rect 263777 230286 334867 230288
rect 263777 230283 263843 230286
rect 334249 230283 334315 230286
rect 334801 230283 334867 230286
rect 263409 230210 263475 230213
rect 322657 230210 322723 230213
rect 263409 230208 322723 230210
rect 263409 230152 263414 230208
rect 263470 230152 322662 230208
rect 322718 230152 322723 230208
rect 263409 230150 322723 230152
rect 263409 230147 263475 230150
rect 322657 230147 322723 230150
rect 259085 230074 259151 230077
rect 309869 230074 309935 230077
rect 259085 230072 309935 230074
rect 259085 230016 259090 230072
rect 259146 230016 309874 230072
rect 309930 230016 309935 230072
rect 259085 230014 309935 230016
rect 259085 230011 259151 230014
rect 309869 230011 309935 230014
rect 110413 229938 110479 229941
rect 214833 229938 214899 229941
rect 110413 229936 214899 229938
rect 110413 229880 110418 229936
rect 110474 229880 214838 229936
rect 214894 229880 214899 229936
rect 110413 229878 214899 229880
rect 110413 229875 110479 229878
rect 214833 229875 214899 229878
rect 258993 229938 259059 229941
rect 302969 229938 303035 229941
rect 336917 229938 336983 229941
rect 440233 229938 440299 229941
rect 258993 229936 303035 229938
rect 258993 229880 258998 229936
rect 259054 229880 302974 229936
rect 303030 229880 303035 229936
rect 258993 229878 303035 229880
rect 258993 229875 259059 229878
rect 302969 229875 303035 229878
rect 315990 229936 440299 229938
rect 315990 229880 336922 229936
rect 336978 229880 440238 229936
rect 440294 229880 440299 229936
rect 315990 229878 440299 229880
rect 71037 229802 71103 229805
rect 217225 229802 217291 229805
rect 71037 229800 217291 229802
rect 71037 229744 71042 229800
rect 71098 229744 217230 229800
rect 217286 229744 217291 229800
rect 71037 229742 217291 229744
rect 71037 229739 71103 229742
rect 217225 229739 217291 229742
rect 242382 229740 242388 229804
rect 242452 229802 242458 229804
rect 271505 229802 271571 229805
rect 242452 229800 271571 229802
rect 242452 229744 271510 229800
rect 271566 229744 271571 229800
rect 242452 229742 271571 229744
rect 242452 229740 242458 229742
rect 271505 229739 271571 229742
rect 257981 229666 258047 229669
rect 315990 229666 316050 229878
rect 336917 229875 336983 229878
rect 440233 229875 440299 229878
rect 334801 229802 334867 229805
rect 536097 229802 536163 229805
rect 334801 229800 536163 229802
rect 334801 229744 334806 229800
rect 334862 229744 536102 229800
rect 536158 229744 536163 229800
rect 334801 229742 536163 229744
rect 334801 229739 334867 229742
rect 536097 229739 536163 229742
rect 257981 229664 316050 229666
rect 257981 229608 257986 229664
rect 258042 229608 316050 229664
rect 257981 229606 316050 229608
rect 257981 229603 258047 229606
rect 306097 229260 306163 229261
rect 306046 229196 306052 229260
rect 306116 229258 306163 229260
rect 306116 229256 306208 229258
rect 306158 229200 306208 229256
rect 306116 229198 306208 229200
rect 306116 229196 306163 229198
rect 306097 229195 306163 229196
rect 260414 228924 260420 228988
rect 260484 228986 260490 228988
rect 260741 228986 260807 228989
rect 260484 228984 260807 228986
rect 260484 228928 260746 228984
rect 260802 228928 260807 228984
rect 260484 228926 260807 228928
rect 260484 228924 260490 228926
rect 260741 228923 260807 228926
rect 263041 228986 263107 228989
rect 335629 228986 335695 228989
rect 263041 228984 335695 228986
rect 263041 228928 263046 228984
rect 263102 228928 335634 228984
rect 335690 228928 335695 228984
rect 263041 228926 335695 228928
rect 263041 228923 263107 228926
rect 265617 228850 265683 228853
rect 265617 228848 316050 228850
rect 265617 228792 265622 228848
rect 265678 228792 316050 228848
rect 265617 228790 316050 228792
rect 265617 228787 265683 228790
rect 253054 228652 253060 228716
rect 253124 228714 253130 228716
rect 253657 228714 253723 228717
rect 278405 228714 278471 228717
rect 253124 228712 278471 228714
rect 253124 228656 253662 228712
rect 253718 228656 278410 228712
rect 278466 228656 278471 228712
rect 253124 228654 278471 228656
rect 253124 228652 253130 228654
rect 253657 228651 253723 228654
rect 278405 228651 278471 228654
rect 257521 228578 257587 228581
rect 280981 228578 281047 228581
rect 257521 228576 281047 228578
rect 257521 228520 257526 228576
rect 257582 228520 280986 228576
rect 281042 228520 281047 228576
rect 257521 228518 281047 228520
rect 257521 228515 257587 228518
rect 280981 228515 281047 228518
rect 71773 228306 71839 228309
rect 213637 228306 213703 228309
rect 71773 228304 213703 228306
rect 71773 228248 71778 228304
rect 71834 228248 213642 228304
rect 213698 228248 213703 228304
rect 71773 228246 213703 228248
rect 71773 228243 71839 228246
rect 213637 228243 213703 228246
rect 243486 228244 243492 228308
rect 243556 228306 243562 228308
rect 269113 228306 269179 228309
rect 243556 228304 269179 228306
rect 243556 228248 269118 228304
rect 269174 228248 269179 228304
rect 243556 228246 269179 228248
rect 315990 228306 316050 228790
rect 335310 228442 335370 228926
rect 335629 228923 335695 228926
rect 523125 228442 523191 228445
rect 335310 228440 523191 228442
rect 335310 228384 523130 228440
rect 523186 228384 523191 228440
rect 335310 228382 523191 228384
rect 523125 228379 523191 228382
rect 335721 228306 335787 228309
rect 557533 228306 557599 228309
rect 315990 228304 557599 228306
rect 315990 228248 335726 228304
rect 335782 228248 557538 228304
rect 557594 228248 557599 228304
rect 315990 228246 557599 228248
rect 243556 228244 243562 228246
rect 269113 228243 269179 228246
rect 335721 228243 335787 228246
rect 557533 228243 557599 228246
rect -960 227884 480 228124
rect 302049 227628 302115 227629
rect 301998 227626 302004 227628
rect 301958 227566 302004 227626
rect 302068 227624 302115 227628
rect 302110 227568 302115 227624
rect 301998 227564 302004 227566
rect 302068 227564 302115 227568
rect 302049 227563 302115 227564
rect 262121 227490 262187 227493
rect 322289 227490 322355 227493
rect 262121 227488 322355 227490
rect 262121 227432 262126 227488
rect 262182 227432 322294 227488
rect 322350 227432 322355 227488
rect 262121 227430 322355 227432
rect 262121 227427 262187 227430
rect 322289 227427 322355 227430
rect 242566 227292 242572 227356
rect 242636 227354 242642 227356
rect 302182 227354 302188 227356
rect 242636 227294 302188 227354
rect 242636 227292 242642 227294
rect 302182 227292 302188 227294
rect 302252 227292 302258 227356
rect 253197 227218 253263 227221
rect 311014 227218 311020 227220
rect 253197 227216 311020 227218
rect 253197 227160 253202 227216
rect 253258 227160 311020 227216
rect 253197 227158 311020 227160
rect 253197 227155 253263 227158
rect 311014 227156 311020 227158
rect 311084 227156 311090 227220
rect 233734 227020 233740 227084
rect 233804 227082 233810 227084
rect 289169 227082 289235 227085
rect 233804 227080 289235 227082
rect 233804 227024 289174 227080
rect 289230 227024 289235 227080
rect 233804 227022 289235 227024
rect 233804 227020 233810 227022
rect 289169 227019 289235 227022
rect 25497 226946 25563 226949
rect 213729 226946 213795 226949
rect 25497 226944 213795 226946
rect 25497 226888 25502 226944
rect 25558 226888 213734 226944
rect 213790 226888 213795 226944
rect 25497 226886 213795 226888
rect 25497 226883 25563 226886
rect 213729 226883 213795 226886
rect 216673 226946 216739 226949
rect 239070 226946 239076 226948
rect 216673 226944 239076 226946
rect 216673 226888 216678 226944
rect 216734 226888 239076 226944
rect 216673 226886 239076 226888
rect 216673 226883 216739 226886
rect 239070 226884 239076 226886
rect 239140 226884 239146 226948
rect 266537 226946 266603 226949
rect 328637 226946 328703 226949
rect 562317 226946 562383 226949
rect 266537 226944 562383 226946
rect 266537 226888 266542 226944
rect 266598 226888 328642 226944
rect 328698 226888 562322 226944
rect 562378 226888 562383 226944
rect 266537 226886 562383 226888
rect 266537 226883 266603 226886
rect 328637 226883 328703 226886
rect 562317 226883 562383 226886
rect 250110 226204 250116 226268
rect 250180 226266 250186 226268
rect 250989 226266 251055 226269
rect 250180 226264 251055 226266
rect 250180 226208 250994 226264
rect 251050 226208 251055 226264
rect 250180 226206 251055 226208
rect 250180 226204 250186 226206
rect 250989 226203 251055 226206
rect 305269 226266 305335 226269
rect 306230 226266 306236 226268
rect 305269 226264 306236 226266
rect 305269 226208 305274 226264
rect 305330 226208 306236 226264
rect 305269 226206 306236 226208
rect 305269 226203 305335 226206
rect 306230 226204 306236 226206
rect 306300 226204 306306 226268
rect 261845 226130 261911 226133
rect 322381 226130 322447 226133
rect 261845 226128 322447 226130
rect 261845 226072 261850 226128
rect 261906 226072 322386 226128
rect 322442 226072 322447 226128
rect 261845 226070 322447 226072
rect 261845 226067 261911 226070
rect 322381 226067 322447 226070
rect 255078 225932 255084 225996
rect 255148 225994 255154 225996
rect 282269 225994 282335 225997
rect 255148 225992 282335 225994
rect 255148 225936 282274 225992
rect 282330 225936 282335 225992
rect 255148 225934 282335 225936
rect 255148 225932 255154 225934
rect 282269 225931 282335 225934
rect 263174 225796 263180 225860
rect 263244 225858 263250 225860
rect 286685 225858 286751 225861
rect 263244 225856 286751 225858
rect 263244 225800 286690 225856
rect 286746 225800 286751 225856
rect 263244 225798 286751 225800
rect 263244 225796 263250 225798
rect 286685 225795 286751 225798
rect 263225 225722 263291 225725
rect 263225 225720 335370 225722
rect 263225 225664 263230 225720
rect 263286 225664 335370 225720
rect 263225 225662 335370 225664
rect 263225 225659 263291 225662
rect 57973 225586 58039 225589
rect 213085 225586 213151 225589
rect 57973 225584 213151 225586
rect 57973 225528 57978 225584
rect 58034 225528 213090 225584
rect 213146 225528 213151 225584
rect 57973 225526 213151 225528
rect 335310 225586 335370 225662
rect 335445 225586 335511 225589
rect 525793 225586 525859 225589
rect 335310 225584 525859 225586
rect 335310 225528 335450 225584
rect 335506 225528 525798 225584
rect 525854 225528 525859 225584
rect 335310 225526 525859 225528
rect 57973 225523 58039 225526
rect 213085 225523 213151 225526
rect 335445 225523 335511 225526
rect 525793 225523 525859 225526
rect 214741 224906 214807 224909
rect 215201 224906 215267 224909
rect 229870 224906 229876 224908
rect 214741 224904 229876 224906
rect 214741 224848 214746 224904
rect 214802 224848 215206 224904
rect 215262 224848 229876 224904
rect 214741 224846 229876 224848
rect 214741 224843 214807 224846
rect 215201 224843 215267 224846
rect 229870 224844 229876 224846
rect 229940 224844 229946 224908
rect 233601 224906 233667 224909
rect 294638 224906 294644 224908
rect 233601 224904 294644 224906
rect 233601 224848 233606 224904
rect 233662 224848 294644 224904
rect 233601 224846 294644 224848
rect 233601 224843 233667 224846
rect 294638 224844 294644 224846
rect 294708 224844 294714 224908
rect 294321 224770 294387 224773
rect 238710 224768 294387 224770
rect 238710 224712 294326 224768
rect 294382 224712 294387 224768
rect 238710 224710 294387 224712
rect 209865 224498 209931 224501
rect 237414 224498 237420 224500
rect 209865 224496 237420 224498
rect 209865 224440 209870 224496
rect 209926 224440 237420 224496
rect 209865 224438 237420 224440
rect 209865 224435 209931 224438
rect 237414 224436 237420 224438
rect 237484 224436 237490 224500
rect 158713 224362 158779 224365
rect 235574 224362 235580 224364
rect 158713 224360 235580 224362
rect 158713 224304 158718 224360
rect 158774 224304 235580 224360
rect 158713 224302 235580 224304
rect 158713 224299 158779 224302
rect 235574 224300 235580 224302
rect 235644 224362 235650 224364
rect 238710 224362 238770 224710
rect 294321 224707 294387 224710
rect 260230 224572 260236 224636
rect 260300 224634 260306 224636
rect 318057 224634 318123 224637
rect 260300 224632 318123 224634
rect 260300 224576 318062 224632
rect 318118 224576 318123 224632
rect 260300 224574 318123 224576
rect 260300 224572 260306 224574
rect 318057 224571 318123 224574
rect 262806 224436 262812 224500
rect 262876 224498 262882 224500
rect 319294 224498 319300 224500
rect 262876 224438 319300 224498
rect 262876 224436 262882 224438
rect 319294 224436 319300 224438
rect 319364 224436 319370 224500
rect 235644 224302 238770 224362
rect 235644 224300 235650 224302
rect 262070 224300 262076 224364
rect 262140 224362 262146 224364
rect 318241 224362 318307 224365
rect 262140 224360 318307 224362
rect 262140 224304 318246 224360
rect 318302 224304 318307 224360
rect 262140 224302 318307 224304
rect 262140 224300 262146 224302
rect 318241 224299 318307 224302
rect 93853 224226 93919 224229
rect 214741 224226 214807 224229
rect 93853 224224 214807 224226
rect 93853 224168 93858 224224
rect 93914 224168 214746 224224
rect 214802 224168 214807 224224
rect 93853 224166 214807 224168
rect 93853 224163 93919 224166
rect 214741 224163 214807 224166
rect 247718 224164 247724 224228
rect 247788 224226 247794 224228
rect 327073 224226 327139 224229
rect 247788 224224 327139 224226
rect 247788 224168 327078 224224
rect 327134 224168 327139 224224
rect 247788 224166 327139 224168
rect 247788 224164 247794 224166
rect 327073 224163 327139 224166
rect 256734 224028 256740 224092
rect 256804 224090 256810 224092
rect 272517 224090 272583 224093
rect 256804 224088 272583 224090
rect 256804 224032 272522 224088
rect 272578 224032 272583 224088
rect 256804 224030 272583 224032
rect 256804 224028 256810 224030
rect 272517 224027 272583 224030
rect 254894 223756 254900 223820
rect 254964 223818 254970 223820
rect 255129 223818 255195 223821
rect 254964 223816 255195 223818
rect 254964 223760 255134 223816
rect 255190 223760 255195 223816
rect 254964 223758 255195 223760
rect 254964 223756 254970 223758
rect 255129 223755 255195 223758
rect 213821 223546 213887 223549
rect 227662 223546 227668 223548
rect 213821 223544 227668 223546
rect 213821 223488 213826 223544
rect 213882 223488 227668 223544
rect 213821 223486 227668 223488
rect 213821 223483 213887 223486
rect 227662 223484 227668 223486
rect 227732 223484 227738 223548
rect 287421 223546 287487 223549
rect 287830 223546 287836 223548
rect 287421 223544 287836 223546
rect 287421 223488 287426 223544
rect 287482 223488 287836 223544
rect 287421 223486 287836 223488
rect 287421 223483 287487 223486
rect 287830 223484 287836 223486
rect 287900 223484 287906 223548
rect 246798 223348 246804 223412
rect 246868 223410 246874 223412
rect 306414 223410 306420 223412
rect 246868 223350 306420 223410
rect 246868 223348 246874 223350
rect 306414 223348 306420 223350
rect 306484 223348 306490 223412
rect 248270 223212 248276 223276
rect 248340 223274 248346 223276
rect 308857 223274 308923 223277
rect 248340 223272 308923 223274
rect 248340 223216 308862 223272
rect 308918 223216 308923 223272
rect 248340 223214 308923 223216
rect 248340 223212 248346 223214
rect 308857 223211 308923 223214
rect 245142 223076 245148 223140
rect 245212 223138 245218 223140
rect 245561 223138 245627 223141
rect 303838 223138 303844 223140
rect 245212 223136 303844 223138
rect 245212 223080 245566 223136
rect 245622 223080 303844 223136
rect 245212 223078 303844 223080
rect 245212 223076 245218 223078
rect 245561 223075 245627 223078
rect 303838 223076 303844 223078
rect 303908 223076 303914 223140
rect 250846 222940 250852 223004
rect 250916 223002 250922 223004
rect 310053 223002 310119 223005
rect 250916 223000 310119 223002
rect 250916 222944 310058 223000
rect 310114 222944 310119 223000
rect 250916 222942 310119 222944
rect 250916 222940 250922 222942
rect 310053 222939 310119 222942
rect 313273 223002 313339 223005
rect 313774 223002 313780 223004
rect 313273 223000 313780 223002
rect 313273 222944 313278 223000
rect 313334 222944 313780 223000
rect 313273 222942 313780 222944
rect 313273 222939 313339 222942
rect 313774 222940 313780 222942
rect 313844 222940 313850 223004
rect 82813 222866 82879 222869
rect 213821 222866 213887 222869
rect 82813 222864 213887 222866
rect 82813 222808 82818 222864
rect 82874 222808 213826 222864
rect 213882 222808 213887 222864
rect 82813 222806 213887 222808
rect 82813 222803 82879 222806
rect 213821 222803 213887 222806
rect 249374 222804 249380 222868
rect 249444 222866 249450 222868
rect 308581 222866 308647 222869
rect 249444 222864 308647 222866
rect 249444 222808 308586 222864
rect 308642 222808 308647 222864
rect 249444 222806 308647 222808
rect 249444 222804 249450 222806
rect 308581 222803 308647 222806
rect 234286 222668 234292 222732
rect 234356 222730 234362 222732
rect 291929 222730 291995 222733
rect 234356 222728 291995 222730
rect 234356 222672 291934 222728
rect 291990 222672 291995 222728
rect 234356 222670 291995 222672
rect 234356 222668 234362 222670
rect 291929 222667 291995 222670
rect 245326 222532 245332 222596
rect 245396 222594 245402 222596
rect 305494 222594 305500 222596
rect 245396 222534 305500 222594
rect 245396 222532 245402 222534
rect 305494 222532 305500 222534
rect 305564 222532 305570 222596
rect 232037 222186 232103 222189
rect 232865 222186 232931 222189
rect 237373 222186 237439 222189
rect 238477 222186 238543 222189
rect 301814 222186 301820 222188
rect 232037 222184 234538 222186
rect 232037 222128 232042 222184
rect 232098 222128 232870 222184
rect 232926 222128 234538 222184
rect 232037 222126 234538 222128
rect 232037 222123 232103 222126
rect 232865 222123 232931 222126
rect 234478 222050 234538 222126
rect 237373 222184 301820 222186
rect 237373 222128 237378 222184
rect 237434 222128 238482 222184
rect 238538 222128 301820 222184
rect 237373 222126 301820 222128
rect 237373 222123 237439 222126
rect 238477 222123 238543 222126
rect 301814 222124 301820 222126
rect 301884 222124 301890 222188
rect 294454 222050 294460 222052
rect 234478 221990 294460 222050
rect 294454 221988 294460 221990
rect 294524 221988 294530 222052
rect 232446 221852 232452 221916
rect 232516 221914 232522 221916
rect 292614 221914 292620 221916
rect 232516 221854 292620 221914
rect 232516 221852 232522 221854
rect 292614 221852 292620 221854
rect 292684 221852 292690 221916
rect 238845 221778 238911 221781
rect 298134 221778 298140 221780
rect 238710 221776 298140 221778
rect 238710 221720 238850 221776
rect 238906 221720 298140 221776
rect 238710 221718 298140 221720
rect 212533 221642 212599 221645
rect 238710 221642 238770 221718
rect 238845 221715 238911 221718
rect 298134 221716 298140 221718
rect 298204 221716 298210 221780
rect 212533 221640 238770 221642
rect 212533 221584 212538 221640
rect 212594 221584 238770 221640
rect 212533 221582 238770 221584
rect 212533 221579 212599 221582
rect 251950 221580 251956 221644
rect 252020 221642 252026 221644
rect 252277 221642 252343 221645
rect 311433 221642 311499 221645
rect 252020 221640 311499 221642
rect 252020 221584 252282 221640
rect 252338 221584 311438 221640
rect 311494 221584 311499 221640
rect 252020 221582 311499 221584
rect 252020 221580 252026 221582
rect 252277 221579 252343 221582
rect 311433 221579 311499 221582
rect 131113 221506 131179 221509
rect 232446 221506 232452 221508
rect 131113 221504 232452 221506
rect 131113 221448 131118 221504
rect 131174 221448 232452 221504
rect 131113 221446 232452 221448
rect 131113 221443 131179 221446
rect 232446 221444 232452 221446
rect 232516 221444 232522 221508
rect 256182 221444 256188 221508
rect 256252 221506 256258 221508
rect 290457 221506 290523 221509
rect 256252 221504 290523 221506
rect 256252 221448 290462 221504
rect 290518 221448 290523 221504
rect 256252 221446 290523 221448
rect 256252 221444 256258 221446
rect 290457 221443 290523 221446
rect 256918 221308 256924 221372
rect 256988 221370 256994 221372
rect 275369 221370 275435 221373
rect 256988 221368 275435 221370
rect 256988 221312 275374 221368
rect 275430 221312 275435 221368
rect 256988 221310 275435 221312
rect 256988 221308 256994 221310
rect 275369 221307 275435 221310
rect 264462 221172 264468 221236
rect 264532 221234 264538 221236
rect 264605 221234 264671 221237
rect 264532 221232 264671 221234
rect 264532 221176 264610 221232
rect 264666 221176 264671 221232
rect 264532 221174 264671 221176
rect 264532 221172 264538 221174
rect 264605 221171 264671 221174
rect 223757 220826 223823 220829
rect 224493 220826 224559 220829
rect 223757 220824 224559 220826
rect 223757 220768 223762 220824
rect 223818 220768 224498 220824
rect 224554 220768 224559 220824
rect 223757 220766 224559 220768
rect 223757 220763 223823 220766
rect 224493 220763 224559 220766
rect 228265 220826 228331 220829
rect 228725 220826 228791 220829
rect 228265 220824 228791 220826
rect 228265 220768 228270 220824
rect 228326 220768 228730 220824
rect 228786 220768 228791 220824
rect 228265 220766 228791 220768
rect 228265 220763 228331 220766
rect 228725 220763 228791 220766
rect 242750 220764 242756 220828
rect 242820 220826 242826 220828
rect 244917 220826 244983 220829
rect 242820 220824 244983 220826
rect 242820 220768 244922 220824
rect 244978 220768 244983 220824
rect 242820 220766 244983 220768
rect 242820 220764 242826 220766
rect 244917 220763 244983 220766
rect 225229 220690 225295 220693
rect 285622 220690 285628 220692
rect 225229 220688 285628 220690
rect 225229 220632 225234 220688
rect 225290 220632 285628 220688
rect 225229 220630 285628 220632
rect 225229 220627 225295 220630
rect 285622 220628 285628 220630
rect 285692 220628 285698 220692
rect 224493 220554 224559 220557
rect 282862 220554 282868 220556
rect 224493 220552 282868 220554
rect 224493 220496 224498 220552
rect 224554 220496 282868 220552
rect 224493 220494 282868 220496
rect 224493 220491 224559 220494
rect 282862 220492 282868 220494
rect 282932 220492 282938 220556
rect 228582 220356 228588 220420
rect 228652 220418 228658 220420
rect 228652 220358 283666 220418
rect 228652 220356 228658 220358
rect 114553 220282 114619 220285
rect 231342 220282 231348 220284
rect 114553 220280 231348 220282
rect 114553 220224 114558 220280
rect 114614 220224 231348 220280
rect 114553 220222 231348 220224
rect 114553 220219 114619 220222
rect 231342 220220 231348 220222
rect 231412 220282 231418 220284
rect 282913 220282 282979 220285
rect 283414 220282 283420 220284
rect 231412 220222 277410 220282
rect 231412 220220 231418 220222
rect 231526 220084 231532 220148
rect 231596 220146 231602 220148
rect 276657 220146 276723 220149
rect 231596 220144 276723 220146
rect 231596 220088 276662 220144
rect 276718 220088 276723 220144
rect 231596 220086 276723 220088
rect 277350 220146 277410 220222
rect 282913 220280 283420 220282
rect 282913 220224 282918 220280
rect 282974 220224 283420 220280
rect 282913 220222 283420 220224
rect 282913 220219 282979 220222
rect 283414 220220 283420 220222
rect 283484 220220 283490 220284
rect 283606 220282 283666 220358
rect 287094 220282 287100 220284
rect 283606 220222 287100 220282
rect 287094 220220 287100 220222
rect 287164 220220 287170 220284
rect 289077 220146 289143 220149
rect 277350 220144 289143 220146
rect 277350 220088 289082 220144
rect 289138 220088 289143 220144
rect 277350 220086 289143 220088
rect 231596 220084 231602 220086
rect 276657 220083 276723 220086
rect 289077 220083 289143 220086
rect 228725 219874 228791 219877
rect 291142 219874 291148 219876
rect 228725 219872 291148 219874
rect 228725 219816 228730 219872
rect 228786 219816 291148 219872
rect 228725 219814 291148 219816
rect 228725 219811 228791 219814
rect 291142 219812 291148 219814
rect 291212 219812 291218 219876
rect 224033 219330 224099 219333
rect 284334 219330 284340 219332
rect 224033 219328 284340 219330
rect 224033 219272 224038 219328
rect 224094 219272 284340 219328
rect 224033 219270 284340 219272
rect 224033 219267 224099 219270
rect 284334 219268 284340 219270
rect 284404 219268 284410 219332
rect 227989 219194 228055 219197
rect 303429 219196 303495 219197
rect 288382 219194 288388 219196
rect 227989 219192 288388 219194
rect 227989 219136 227994 219192
rect 228050 219136 288388 219192
rect 227989 219134 288388 219136
rect 227989 219131 228055 219134
rect 288382 219132 288388 219134
rect 288452 219132 288458 219196
rect 303429 219192 303476 219196
rect 303540 219194 303546 219196
rect 303429 219136 303434 219192
rect 303429 219132 303476 219136
rect 303540 219134 303586 219194
rect 303540 219132 303546 219134
rect 303429 219131 303495 219132
rect 260046 218996 260052 219060
rect 260116 219058 260122 219060
rect 317454 219058 317460 219060
rect 260116 218998 317460 219058
rect 260116 218996 260122 218998
rect 317454 218996 317460 218998
rect 317524 218996 317530 219060
rect 580533 219058 580599 219061
rect 583520 219058 584960 219148
rect 580533 219056 584960 219058
rect 580533 219000 580538 219056
rect 580594 219000 584960 219056
rect 580533 218998 584960 219000
rect 580533 218995 580599 218998
rect 235758 218860 235764 218924
rect 235828 218922 235834 218924
rect 287789 218922 287855 218925
rect 235828 218920 287855 218922
rect 235828 218864 287794 218920
rect 287850 218864 287855 218920
rect 583520 218908 584960 218998
rect 235828 218862 287855 218864
rect 235828 218860 235834 218862
rect 287789 218859 287855 218862
rect 231710 218724 231716 218788
rect 231780 218786 231786 218788
rect 279509 218786 279575 218789
rect 231780 218784 279575 218786
rect 231780 218728 279514 218784
rect 279570 218728 279575 218784
rect 231780 218726 279575 218728
rect 231780 218724 231786 218726
rect 279509 218723 279575 218726
rect 257102 218588 257108 218652
rect 257172 218650 257178 218652
rect 285029 218650 285095 218653
rect 257172 218648 285095 218650
rect 257172 218592 285034 218648
rect 285090 218592 285095 218648
rect 257172 218590 285095 218592
rect 257172 218588 257178 218590
rect 285029 218587 285095 218590
rect 258942 218452 258948 218516
rect 259012 218514 259018 218516
rect 286501 218514 286567 218517
rect 259012 218512 286567 218514
rect 259012 218456 286506 218512
rect 286562 218456 286567 218512
rect 259012 218454 286567 218456
rect 259012 218452 259018 218454
rect 286501 218451 286567 218454
rect 230974 218044 230980 218108
rect 231044 218106 231050 218108
rect 231710 218106 231716 218108
rect 231044 218046 231716 218106
rect 231044 218044 231050 218046
rect 231710 218044 231716 218046
rect 231780 218044 231786 218108
rect 235257 218106 235323 218109
rect 235758 218106 235764 218108
rect 235257 218104 235764 218106
rect 235257 218048 235262 218104
rect 235318 218048 235764 218104
rect 235257 218046 235764 218048
rect 235257 218043 235323 218046
rect 235758 218044 235764 218046
rect 235828 218044 235834 218108
rect 259361 218106 259427 218109
rect 260046 218106 260052 218108
rect 259361 218104 260052 218106
rect 259361 218048 259366 218104
rect 259422 218048 260052 218104
rect 259361 218046 260052 218048
rect 259361 218043 259427 218046
rect 260046 218044 260052 218046
rect 260116 218044 260122 218108
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 243302 214508 243308 214572
rect 243372 214570 243378 214572
rect 280153 214570 280219 214573
rect 281165 214570 281231 214573
rect 243372 214568 281231 214570
rect 243372 214512 280158 214568
rect 280214 214512 281170 214568
rect 281226 214512 281231 214568
rect 243372 214510 281231 214512
rect 243372 214508 243378 214510
rect 280153 214507 280219 214510
rect 281165 214507 281231 214510
rect 281165 213890 281231 213893
rect 303654 213890 303660 213892
rect 281165 213888 303660 213890
rect 281165 213832 281170 213888
rect 281226 213832 303660 213888
rect 281165 213830 303660 213832
rect 281165 213827 281231 213830
rect 303654 213828 303660 213830
rect 303724 213828 303730 213892
rect 69013 213210 69079 213213
rect 228582 213210 228588 213212
rect 69013 213208 228588 213210
rect 69013 213152 69018 213208
rect 69074 213152 228588 213208
rect 69013 213150 228588 213152
rect 69013 213147 69079 213150
rect 228582 213148 228588 213150
rect 228652 213148 228658 213212
rect 246246 213148 246252 213212
rect 246316 213210 246322 213212
rect 304993 213210 305059 213213
rect 246316 213208 305059 213210
rect 246316 213152 304998 213208
rect 305054 213152 305059 213208
rect 246316 213150 305059 213152
rect 246316 213148 246322 213150
rect 304993 213147 305059 213150
rect 244958 211788 244964 211852
rect 245028 211850 245034 211852
rect 289169 211850 289235 211853
rect 245028 211848 289235 211850
rect 245028 211792 289174 211848
rect 289230 211792 289235 211848
rect 245028 211790 289235 211792
rect 245028 211788 245034 211790
rect 289169 211787 289235 211790
rect 292573 208314 292639 208317
rect 304206 208314 304212 208316
rect 292573 208312 304212 208314
rect 292573 208256 292578 208312
rect 292634 208256 304212 208312
rect 292573 208254 304212 208256
rect 292573 208251 292639 208254
rect 304206 208252 304212 208254
rect 304276 208252 304282 208316
rect 142153 207634 142219 207637
rect 233918 207634 233924 207636
rect 142153 207632 233924 207634
rect 142153 207576 142158 207632
rect 142214 207576 233924 207632
rect 142153 207574 233924 207576
rect 142153 207571 142219 207574
rect 233918 207572 233924 207574
rect 233988 207572 233994 207636
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 242382 204852 242388 204916
rect 242452 204914 242458 204916
rect 258073 204914 258139 204917
rect 242452 204912 258139 204914
rect 242452 204856 258078 204912
rect 258134 204856 258139 204912
rect 242452 204854 258139 204856
rect 242452 204852 242458 204854
rect 258073 204851 258139 204854
rect 104893 203554 104959 203557
rect 231158 203554 231164 203556
rect 104893 203552 231164 203554
rect 104893 203496 104898 203552
rect 104954 203496 231164 203552
rect 104893 203494 231164 203496
rect 104893 203491 104959 203494
rect 231158 203492 231164 203494
rect 231228 203492 231234 203556
rect 250846 202132 250852 202196
rect 250916 202194 250922 202196
rect 354673 202194 354739 202197
rect 250916 202192 354739 202194
rect 250916 202136 354678 202192
rect 354734 202136 354739 202192
rect 250916 202134 354739 202136
rect 250916 202132 250922 202134
rect 354673 202131 354739 202134
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 62113 200698 62179 200701
rect 227294 200698 227300 200700
rect 62113 200696 227300 200698
rect 62113 200640 62118 200696
rect 62174 200640 227300 200696
rect 62113 200638 227300 200640
rect 62113 200635 62179 200638
rect 227294 200636 227300 200638
rect 227364 200636 227370 200700
rect 242566 200636 242572 200700
rect 242636 200698 242642 200700
rect 260097 200698 260163 200701
rect 242636 200696 260163 200698
rect 242636 200640 260102 200696
rect 260158 200640 260163 200696
rect 242636 200638 260163 200640
rect 242636 200636 242642 200638
rect 260097 200635 260163 200638
rect 226977 199474 227043 199477
rect 238886 199474 238892 199476
rect 226977 199472 238892 199474
rect 226977 199416 226982 199472
rect 227038 199416 238892 199472
rect 226977 199414 238892 199416
rect 226977 199411 227043 199414
rect 238886 199412 238892 199414
rect 238956 199412 238962 199476
rect 102133 199338 102199 199341
rect 230054 199338 230060 199340
rect 102133 199336 230060 199338
rect 102133 199280 102138 199336
rect 102194 199280 230060 199336
rect 102133 199278 230060 199280
rect 102133 199275 102199 199278
rect 230054 199276 230060 199278
rect 230124 199276 230130 199340
rect 247534 199276 247540 199340
rect 247604 199338 247610 199340
rect 324957 199338 325023 199341
rect 247604 199336 325023 199338
rect 247604 199280 324962 199336
rect 325018 199280 325023 199336
rect 247604 199278 325023 199280
rect 247604 199276 247610 199278
rect 324957 199275 325023 199278
rect 249374 197916 249380 197980
rect 249444 197978 249450 197980
rect 336733 197978 336799 197981
rect 249444 197976 336799 197978
rect 249444 197920 336738 197976
rect 336794 197920 336799 197976
rect 249444 197918 336799 197920
rect 249444 197916 249450 197918
rect 336733 197915 336799 197918
rect 66253 196618 66319 196621
rect 226926 196618 226932 196620
rect 66253 196616 226932 196618
rect 66253 196560 66258 196616
rect 66314 196560 226932 196616
rect 66253 196558 226932 196560
rect 66253 196555 66319 196558
rect 226926 196556 226932 196558
rect 226996 196556 227002 196620
rect 143625 193898 143691 193901
rect 233734 193898 233740 193900
rect 143625 193896 233740 193898
rect 143625 193840 143630 193896
rect 143686 193840 233740 193896
rect 143625 193838 233740 193840
rect 143625 193835 143691 193838
rect 233734 193836 233740 193838
rect 233804 193836 233810 193900
rect 246062 192476 246068 192540
rect 246132 192538 246138 192540
rect 311157 192538 311223 192541
rect 246132 192536 311223 192538
rect 246132 192480 311162 192536
rect 311218 192480 311223 192536
rect 246132 192478 311223 192480
rect 246132 192476 246138 192478
rect 311157 192475 311223 192478
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 262990 190980 262996 191044
rect 263060 191042 263066 191044
rect 514845 191042 514911 191045
rect 263060 191040 514911 191042
rect 263060 190984 514850 191040
rect 514906 190984 514911 191040
rect 263060 190982 514911 190984
rect 263060 190980 263066 190982
rect 514845 190979 514911 190982
rect 263174 189620 263180 189684
rect 263244 189682 263250 189684
rect 517513 189682 517579 189685
rect 263244 189680 517579 189682
rect 263244 189624 517518 189680
rect 517574 189624 517579 189680
rect 263244 189622 517579 189624
rect 263244 189620 263250 189622
rect 517513 189619 517579 189622
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 144913 188322 144979 188325
rect 233550 188322 233556 188324
rect 144913 188320 233556 188322
rect 144913 188264 144918 188320
rect 144974 188264 233556 188320
rect 144913 188262 233556 188264
rect 144913 188259 144979 188262
rect 233550 188260 233556 188262
rect 233620 188260 233626 188324
rect 245326 188260 245332 188324
rect 245396 188322 245402 188324
rect 298093 188322 298159 188325
rect 245396 188320 298159 188322
rect 245396 188264 298098 188320
rect 298154 188264 298159 188320
rect 245396 188262 298159 188264
rect 245396 188260 245402 188262
rect 298093 188259 298159 188262
rect 247350 186900 247356 186964
rect 247420 186962 247426 186964
rect 329833 186962 329899 186965
rect 247420 186960 329899 186962
rect 247420 186904 329838 186960
rect 329894 186904 329899 186960
rect 247420 186902 329899 186904
rect 247420 186900 247426 186902
rect 329833 186899 329899 186902
rect 118785 182882 118851 182885
rect 230974 182882 230980 182884
rect 118785 182880 230980 182882
rect 118785 182824 118790 182880
rect 118846 182824 230980 182880
rect 118785 182822 230980 182824
rect 118785 182819 118851 182822
rect 230974 182820 230980 182822
rect 231044 182820 231050 182884
rect 263726 182820 263732 182884
rect 263796 182882 263802 182884
rect 546493 182882 546559 182885
rect 263796 182880 546559 182882
rect 263796 182824 546498 182880
rect 546554 182824 546559 182880
rect 263796 182822 546559 182824
rect 263796 182820 263802 182822
rect 546493 182819 546559 182822
rect 579705 179210 579771 179213
rect 583520 179210 584960 179300
rect 579705 179208 584960 179210
rect 579705 179152 579710 179208
rect 579766 179152 584960 179208
rect 579705 179150 584960 179152
rect 579705 179147 579771 179150
rect 583520 179060 584960 179150
rect 249006 178604 249012 178668
rect 249076 178666 249082 178668
rect 350533 178666 350599 178669
rect 249076 178664 350599 178666
rect 249076 178608 350538 178664
rect 350594 178608 350599 178664
rect 249076 178606 350599 178608
rect 249076 178604 249082 178606
rect 350533 178603 350599 178606
rect -960 175796 480 176036
rect 256734 168948 256740 169012
rect 256804 169010 256810 169012
rect 447133 169010 447199 169013
rect 256804 169008 447199 169010
rect 256804 168952 447138 169008
rect 447194 168952 447199 169008
rect 256804 168950 447199 168952
rect 256804 168948 256810 168950
rect 447133 168947 447199 168950
rect 249190 167588 249196 167652
rect 249260 167650 249266 167652
rect 347773 167650 347839 167653
rect 249260 167648 347839 167650
rect 249260 167592 347778 167648
rect 347834 167592 347839 167648
rect 249260 167590 347839 167592
rect 249260 167588 249266 167590
rect 347773 167587 347839 167590
rect 245510 166228 245516 166292
rect 245580 166290 245586 166292
rect 293953 166290 294019 166293
rect 245580 166288 294019 166290
rect 245580 166232 293958 166288
rect 294014 166232 294019 166288
rect 245580 166230 294019 166232
rect 245580 166228 245586 166230
rect 293953 166227 294019 166230
rect 580625 165882 580691 165885
rect 583520 165882 584960 165972
rect 580625 165880 584960 165882
rect 580625 165824 580630 165880
rect 580686 165824 584960 165880
rect 580625 165822 584960 165824
rect 580625 165819 580691 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 226333 156634 226399 156637
rect 239438 156634 239444 156636
rect 226333 156632 239444 156634
rect 226333 156576 226338 156632
rect 226394 156576 239444 156632
rect 226333 156574 239444 156576
rect 226333 156571 226399 156574
rect 239438 156572 239444 156574
rect 239508 156572 239514 156636
rect 255078 156572 255084 156636
rect 255148 156634 255154 156636
rect 418153 156634 418219 156637
rect 255148 156632 418219 156634
rect 255148 156576 418158 156632
rect 418214 156576 418219 156632
rect 255148 156574 418219 156576
rect 255148 156572 255154 156574
rect 418153 156571 418219 156574
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 246798 152356 246804 152420
rect 246868 152418 246874 152420
rect 316125 152418 316191 152421
rect 246868 152416 316191 152418
rect 246868 152360 316130 152416
rect 316186 152360 316191 152416
rect 246868 152358 316191 152360
rect 246868 152356 246874 152358
rect 316125 152355 316191 152358
rect 256918 150996 256924 151060
rect 256988 151058 256994 151060
rect 449893 151058 449959 151061
rect 256988 151056 449959 151058
rect 256988 151000 449898 151056
rect 449954 151000 449959 151056
rect 256988 150998 449959 151000
rect 256988 150996 256994 150998
rect 449893 150995 449959 150998
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 258942 146916 258948 146980
rect 259012 146978 259018 146980
rect 471973 146978 472039 146981
rect 259012 146976 472039 146978
rect 259012 146920 471978 146976
rect 472034 146920 472039 146976
rect 259012 146918 472039 146920
rect 259012 146916 259018 146918
rect 471973 146915 472039 146918
rect 242198 141340 242204 141404
rect 242268 141402 242274 141404
rect 262213 141402 262279 141405
rect 242268 141400 262279 141402
rect 242268 141344 262218 141400
rect 262274 141344 262279 141400
rect 242268 141342 262279 141344
rect 242268 141340 242274 141342
rect 262213 141339 262279 141342
rect 580349 139362 580415 139365
rect 583520 139362 584960 139452
rect 580349 139360 584960 139362
rect 580349 139304 580354 139360
rect 580410 139304 584960 139360
rect 580349 139302 584960 139304
rect 580349 139299 580415 139302
rect 583520 139212 584960 139302
rect 251030 138620 251036 138684
rect 251100 138682 251106 138684
rect 365805 138682 365871 138685
rect 251100 138680 365871 138682
rect 251100 138624 365810 138680
rect 365866 138624 365871 138680
rect 251100 138622 365871 138624
rect 251100 138620 251106 138622
rect 365805 138619 365871 138622
rect -960 136778 480 136868
rect 2865 136778 2931 136781
rect -960 136776 2931 136778
rect -960 136720 2870 136776
rect 2926 136720 2931 136776
rect -960 136718 2931 136720
rect -960 136628 480 136718
rect 2865 136715 2931 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 269614 125564 269620 125628
rect 269684 125626 269690 125628
rect 583526 125626 583586 125838
rect 269684 125566 583586 125626
rect 269684 125564 269690 125566
rect -960 123572 480 123812
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580441 86186 580507 86189
rect 583520 86186 584960 86276
rect 580441 86184 584960 86186
rect 580441 86128 580446 86184
rect 580502 86128 584960 86184
rect 580441 86126 584960 86128
rect 580441 86123 580507 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580349 46338 580415 46341
rect 583520 46338 584960 46428
rect 580349 46336 584960 46338
rect 580349 46280 580354 46336
rect 580410 46280 584960 46336
rect 580349 46278 584960 46280
rect 580349 46275 580415 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 281390 31724 281396 31788
rect 281460 31786 281466 31788
rect 583526 31786 583586 32950
rect 281460 31726 583586 31786
rect 281460 31724 281466 31726
rect 259126 25468 259132 25532
rect 259196 25530 259202 25532
rect 474733 25530 474799 25533
rect 259196 25528 474799 25530
rect 259196 25472 474738 25528
rect 474794 25472 474799 25528
rect 259196 25470 474799 25472
rect 259196 25468 259202 25470
rect 474733 25467 474799 25470
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 257102 15812 257108 15876
rect 257172 15874 257178 15876
rect 456885 15874 456951 15877
rect 257172 15872 456951 15874
rect 257172 15816 456890 15872
rect 456946 15816 456951 15872
rect 257172 15814 456951 15816
rect 257172 15812 257178 15814
rect 456885 15811 456951 15814
rect 262622 10236 262628 10300
rect 262692 10298 262698 10300
rect 528553 10298 528619 10301
rect 262692 10296 528619 10298
rect 262692 10240 528558 10296
rect 528614 10240 528619 10296
rect 262692 10238 528619 10240
rect 262692 10236 262698 10238
rect 528553 10235 528619 10238
rect 252686 6836 252692 6900
rect 252756 6898 252762 6900
rect 401317 6898 401383 6901
rect 252756 6896 401383 6898
rect 252756 6840 401322 6896
rect 401378 6840 401383 6896
rect 252756 6838 401383 6840
rect 252756 6836 252762 6838
rect 401317 6835 401383 6838
rect 253238 6700 253244 6764
rect 253308 6762 253314 6764
rect 404813 6762 404879 6765
rect 253308 6760 404879 6762
rect 253308 6704 404818 6760
rect 404874 6704 404879 6760
rect 253308 6702 404879 6704
rect 253308 6700 253314 6702
rect 404813 6699 404879 6702
rect -960 6490 480 6580
rect 256182 6564 256188 6628
rect 256252 6626 256258 6628
rect 426157 6626 426223 6629
rect 256252 6624 426223 6626
rect 256252 6568 426162 6624
rect 426218 6568 426223 6624
rect 256252 6566 426223 6568
rect 256252 6564 256258 6566
rect 426157 6563 426223 6566
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 256366 6428 256372 6492
rect 256436 6490 256442 6492
rect 436645 6490 436711 6493
rect 256436 6488 436711 6490
rect 256436 6432 436650 6488
rect 436706 6432 436711 6488
rect 583520 6476 584960 6566
rect 256436 6430 436711 6432
rect 256436 6428 256442 6430
rect 436645 6427 436711 6430
rect 255998 6292 256004 6356
rect 256068 6354 256074 6356
rect 440325 6354 440391 6357
rect 256068 6352 440391 6354
rect 256068 6296 440330 6352
rect 440386 6296 440391 6352
rect 256068 6294 440391 6296
rect 256068 6292 256074 6294
rect 440325 6291 440391 6294
rect 259310 6156 259316 6220
rect 259380 6218 259386 6220
rect 465165 6218 465231 6221
rect 259380 6216 465231 6218
rect 259380 6160 465170 6216
rect 465226 6160 465231 6216
rect 259380 6158 465231 6160
rect 259380 6156 259386 6158
rect 465165 6155 465231 6158
rect 248270 6020 248276 6084
rect 248340 6082 248346 6084
rect 333881 6082 333947 6085
rect 248340 6080 333947 6082
rect 248340 6024 333886 6080
rect 333942 6024 333947 6080
rect 248340 6022 333947 6024
rect 248340 6020 248346 6022
rect 333881 6019 333947 6022
rect 251582 3572 251588 3636
rect 251652 3634 251658 3636
rect 379973 3634 380039 3637
rect 251652 3632 380039 3634
rect 251652 3576 379978 3632
rect 380034 3576 380039 3632
rect 251652 3574 380039 3576
rect 251652 3572 251658 3574
rect 379973 3571 380039 3574
rect 252134 3436 252140 3500
rect 252204 3498 252210 3500
rect 383561 3498 383627 3501
rect 252204 3496 383627 3498
rect 252204 3440 383566 3496
rect 383622 3440 383627 3496
rect 252204 3438 383627 3440
rect 252204 3436 252210 3438
rect 383561 3435 383627 3438
rect 260598 3300 260604 3364
rect 260668 3362 260674 3364
rect 486417 3362 486483 3365
rect 260668 3360 486483 3362
rect 260668 3304 486422 3360
rect 486478 3304 486483 3360
rect 260668 3302 486483 3304
rect 260668 3300 260674 3302
rect 486417 3299 486483 3302
<< via3 >>
rect 309180 403548 309244 403612
rect 313412 389812 313476 389876
rect 305500 386276 305564 386340
rect 316724 385596 316788 385660
rect 314700 381516 314764 381580
rect 313228 380156 313292 380220
rect 309364 378660 309428 378724
rect 306420 377300 306484 377364
rect 277900 375668 277964 375732
rect 275324 375532 275388 375596
rect 275140 375396 275204 375460
rect 307708 374580 307772 374644
rect 278084 374172 278148 374236
rect 307524 372540 307588 372604
rect 309364 372540 309428 372604
rect 285628 371860 285692 371924
rect 296484 371316 296548 371380
rect 288020 369880 288084 369884
rect 288020 369824 288024 369880
rect 288024 369824 288080 369880
rect 288080 369824 288084 369880
rect 288020 369820 288084 369824
rect 308076 369684 308140 369748
rect 309364 369744 309428 369748
rect 309364 369688 309368 369744
rect 309368 369688 309424 369744
rect 309424 369688 309428 369744
rect 309364 369684 309428 369688
rect 311572 369684 311636 369748
rect 283788 369548 283852 369612
rect 283052 369412 283116 369476
rect 283972 369412 284036 369476
rect 284892 369472 284956 369476
rect 284892 369416 284942 369472
rect 284942 369416 284956 369472
rect 284892 369412 284956 369416
rect 287284 369412 287348 369476
rect 282684 369140 282748 369204
rect 299980 369412 300044 369476
rect 302740 369412 302804 369476
rect 303660 369412 303724 369476
rect 305500 369472 305564 369476
rect 305500 369416 305514 369472
rect 305514 369416 305564 369472
rect 305500 369412 305564 369416
rect 306420 369412 306484 369476
rect 309916 369472 309980 369476
rect 309916 369416 309930 369472
rect 309930 369416 309980 369472
rect 309916 369412 309980 369416
rect 311020 369472 311084 369476
rect 311020 369416 311034 369472
rect 311034 369416 311084 369472
rect 311020 369412 311084 369416
rect 311756 369412 311820 369476
rect 307524 369276 307588 369340
rect 310100 369336 310164 369340
rect 310100 369280 310104 369336
rect 310104 369280 310160 369336
rect 310160 369280 310164 369336
rect 310100 369276 310164 369280
rect 313228 369412 313292 369476
rect 314700 369412 314764 369476
rect 320220 369412 320284 369476
rect 322796 369412 322860 369476
rect 313412 369336 313476 369340
rect 313412 369280 313416 369336
rect 313416 369280 313472 369336
rect 313472 369280 313476 369336
rect 313412 369276 313476 369280
rect 316724 369336 316788 369340
rect 316724 369280 316728 369336
rect 316728 369280 316784 369336
rect 316784 369280 316788 369336
rect 316724 369276 316788 369280
rect 310100 368596 310164 368660
rect 285628 367780 285692 367844
rect 288020 367644 288084 367708
rect 284892 367508 284956 367572
rect 283788 362204 283852 362268
rect 281396 360164 281460 360228
rect 283972 360164 284036 360228
rect 283972 321812 284036 321876
rect 293172 321676 293236 321740
rect 288020 321540 288084 321604
rect 319300 321540 319364 321604
rect 306420 321268 306484 321332
rect 317460 321268 317524 321332
rect 307708 321132 307772 321196
rect 310652 321132 310716 321196
rect 314700 321132 314764 321196
rect 303660 320996 303724 321060
rect 313412 320860 313476 320924
rect 325372 320860 325436 320924
rect 287284 320724 287348 320788
rect 288020 320784 288084 320788
rect 288020 320728 288024 320784
rect 288024 320728 288080 320784
rect 288080 320728 288084 320784
rect 288020 320724 288084 320728
rect 291884 320724 291948 320788
rect 292620 320724 292684 320788
rect 294460 320724 294524 320788
rect 295748 320724 295812 320788
rect 299244 320724 299308 320788
rect 322244 320724 322308 320788
rect 299980 320588 300044 320652
rect 312860 320588 312924 320652
rect 313412 320588 313476 320652
rect 313228 320452 313292 320516
rect 317460 320452 317524 320516
rect 318564 320452 318628 320516
rect 319116 320452 319180 320516
rect 325372 320452 325436 320516
rect 283420 320316 283484 320380
rect 283788 320376 283852 320380
rect 283788 320320 283792 320376
rect 283792 320320 283848 320376
rect 283848 320320 283852 320376
rect 283788 320316 283852 320320
rect 288940 320316 289004 320380
rect 290780 320316 290844 320380
rect 292804 320316 292868 320380
rect 299612 320316 299676 320380
rect 299796 320316 299860 320380
rect 307708 320316 307772 320380
rect 313228 320376 313292 320380
rect 313228 320320 313232 320376
rect 313232 320320 313288 320376
rect 313288 320320 313292 320376
rect 285628 320180 285692 320244
rect 287836 320180 287900 320244
rect 288756 320180 288820 320244
rect 289492 320180 289556 320244
rect 290964 320240 291028 320244
rect 290964 320184 290968 320240
rect 290968 320184 291024 320240
rect 291024 320184 291028 320240
rect 290964 320180 291028 320184
rect 291332 320240 291396 320244
rect 291332 320184 291336 320240
rect 291336 320184 291392 320240
rect 291392 320184 291396 320240
rect 291332 320180 291396 320184
rect 293356 320180 293420 320244
rect 294644 320180 294708 320244
rect 294828 320180 294892 320244
rect 297956 320180 298020 320244
rect 283236 320044 283300 320108
rect 284340 320044 284404 320108
rect 285812 320044 285876 320108
rect 286732 320044 286796 320108
rect 287652 320104 287716 320108
rect 287652 320048 287656 320104
rect 287656 320048 287712 320104
rect 287712 320048 287716 320104
rect 287652 320044 287716 320048
rect 288020 320044 288084 320108
rect 288204 320044 288268 320108
rect 288572 320044 288636 320108
rect 289124 320044 289188 320108
rect 290596 320044 290660 320108
rect 291516 320104 291580 320108
rect 291516 320048 291520 320104
rect 291520 320048 291576 320104
rect 291576 320048 291580 320104
rect 291516 320044 291580 320048
rect 291700 320104 291764 320108
rect 291700 320048 291704 320104
rect 291704 320048 291760 320104
rect 291760 320048 291764 320104
rect 291700 320044 291764 320048
rect 292068 320044 292132 320108
rect 292988 320044 293052 320108
rect 294276 320104 294340 320108
rect 294276 320048 294280 320104
rect 294280 320048 294336 320104
rect 294336 320048 294340 320104
rect 294276 320044 294340 320048
rect 295012 320104 295076 320108
rect 295012 320048 295016 320104
rect 295016 320048 295072 320104
rect 295072 320048 295076 320104
rect 295012 320044 295076 320048
rect 295564 320104 295628 320108
rect 295564 320048 295568 320104
rect 295568 320048 295624 320104
rect 295624 320048 295628 320104
rect 295564 320044 295628 320048
rect 295932 320104 295996 320108
rect 295932 320048 295936 320104
rect 295936 320048 295992 320104
rect 295992 320048 295996 320104
rect 295932 320044 295996 320048
rect 297036 320044 297100 320108
rect 283420 319908 283484 319972
rect 285444 319908 285508 319972
rect 289308 319908 289372 319972
rect 291148 319908 291212 319972
rect 292436 319908 292500 319972
rect 295380 319908 295444 319972
rect 296852 319908 296916 319972
rect 299060 320180 299124 320244
rect 300532 320180 300596 320244
rect 303660 320180 303724 320244
rect 308076 320180 308140 320244
rect 310284 320180 310348 320244
rect 310836 320240 310900 320244
rect 310836 320184 310840 320240
rect 310840 320184 310896 320240
rect 310896 320184 310900 320240
rect 310836 320180 310900 320184
rect 311388 320180 311452 320244
rect 298324 320044 298388 320108
rect 299428 320044 299492 320108
rect 299980 320044 300044 320108
rect 300716 320104 300780 320108
rect 300716 320048 300720 320104
rect 300720 320048 300776 320104
rect 300776 320048 300780 320104
rect 300716 320044 300780 320048
rect 301820 320044 301884 320108
rect 302372 320044 302436 320108
rect 303844 320104 303908 320108
rect 303844 320048 303848 320104
rect 303848 320048 303904 320104
rect 303904 320048 303908 320104
rect 303844 320044 303908 320048
rect 304396 320104 304460 320108
rect 304396 320048 304400 320104
rect 304400 320048 304456 320104
rect 304456 320048 304460 320104
rect 304396 320044 304460 320048
rect 305684 320044 305748 320108
rect 306052 320104 306116 320108
rect 306052 320048 306056 320104
rect 306056 320048 306112 320104
rect 306112 320048 306116 320104
rect 306052 320044 306116 320048
rect 306236 320104 306300 320108
rect 306236 320048 306240 320104
rect 306240 320048 306296 320104
rect 306296 320048 306300 320104
rect 306236 320044 306300 320048
rect 306604 320044 306668 320108
rect 307156 320104 307220 320108
rect 307156 320048 307160 320104
rect 307160 320048 307216 320104
rect 307216 320048 307220 320104
rect 307156 320044 307220 320048
rect 307340 320044 307404 320108
rect 307892 320044 307956 320108
rect 309548 320044 309612 320108
rect 309916 320044 309980 320108
rect 310468 320104 310532 320108
rect 310468 320048 310472 320104
rect 310472 320048 310528 320104
rect 310528 320048 310532 320104
rect 310468 320044 310532 320048
rect 311204 320044 311268 320108
rect 313228 320316 313292 320320
rect 317092 320376 317156 320380
rect 317092 320320 317096 320376
rect 317096 320320 317152 320376
rect 317152 320320 317156 320376
rect 317092 320316 317156 320320
rect 318748 320376 318812 320380
rect 318748 320320 318752 320376
rect 318752 320320 318808 320376
rect 318808 320320 318812 320376
rect 318748 320316 318812 320320
rect 323164 320376 323228 320380
rect 323164 320320 323168 320376
rect 323168 320320 323224 320376
rect 323224 320320 323228 320376
rect 306972 319908 307036 319972
rect 310652 319908 310716 319972
rect 306972 319500 307036 319564
rect 307524 319560 307588 319564
rect 307524 319504 307538 319560
rect 307538 319504 307588 319560
rect 307524 319500 307588 319504
rect 307708 319500 307772 319564
rect 309548 319560 309612 319564
rect 309548 319504 309562 319560
rect 309562 319504 309612 319560
rect 309548 319500 309612 319504
rect 311020 319500 311084 319564
rect 311572 319500 311636 319564
rect 283052 319228 283116 319292
rect 283972 319288 284036 319292
rect 283972 319232 284022 319288
rect 284022 319232 284036 319288
rect 283972 319228 284036 319232
rect 285444 319288 285508 319292
rect 285444 319232 285494 319288
rect 285494 319232 285508 319288
rect 285444 319228 285508 319232
rect 287652 319228 287716 319292
rect 289308 319228 289372 319292
rect 290596 319228 290660 319292
rect 290964 319228 291028 319292
rect 291516 319228 291580 319292
rect 293172 319424 293236 319428
rect 293172 319368 293222 319424
rect 293222 319368 293236 319424
rect 293172 319364 293236 319368
rect 294828 319364 294892 319428
rect 296484 319364 296548 319428
rect 299980 319364 300044 319428
rect 300716 319364 300780 319428
rect 301820 319364 301884 319428
rect 302924 319364 302988 319428
rect 304396 319364 304460 319428
rect 306052 319364 306116 319428
rect 306236 319424 306300 319428
rect 306236 319368 306286 319424
rect 306286 319368 306300 319424
rect 306236 319364 306300 319368
rect 306604 319364 306668 319428
rect 308076 319364 308140 319428
rect 310100 319364 310164 319428
rect 311756 319364 311820 319428
rect 314332 320240 314396 320244
rect 314332 320184 314336 320240
rect 314336 320184 314392 320240
rect 314392 320184 314396 320240
rect 314332 320180 314396 320184
rect 314516 320180 314580 320244
rect 316540 320240 316604 320244
rect 316540 320184 316544 320240
rect 316544 320184 316600 320240
rect 316600 320184 316604 320240
rect 316540 320180 316604 320184
rect 314332 319636 314396 319700
rect 313412 319500 313476 319564
rect 316908 320044 316972 320108
rect 318380 320044 318444 320108
rect 316908 319500 316972 319564
rect 316724 319364 316788 319428
rect 319300 320180 319364 320244
rect 319668 320180 319732 320244
rect 323164 320316 323228 320320
rect 321692 320180 321756 320244
rect 322060 320240 322124 320244
rect 322060 320184 322064 320240
rect 322064 320184 322120 320240
rect 322120 320184 322124 320240
rect 322060 320180 322124 320184
rect 324084 320180 324148 320244
rect 323348 320044 323412 320108
rect 323900 320044 323964 320108
rect 322796 319636 322860 319700
rect 322244 319500 322308 319564
rect 323164 319500 323228 319564
rect 318380 319364 318444 319428
rect 319668 319424 319732 319428
rect 319668 319368 319682 319424
rect 319682 319368 319732 319424
rect 319668 319364 319732 319368
rect 305500 319228 305564 319292
rect 307156 319228 307220 319292
rect 309732 319228 309796 319292
rect 309916 319228 309980 319292
rect 310836 319228 310900 319292
rect 311388 319288 311452 319292
rect 311388 319232 311402 319288
rect 311402 319232 311452 319288
rect 311388 319228 311452 319232
rect 320220 319228 320284 319292
rect 323348 319364 323412 319428
rect 323900 319424 323964 319428
rect 323900 319368 323950 319424
rect 323950 319368 323964 319424
rect 323900 319364 323964 319368
rect 324084 319092 324148 319156
rect 246804 318956 246868 319020
rect 310284 318956 310348 319020
rect 311204 318956 311268 319020
rect 313228 318956 313292 319020
rect 316540 318956 316604 319020
rect 319116 319016 319180 319020
rect 319116 318960 319130 319016
rect 319130 318960 319180 319016
rect 319116 318956 319180 318960
rect 232268 318820 232332 318884
rect 292068 318820 292132 318884
rect 293356 318820 293420 318884
rect 294460 318820 294524 318884
rect 295012 318820 295076 318884
rect 295932 318820 295996 318884
rect 296668 318880 296732 318884
rect 296668 318824 296718 318880
rect 296718 318824 296732 318880
rect 296668 318820 296732 318824
rect 296852 318820 296916 318884
rect 299244 318820 299308 318884
rect 299796 318820 299860 318884
rect 300532 318820 300596 318884
rect 305684 318820 305748 318884
rect 312860 318820 312924 318884
rect 321692 318820 321756 318884
rect 286732 318744 286796 318748
rect 286732 318688 286746 318744
rect 286746 318688 286796 318744
rect 286732 318684 286796 318688
rect 287100 318684 287164 318748
rect 288020 318744 288084 318748
rect 288020 318688 288034 318744
rect 288034 318688 288084 318744
rect 288020 318684 288084 318688
rect 288204 318684 288268 318748
rect 288756 318684 288820 318748
rect 289492 318684 289556 318748
rect 291148 318684 291212 318748
rect 220676 318548 220740 318612
rect 282868 318548 282932 318612
rect 298140 318684 298204 318748
rect 299060 318684 299124 318748
rect 302004 318684 302068 318748
rect 304396 318684 304460 318748
rect 307340 318684 307404 318748
rect 310100 318684 310164 318748
rect 314516 318684 314580 318748
rect 295932 318548 295996 318612
rect 317092 318548 317156 318612
rect 292620 318412 292684 318476
rect 297956 318412 298020 318476
rect 307892 318412 307956 318476
rect 283604 318276 283668 318340
rect 292804 318276 292868 318340
rect 299980 318276 300044 318340
rect 303476 318276 303540 318340
rect 282868 318140 282932 318204
rect 291148 318140 291212 318204
rect 292436 318140 292500 318204
rect 303844 318140 303908 318204
rect 291700 318004 291764 318068
rect 283788 317868 283852 317932
rect 285628 317868 285692 317932
rect 291884 317868 291948 317932
rect 294828 317928 294892 317932
rect 294828 317872 294842 317928
rect 294842 317872 294892 317928
rect 294828 317868 294892 317872
rect 298508 317868 298572 317932
rect 302740 317868 302804 317932
rect 306236 317868 306300 317932
rect 319300 317868 319364 317932
rect 302924 317732 302988 317796
rect 306052 317732 306116 317796
rect 314148 317732 314212 317796
rect 318012 317732 318076 317796
rect 318748 317732 318812 317796
rect 284524 317596 284588 317660
rect 285996 317596 286060 317660
rect 291332 317596 291396 317660
rect 294460 317596 294524 317660
rect 303844 317596 303908 317660
rect 305684 317596 305748 317660
rect 306604 317596 306668 317660
rect 285628 317460 285692 317524
rect 287284 317460 287348 317524
rect 287468 317460 287532 317524
rect 288388 317460 288452 317524
rect 291332 317520 291396 317524
rect 291332 317464 291346 317520
rect 291346 317464 291396 317520
rect 291332 317460 291396 317464
rect 291516 317520 291580 317524
rect 291516 317464 291566 317520
rect 291566 317464 291580 317520
rect 291516 317460 291580 317464
rect 292620 317520 292684 317524
rect 292620 317464 292670 317520
rect 292670 317464 292684 317520
rect 292620 317460 292684 317464
rect 295564 317460 295628 317524
rect 299612 317460 299676 317524
rect 301820 317460 301884 317524
rect 304212 317460 304276 317524
rect 305500 317520 305564 317524
rect 305500 317464 305550 317520
rect 305550 317464 305564 317520
rect 305500 317460 305564 317464
rect 306420 317460 306484 317524
rect 311756 317520 311820 317524
rect 311756 317464 311770 317520
rect 311770 317464 311820 317520
rect 311756 317460 311820 317464
rect 313780 317460 313844 317524
rect 317460 317460 317524 317524
rect 328316 317460 328380 317524
rect 226748 317052 226812 317116
rect 299428 315828 299492 315892
rect 232084 315692 232148 315756
rect 253428 315556 253492 315620
rect 223436 315420 223500 315484
rect 243492 315420 243556 315484
rect 294276 315284 294340 315348
rect 299612 315148 299676 315212
rect 294828 315012 294892 315076
rect 314148 315072 314212 315076
rect 314148 315016 314162 315072
rect 314162 315016 314212 315072
rect 314148 315012 314212 315016
rect 222700 314604 222764 314668
rect 310468 314876 310532 314940
rect 311020 314740 311084 314804
rect 285812 314468 285876 314532
rect 289124 314332 289188 314396
rect 295380 314196 295444 314260
rect 296668 314060 296732 314124
rect 297036 313924 297100 313988
rect 241284 312972 241348 313036
rect 238156 312836 238220 312900
rect 238340 312700 238404 312764
rect 238708 312564 238772 312628
rect 298508 312428 298572 312492
rect 242204 312292 242268 312356
rect 243308 312156 243372 312220
rect 288572 312020 288636 312084
rect 292988 312020 293052 312084
rect 311756 312020 311820 312084
rect 322060 311884 322124 311948
rect 249380 311748 249444 311812
rect 247724 311612 247788 311676
rect 249564 311476 249628 311540
rect 246436 311340 246500 311404
rect 248092 311204 248156 311268
rect 249196 311068 249260 311132
rect 234476 310932 234540 310996
rect 288940 310388 289004 310452
rect 254716 310252 254780 310316
rect 253244 310116 253308 310180
rect 253060 309980 253124 310044
rect 285996 309844 286060 309908
rect 290596 309708 290660 309772
rect 291516 309572 291580 309636
rect 252140 309436 252204 309500
rect 287468 309300 287532 309364
rect 230980 308620 231044 308684
rect 259316 308484 259380 308548
rect 259132 308348 259196 308412
rect 245516 307668 245580 307732
rect 302924 307668 302988 307732
rect 230244 307532 230308 307596
rect 223068 307396 223132 307460
rect 230060 307260 230124 307324
rect 284524 307124 284588 307188
rect 295748 307124 295812 307188
rect 298324 306988 298388 307052
rect 238156 306852 238220 306916
rect 238524 306852 238588 306916
rect 238892 306308 238956 306372
rect 240916 305628 240980 305692
rect 228220 304268 228284 304332
rect 287284 304268 287348 304332
rect 227852 304132 227916 304196
rect 318564 304056 318628 304060
rect 318564 304000 318614 304056
rect 318614 304000 318628 304056
rect 318564 303996 318628 304000
rect 228036 302772 228100 302836
rect 327580 302228 327644 302292
rect 242020 300324 242084 300388
rect 251588 300188 251652 300252
rect 239260 300052 239324 300116
rect 227300 298692 227364 298756
rect 231532 297740 231596 297804
rect 224724 297604 224788 297668
rect 247908 297468 247972 297532
rect 306604 297468 306668 297532
rect 231716 297332 231780 297396
rect 291332 297332 291396 297396
rect 238892 296788 238956 296852
rect 238708 296516 238772 296580
rect 226564 296108 226628 296172
rect 228404 295972 228468 296036
rect 275324 294748 275388 294812
rect 229876 294612 229940 294676
rect 252876 294476 252940 294540
rect 277900 293252 277964 293316
rect 278084 293116 278148 293180
rect 275140 292028 275204 292092
rect 231164 291892 231228 291956
rect 242388 291756 242452 291820
rect 263548 291484 263612 291548
rect 260604 290804 260668 290868
rect 226932 290668 226996 290732
rect 245332 290532 245396 290596
rect 305684 290532 305748 290596
rect 257108 290396 257172 290460
rect 238892 290260 238956 290324
rect 249012 289988 249076 290052
rect 250484 289988 250548 290052
rect 255452 289988 255516 290052
rect 223620 289716 223684 289780
rect 269620 289852 269684 289916
rect 231900 289716 231964 289780
rect 235212 289716 235276 289780
rect 250668 289716 250732 289780
rect 255636 289716 255700 289780
rect 223988 289580 224052 289644
rect 235396 289580 235460 289644
rect 250300 289444 250364 289508
rect 251772 289580 251836 289644
rect 255820 289580 255884 289644
rect 282684 289036 282748 289100
rect 256188 287676 256252 287740
rect 263548 286996 263612 287060
rect 318012 286452 318076 286516
rect 284892 283460 284956 283524
rect 266492 271084 266556 271148
rect 267412 258844 267476 258908
rect 263732 258708 263796 258772
rect 310100 253948 310164 254012
rect 264100 247692 264164 247756
rect 266124 244972 266188 245036
rect 263548 244836 263612 244900
rect 267596 244216 267660 244220
rect 267596 244160 267610 244216
rect 267610 244160 267660 244216
rect 267596 244156 267660 244160
rect 264468 243884 264532 243948
rect 327580 243476 327644 243540
rect 264284 242252 264348 242316
rect 263732 242116 263796 242180
rect 322060 242116 322124 242180
rect 260972 241980 261036 242044
rect 264652 241844 264716 241908
rect 239076 241708 239140 241772
rect 258764 241572 258828 241636
rect 246620 241436 246684 241500
rect 302740 241436 302804 241500
rect 223252 241300 223316 241364
rect 226196 241300 226260 241364
rect 227668 241164 227732 241228
rect 223804 241028 223868 241092
rect 226012 241028 226076 241092
rect 234292 241028 234356 241092
rect 232452 240892 232516 240956
rect 265940 240892 266004 240956
rect 226932 240756 226996 240820
rect 228588 240756 228652 240820
rect 231164 240756 231228 240820
rect 229692 240620 229756 240684
rect 248276 240620 248340 240684
rect 295932 240620 295996 240684
rect 227484 240484 227548 240548
rect 223804 240348 223868 240412
rect 226012 240212 226076 240276
rect 223436 240076 223500 240140
rect 222516 239804 222580 239868
rect 224172 239842 224176 239868
rect 224176 239842 224232 239868
rect 224232 239842 224236 239868
rect 224172 239804 224236 239842
rect 224540 239804 224604 239868
rect 226012 239864 226076 239868
rect 226012 239808 226016 239864
rect 226016 239808 226072 239864
rect 226072 239808 226076 239864
rect 226012 239804 226076 239808
rect 230060 240348 230124 240412
rect 230428 240348 230492 240412
rect 230796 240348 230860 240412
rect 238340 240348 238404 240412
rect 226380 239940 226444 240004
rect 228220 240076 228284 240140
rect 227852 239940 227916 240004
rect 226564 239804 226628 239868
rect 227300 239842 227304 239868
rect 227304 239842 227360 239868
rect 227360 239842 227364 239868
rect 227300 239804 227364 239842
rect 230980 240212 231044 240276
rect 231900 240076 231964 240140
rect 231532 239940 231596 240004
rect 228220 239804 228284 239868
rect 230612 239804 230676 239868
rect 232268 239804 232332 239868
rect 237236 240076 237300 240140
rect 237420 239940 237484 240004
rect 238156 239940 238220 240004
rect 222700 239728 222764 239732
rect 222700 239672 222750 239728
rect 222750 239672 222764 239728
rect 222700 239668 222764 239672
rect 223068 239728 223132 239732
rect 223068 239672 223118 239728
rect 223118 239672 223132 239728
rect 223068 239668 223132 239672
rect 223252 239668 223316 239732
rect 223804 239728 223868 239732
rect 223804 239672 223854 239728
rect 223854 239672 223868 239728
rect 223804 239668 223868 239672
rect 224724 239668 224788 239732
rect 224908 239668 224972 239732
rect 226748 239728 226812 239732
rect 226748 239672 226762 239728
rect 226762 239672 226812 239728
rect 226748 239668 226812 239672
rect 226932 239728 226996 239732
rect 226932 239672 226946 239728
rect 226946 239672 226996 239728
rect 226932 239668 226996 239672
rect 228036 239668 228100 239732
rect 229876 239668 229940 239732
rect 230428 239728 230492 239732
rect 230428 239672 230442 239728
rect 230442 239672 230492 239728
rect 230428 239668 230492 239672
rect 230980 239668 231044 239732
rect 232084 239668 232148 239732
rect 232452 239668 232516 239732
rect 220676 239396 220740 239460
rect 223988 239592 224052 239596
rect 223988 239536 224002 239592
rect 224002 239536 224052 239592
rect 223988 239532 224052 239536
rect 226196 239532 226260 239596
rect 227116 239532 227180 239596
rect 227484 239532 227548 239596
rect 230796 239532 230860 239596
rect 231716 239532 231780 239596
rect 231900 239532 231964 239596
rect 233924 239842 233928 239868
rect 233928 239842 233984 239868
rect 233984 239842 233988 239868
rect 233924 239804 233988 239842
rect 234292 239864 234356 239868
rect 234292 239808 234296 239864
rect 234296 239808 234352 239864
rect 234352 239808 234356 239864
rect 234292 239804 234356 239808
rect 234660 239864 234724 239868
rect 234660 239808 234664 239864
rect 234664 239808 234720 239864
rect 234720 239808 234724 239864
rect 234660 239804 234724 239808
rect 235212 239804 235276 239868
rect 236132 239804 236196 239868
rect 243124 239940 243188 240004
rect 238524 239804 238588 239868
rect 239076 239804 239140 239868
rect 240916 239804 240980 239868
rect 242020 239804 242084 239868
rect 242756 239864 242820 239868
rect 242756 239808 242760 239864
rect 242760 239808 242816 239864
rect 242816 239808 242820 239864
rect 242756 239804 242820 239808
rect 246252 239864 246316 239868
rect 246252 239808 246266 239864
rect 246266 239808 246316 239864
rect 246252 239804 246316 239808
rect 246804 239804 246868 239868
rect 247540 239804 247604 239868
rect 248092 239804 248156 239868
rect 249012 239804 249076 239868
rect 250300 239804 250364 239868
rect 251036 239804 251100 239868
rect 251588 239804 251652 239868
rect 252876 239804 252940 239868
rect 233740 239668 233804 239732
rect 235396 239668 235460 239732
rect 233556 239532 233620 239596
rect 234476 239532 234540 239596
rect 238892 239668 238956 239732
rect 242388 239668 242452 239732
rect 244964 239668 245028 239732
rect 246068 239668 246132 239732
rect 247908 239728 247972 239732
rect 247908 239672 247922 239728
rect 247922 239672 247972 239728
rect 247908 239668 247972 239672
rect 248276 239668 248340 239732
rect 249564 239668 249628 239732
rect 250668 239668 250732 239732
rect 251956 239668 252020 239732
rect 252140 239668 252204 239732
rect 238708 239532 238772 239596
rect 239444 239532 239508 239596
rect 241284 239592 241348 239596
rect 241284 239536 241334 239592
rect 241334 239536 241348 239592
rect 241284 239532 241348 239536
rect 242204 239532 242268 239596
rect 243308 239532 243372 239596
rect 245516 239532 245580 239596
rect 246620 239532 246684 239596
rect 247724 239532 247788 239596
rect 253244 239668 253308 239732
rect 249380 239532 249444 239596
rect 251772 239532 251836 239596
rect 253060 239532 253124 239596
rect 227668 239396 227732 239460
rect 228588 239396 228652 239460
rect 236132 239396 236196 239460
rect 243492 239396 243556 239460
rect 247356 239396 247420 239460
rect 249196 239396 249260 239460
rect 250852 239396 250916 239460
rect 255636 239804 255700 239868
rect 256188 239804 256252 239868
rect 256924 239804 256988 239868
rect 259316 239940 259380 240004
rect 263916 239940 263980 240004
rect 256740 239668 256804 239732
rect 258948 239804 259012 239868
rect 260788 239804 260852 239868
rect 262076 239842 262080 239868
rect 262080 239842 262136 239868
rect 262136 239842 262140 239868
rect 262076 239804 262140 239842
rect 254716 239532 254780 239596
rect 255452 239532 255516 239596
rect 255820 239532 255884 239596
rect 256372 239592 256436 239596
rect 256372 239536 256386 239592
rect 256386 239536 256436 239592
rect 256372 239532 256436 239536
rect 257108 239532 257172 239596
rect 256740 239396 256804 239460
rect 258764 239532 258828 239596
rect 260604 239532 260668 239596
rect 260972 239592 261036 239596
rect 260972 239536 260986 239592
rect 260986 239536 261036 239592
rect 260972 239532 261036 239536
rect 238340 239260 238404 239324
rect 259132 239456 259196 239460
rect 262628 239668 262692 239732
rect 264284 239804 264348 239868
rect 263548 239728 263612 239732
rect 263548 239672 263562 239728
rect 263562 239672 263612 239728
rect 263548 239668 263612 239672
rect 264468 239668 264532 239732
rect 266492 239940 266556 240004
rect 267596 240000 267660 240004
rect 267596 239944 267610 240000
rect 267610 239944 267660 240000
rect 267596 239940 267660 239944
rect 265940 239864 266004 239868
rect 265940 239808 265944 239864
rect 265944 239808 266000 239864
rect 266000 239808 266004 239864
rect 265940 239804 266004 239808
rect 267412 239804 267476 239868
rect 265940 239668 266004 239732
rect 266124 239728 266188 239732
rect 266124 239672 266138 239728
rect 266138 239672 266188 239728
rect 266124 239668 266188 239672
rect 262628 239532 262692 239596
rect 259132 239400 259182 239456
rect 259182 239400 259196 239456
rect 259132 239396 259196 239400
rect 260236 239260 260300 239324
rect 262076 239260 262140 239324
rect 263548 239260 263612 239324
rect 229692 239184 229756 239188
rect 229692 239128 229742 239184
rect 229742 239128 229756 239184
rect 229692 239124 229756 239128
rect 241652 239124 241716 239188
rect 253428 239184 253492 239188
rect 253428 239128 253478 239184
rect 253478 239128 253492 239184
rect 253428 239124 253492 239128
rect 262076 239124 262140 239188
rect 264652 239124 264716 239188
rect 265940 239124 266004 239188
rect 227852 238716 227916 238780
rect 230244 238716 230308 238780
rect 231900 238580 231964 238644
rect 233924 238580 233988 238644
rect 234660 238640 234724 238644
rect 234660 238584 234674 238640
rect 234674 238584 234724 238640
rect 234660 238580 234724 238584
rect 242756 238580 242820 238644
rect 243308 238580 243372 238644
rect 245148 238580 245212 238644
rect 245332 238580 245396 238644
rect 246804 238580 246868 238644
rect 248276 238580 248340 238644
rect 249380 238580 249444 238644
rect 250116 238580 250180 238644
rect 253060 238640 253124 238644
rect 253060 238584 253110 238640
rect 253110 238584 253124 238640
rect 253060 238580 253124 238584
rect 226012 238444 226076 238508
rect 226564 238504 226628 238508
rect 226564 238448 226578 238504
rect 226578 238448 226628 238504
rect 226564 238444 226628 238448
rect 231532 238444 231596 238508
rect 232452 238444 232516 238508
rect 264284 238444 264348 238508
rect 267596 238368 267660 238372
rect 267596 238312 267610 238368
rect 267610 238312 267660 238368
rect 267596 238308 267660 238312
rect 226380 238172 226444 238236
rect 228588 238172 228652 238236
rect 230612 238172 230676 238236
rect 264100 238172 264164 238236
rect 224540 238036 224604 238100
rect 226748 238036 226812 238100
rect 228588 238036 228652 238100
rect 231716 238096 231780 238100
rect 231716 238040 231730 238096
rect 231730 238040 231780 238096
rect 231716 238036 231780 238040
rect 237236 238036 237300 238100
rect 227668 237900 227732 237964
rect 231348 237900 231412 237964
rect 240916 237900 240980 237964
rect 250484 237960 250548 237964
rect 250484 237904 250534 237960
rect 250534 237904 250548 237960
rect 250484 237900 250548 237904
rect 254716 237900 254780 237964
rect 256188 237900 256252 237964
rect 264468 237900 264532 237964
rect 222700 237492 222764 237556
rect 231532 237492 231596 237556
rect 229876 237356 229940 237420
rect 256740 237628 256804 237692
rect 260420 237552 260484 237556
rect 260420 237496 260434 237552
rect 260434 237496 260484 237552
rect 260420 237492 260484 237496
rect 235212 236812 235276 236876
rect 242388 236736 242452 236740
rect 242388 236680 242402 236736
rect 242402 236680 242452 236736
rect 242388 236676 242452 236680
rect 257108 236676 257172 236740
rect 260788 236676 260852 236740
rect 222516 236268 222580 236332
rect 224172 236268 224236 236332
rect 224908 236192 224972 236196
rect 224908 236136 224958 236192
rect 224958 236136 224972 236192
rect 224908 236132 224972 236136
rect 249564 236192 249628 236196
rect 249564 236136 249614 236192
rect 249614 236136 249628 236192
rect 249564 236132 249628 236136
rect 250668 236132 250732 236196
rect 228404 235996 228468 236060
rect 255084 235996 255148 236060
rect 241652 235920 241716 235924
rect 241652 235864 241666 235920
rect 241666 235864 241716 235920
rect 241652 235860 241716 235864
rect 254900 235860 254964 235924
rect 223436 235588 223500 235652
rect 234292 235316 234356 235380
rect 232268 235180 232332 235244
rect 256740 235180 256804 235244
rect 260052 235180 260116 235244
rect 263180 235180 263244 235244
rect 235764 234772 235828 234836
rect 235580 234500 235644 234564
rect 243124 234500 243188 234564
rect 230244 233956 230308 234020
rect 304396 233140 304460 233204
rect 256556 232868 256620 232932
rect 242756 232596 242820 232660
rect 299980 232596 300044 232660
rect 299796 231236 299860 231300
rect 246620 231100 246684 231164
rect 266124 230964 266188 231028
rect 242388 229740 242452 229804
rect 306052 229256 306116 229260
rect 306052 229200 306102 229256
rect 306102 229200 306116 229256
rect 306052 229196 306116 229200
rect 260420 228924 260484 228988
rect 253060 228652 253124 228716
rect 243492 228244 243556 228308
rect 302004 227624 302068 227628
rect 302004 227568 302054 227624
rect 302054 227568 302068 227624
rect 302004 227564 302068 227568
rect 242572 227292 242636 227356
rect 302188 227292 302252 227356
rect 311020 227156 311084 227220
rect 233740 227020 233804 227084
rect 239076 226884 239140 226948
rect 250116 226204 250180 226268
rect 306236 226204 306300 226268
rect 255084 225932 255148 225996
rect 263180 225796 263244 225860
rect 229876 224844 229940 224908
rect 294644 224844 294708 224908
rect 237420 224436 237484 224500
rect 235580 224300 235644 224364
rect 260236 224572 260300 224636
rect 262812 224436 262876 224500
rect 319300 224436 319364 224500
rect 262076 224300 262140 224364
rect 247724 224164 247788 224228
rect 256740 224028 256804 224092
rect 254900 223756 254964 223820
rect 227668 223484 227732 223548
rect 287836 223484 287900 223548
rect 246804 223348 246868 223412
rect 306420 223348 306484 223412
rect 248276 223212 248340 223276
rect 245148 223076 245212 223140
rect 303844 223076 303908 223140
rect 250852 222940 250916 223004
rect 313780 222940 313844 223004
rect 249380 222804 249444 222868
rect 234292 222668 234356 222732
rect 245332 222532 245396 222596
rect 305500 222532 305564 222596
rect 301820 222124 301884 222188
rect 294460 221988 294524 222052
rect 232452 221852 232516 221916
rect 292620 221852 292684 221916
rect 298140 221716 298204 221780
rect 251956 221580 252020 221644
rect 232452 221444 232516 221508
rect 256188 221444 256252 221508
rect 256924 221308 256988 221372
rect 264468 221172 264532 221236
rect 242756 220764 242820 220828
rect 285628 220628 285692 220692
rect 282868 220492 282932 220556
rect 228588 220356 228652 220420
rect 231348 220220 231412 220284
rect 231532 220084 231596 220148
rect 283420 220220 283484 220284
rect 287100 220220 287164 220284
rect 291148 219812 291212 219876
rect 284340 219268 284404 219332
rect 288388 219132 288452 219196
rect 303476 219192 303540 219196
rect 303476 219136 303490 219192
rect 303490 219136 303540 219192
rect 303476 219132 303540 219136
rect 260052 218996 260116 219060
rect 317460 218996 317524 219060
rect 235764 218860 235828 218924
rect 231716 218724 231780 218788
rect 257108 218588 257172 218652
rect 258948 218452 259012 218516
rect 230980 218044 231044 218108
rect 231716 218044 231780 218108
rect 235764 218044 235828 218108
rect 260052 218044 260116 218108
rect 243308 214508 243372 214572
rect 303660 213828 303724 213892
rect 228588 213148 228652 213212
rect 246252 213148 246316 213212
rect 244964 211788 245028 211852
rect 304212 208252 304276 208316
rect 233924 207572 233988 207636
rect 242388 204852 242452 204916
rect 231164 203492 231228 203556
rect 250852 202132 250916 202196
rect 227300 200636 227364 200700
rect 242572 200636 242636 200700
rect 238892 199412 238956 199476
rect 230060 199276 230124 199340
rect 247540 199276 247604 199340
rect 249380 197916 249444 197980
rect 226932 196556 226996 196620
rect 233740 193836 233804 193900
rect 246068 192476 246132 192540
rect 262996 190980 263060 191044
rect 263180 189620 263244 189684
rect 233556 188260 233620 188324
rect 245332 188260 245396 188324
rect 247356 186900 247420 186964
rect 230980 182820 231044 182884
rect 263732 182820 263796 182884
rect 249012 178604 249076 178668
rect 256740 168948 256804 169012
rect 249196 167588 249260 167652
rect 245516 166228 245580 166292
rect 239444 156572 239508 156636
rect 255084 156572 255148 156636
rect 246804 152356 246868 152420
rect 256924 150996 256988 151060
rect 258948 146916 259012 146980
rect 242204 141340 242268 141404
rect 251036 138620 251100 138684
rect 269620 125564 269684 125628
rect 281396 31724 281460 31788
rect 259132 25468 259196 25532
rect 257108 15812 257172 15876
rect 262628 10236 262692 10300
rect 252692 6836 252756 6900
rect 253244 6700 253308 6764
rect 256188 6564 256252 6628
rect 256372 6428 256436 6492
rect 256004 6292 256068 6356
rect 259316 6156 259380 6220
rect 248276 6020 248340 6084
rect 251588 3572 251652 3636
rect 252140 3436 252204 3500
rect 260604 3300 260668 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52674 522334 53294 557778
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 414334 53294 449778
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 56394 526054 57014 561498
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 56394 490054 57014 525498
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 130054 57014 165498
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 56394 94054 57014 129498
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 56394 58054 57014 93498
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 60114 565774 60734 601218
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 60114 529774 60734 565218
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 60114 493774 60734 529218
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 60114 421774 60734 457218
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 169774 60734 205218
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 97774 60734 133218
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 60114 61774 60734 97218
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 605494 64454 640938
rect 63834 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 64454 605494
rect 63834 605174 64454 605258
rect 63834 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 64454 605174
rect 63834 569494 64454 604938
rect 63834 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 64454 569494
rect 63834 569174 64454 569258
rect 63834 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 64454 569174
rect 63834 533494 64454 568938
rect 63834 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 64454 533494
rect 63834 533174 64454 533258
rect 63834 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 64454 533174
rect 63834 497494 64454 532938
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 63834 461494 64454 496938
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 63834 425494 64454 460938
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 63834 389494 64454 424938
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 281494 64454 316938
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 63834 245494 64454 280938
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 63834 209494 64454 244938
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 63834 173494 64454 208938
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 63834 137494 64454 172938
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 63834 101494 64454 136938
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63834 65494 64454 100938
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 630334 89294 665778
rect 88674 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 89294 630334
rect 88674 630014 89294 630098
rect 88674 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 89294 630014
rect 88674 594334 89294 629778
rect 88674 594098 88706 594334
rect 88942 594098 89026 594334
rect 89262 594098 89294 594334
rect 88674 594014 89294 594098
rect 88674 593778 88706 594014
rect 88942 593778 89026 594014
rect 89262 593778 89294 594014
rect 88674 558334 89294 593778
rect 88674 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 89294 558334
rect 88674 558014 89294 558098
rect 88674 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 89294 558014
rect 88674 522334 89294 557778
rect 88674 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 89294 522334
rect 88674 522014 89294 522098
rect 88674 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 89294 522014
rect 88674 486334 89294 521778
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 88674 450334 89294 485778
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 414334 89294 449778
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 306334 89294 341778
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 88674 270334 89294 305778
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 88674 234334 89294 269778
rect 88674 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 89294 234334
rect 88674 234014 89294 234098
rect 88674 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 89294 234014
rect 88674 198334 89294 233778
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 88674 162334 89294 197778
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 88674 126334 89294 161778
rect 88674 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 89294 126334
rect 88674 126014 89294 126098
rect 88674 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 89294 126014
rect 88674 90334 89294 125778
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 88674 54334 89294 89778
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 598054 93014 633498
rect 92394 597818 92426 598054
rect 92662 597818 92746 598054
rect 92982 597818 93014 598054
rect 92394 597734 93014 597818
rect 92394 597498 92426 597734
rect 92662 597498 92746 597734
rect 92982 597498 93014 597734
rect 92394 562054 93014 597498
rect 92394 561818 92426 562054
rect 92662 561818 92746 562054
rect 92982 561818 93014 562054
rect 92394 561734 93014 561818
rect 92394 561498 92426 561734
rect 92662 561498 92746 561734
rect 92982 561498 93014 561734
rect 92394 526054 93014 561498
rect 92394 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 93014 526054
rect 92394 525734 93014 525818
rect 92394 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 93014 525734
rect 92394 490054 93014 525498
rect 92394 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 93014 490054
rect 92394 489734 93014 489818
rect 92394 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 93014 489734
rect 92394 454054 93014 489498
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 418054 93014 453498
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 310054 93014 345498
rect 92394 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 93014 310054
rect 92394 309734 93014 309818
rect 92394 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 93014 309734
rect 92394 274054 93014 309498
rect 92394 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 93014 274054
rect 92394 273734 93014 273818
rect 92394 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 93014 273734
rect 92394 238054 93014 273498
rect 92394 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 93014 238054
rect 92394 237734 93014 237818
rect 92394 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 93014 237734
rect 92394 202054 93014 237498
rect 92394 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 93014 202054
rect 92394 201734 93014 201818
rect 92394 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 93014 201734
rect 92394 166054 93014 201498
rect 92394 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 93014 166054
rect 92394 165734 93014 165818
rect 92394 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 93014 165734
rect 92394 130054 93014 165498
rect 92394 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 93014 130054
rect 92394 129734 93014 129818
rect 92394 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 93014 129734
rect 92394 94054 93014 129498
rect 92394 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 93014 94054
rect 92394 93734 93014 93818
rect 92394 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 93014 93734
rect 92394 58054 93014 93498
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 96114 601774 96734 637218
rect 96114 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 96734 601774
rect 96114 601454 96734 601538
rect 96114 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 96734 601454
rect 96114 565774 96734 601218
rect 96114 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 96734 565774
rect 96114 565454 96734 565538
rect 96114 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 96734 565454
rect 96114 529774 96734 565218
rect 96114 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 96734 529774
rect 96114 529454 96734 529538
rect 96114 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 96734 529454
rect 96114 493774 96734 529218
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 96114 457774 96734 493218
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 96114 421774 96734 457218
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 313774 96734 349218
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 96114 277774 96734 313218
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 96114 241774 96734 277218
rect 96114 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 96734 241774
rect 96114 241454 96734 241538
rect 96114 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 96734 241454
rect 96114 205774 96734 241218
rect 96114 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 96734 205774
rect 96114 205454 96734 205538
rect 96114 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 96734 205454
rect 96114 169774 96734 205218
rect 96114 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 96734 169774
rect 96114 169454 96734 169538
rect 96114 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 96734 169454
rect 96114 133774 96734 169218
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 96114 97774 96734 133218
rect 96114 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 96734 97774
rect 96114 97454 96734 97538
rect 96114 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 96734 97454
rect 96114 61774 96734 97218
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 96114 25774 96734 61218
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 605494 100454 640938
rect 99834 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 100454 605494
rect 99834 605174 100454 605258
rect 99834 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 100454 605174
rect 99834 569494 100454 604938
rect 99834 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 100454 569494
rect 99834 569174 100454 569258
rect 99834 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 100454 569174
rect 99834 533494 100454 568938
rect 99834 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 100454 533494
rect 99834 533174 100454 533258
rect 99834 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 100454 533174
rect 99834 497494 100454 532938
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 99834 461494 100454 496938
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 425494 100454 460938
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 317494 100454 352938
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 99834 281494 100454 316938
rect 99834 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 100454 281494
rect 99834 281174 100454 281258
rect 99834 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 100454 281174
rect 99834 245494 100454 280938
rect 99834 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 100454 245494
rect 99834 245174 100454 245258
rect 99834 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 100454 245174
rect 99834 209494 100454 244938
rect 99834 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 100454 209494
rect 99834 209174 100454 209258
rect 99834 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 100454 209174
rect 99834 173494 100454 208938
rect 99834 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 100454 173494
rect 99834 173174 100454 173258
rect 99834 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 100454 173174
rect 99834 137494 100454 172938
rect 99834 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 100454 137494
rect 99834 137174 100454 137258
rect 99834 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 100454 137174
rect 99834 101494 100454 136938
rect 99834 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 100454 101494
rect 99834 101174 100454 101258
rect 99834 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 100454 101174
rect 99834 65494 100454 100938
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 99834 29494 100454 64938
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 630334 125294 665778
rect 124674 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 125294 630334
rect 124674 630014 125294 630098
rect 124674 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 125294 630014
rect 124674 594334 125294 629778
rect 124674 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 125294 594334
rect 124674 594014 125294 594098
rect 124674 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 125294 594014
rect 124674 558334 125294 593778
rect 124674 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 125294 558334
rect 124674 558014 125294 558098
rect 124674 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 125294 558014
rect 124674 522334 125294 557778
rect 124674 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 125294 522334
rect 124674 522014 125294 522098
rect 124674 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 125294 522014
rect 124674 486334 125294 521778
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124674 126334 125294 161778
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 124674 90334 125294 125778
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 124674 54334 125294 89778
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 598054 129014 633498
rect 128394 597818 128426 598054
rect 128662 597818 128746 598054
rect 128982 597818 129014 598054
rect 128394 597734 129014 597818
rect 128394 597498 128426 597734
rect 128662 597498 128746 597734
rect 128982 597498 129014 597734
rect 128394 562054 129014 597498
rect 128394 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 129014 562054
rect 128394 561734 129014 561818
rect 128394 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 129014 561734
rect 128394 526054 129014 561498
rect 128394 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 129014 526054
rect 128394 525734 129014 525818
rect 128394 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 129014 525734
rect 128394 490054 129014 525498
rect 128394 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 129014 490054
rect 128394 489734 129014 489818
rect 128394 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 129014 489734
rect 128394 454054 129014 489498
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 128394 418054 129014 453498
rect 128394 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 129014 418054
rect 128394 417734 129014 417818
rect 128394 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 129014 417734
rect 128394 382054 129014 417498
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 128394 130054 129014 165498
rect 128394 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 129014 130054
rect 128394 129734 129014 129818
rect 128394 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 129014 129734
rect 128394 94054 129014 129498
rect 128394 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 129014 94054
rect 128394 93734 129014 93818
rect 128394 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 129014 93734
rect 128394 58054 129014 93498
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 601774 132734 637218
rect 132114 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 132734 601774
rect 132114 601454 132734 601538
rect 132114 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 132734 601454
rect 132114 565774 132734 601218
rect 132114 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 132734 565774
rect 132114 565454 132734 565538
rect 132114 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 132734 565454
rect 132114 529774 132734 565218
rect 132114 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 132734 529774
rect 132114 529454 132734 529538
rect 132114 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 132734 529454
rect 132114 493774 132734 529218
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 132114 457774 132734 493218
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 421774 132734 457218
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 132114 385774 132734 421218
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 97774 132734 133218
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 132114 61774 132734 97218
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 132114 25774 132734 61218
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 135834 605494 136454 640938
rect 135834 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 136454 605494
rect 135834 605174 136454 605258
rect 135834 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 136454 605174
rect 135834 569494 136454 604938
rect 135834 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 136454 569494
rect 135834 569174 136454 569258
rect 135834 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 136454 569174
rect 135834 533494 136454 568938
rect 135834 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 136454 533494
rect 135834 533174 136454 533258
rect 135834 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 136454 533174
rect 135834 497494 136454 532938
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 135834 461494 136454 496938
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 425494 136454 460938
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 135834 389494 136454 424938
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 135834 353494 136454 388938
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 173494 136454 208938
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 135834 137494 136454 172938
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 135834 101494 136454 136938
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 594334 161294 629778
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 160674 558334 161294 593778
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 160674 522334 161294 557778
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 160674 486334 161294 521778
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 160674 450334 161294 485778
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 160674 414334 161294 449778
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 160674 378334 161294 413778
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 598054 165014 633498
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 164394 562054 165014 597498
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 164394 526054 165014 561498
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 164394 490054 165014 525498
rect 164394 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 165014 490054
rect 164394 489734 165014 489818
rect 164394 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 165014 489734
rect 164394 454054 165014 489498
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 418054 165014 453498
rect 164394 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 165014 418054
rect 164394 417734 165014 417818
rect 164394 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 165014 417734
rect 164394 382054 165014 417498
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 168114 529774 168734 565218
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 493774 168734 529218
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 168114 457774 168734 493218
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 421774 168734 457218
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 168114 385774 168734 421218
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171834 569494 172454 604938
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171834 533494 172454 568938
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171834 497494 172454 532938
rect 171834 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 172454 497494
rect 171834 497174 172454 497258
rect 171834 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 172454 497174
rect 171834 461494 172454 496938
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 171834 425494 172454 460938
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 171834 389494 172454 424938
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 171834 353494 172454 388938
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 594334 197294 629778
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 196674 558334 197294 593778
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 486334 197294 521778
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 196674 450334 197294 485778
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 196674 414334 197294 449778
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 196674 378334 197294 413778
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 196674 234334 197294 269778
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 196674 162334 197294 197778
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 598054 201014 633498
rect 200394 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 201014 598054
rect 200394 597734 201014 597818
rect 200394 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 201014 597734
rect 200394 562054 201014 597498
rect 200394 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 201014 562054
rect 200394 561734 201014 561818
rect 200394 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 201014 561734
rect 200394 526054 201014 561498
rect 200394 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 201014 526054
rect 200394 525734 201014 525818
rect 200394 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 201014 525734
rect 200394 490054 201014 525498
rect 200394 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 201014 490054
rect 200394 489734 201014 489818
rect 200394 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 201014 489734
rect 200394 454054 201014 489498
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 418054 201014 453498
rect 200394 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 201014 418054
rect 200394 417734 201014 417818
rect 200394 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 201014 417734
rect 200394 382054 201014 417498
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 200394 238054 201014 273498
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 601774 204734 637218
rect 204114 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 204734 601774
rect 204114 601454 204734 601538
rect 204114 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 204734 601454
rect 204114 565774 204734 601218
rect 204114 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 204734 565774
rect 204114 565454 204734 565538
rect 204114 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 204734 565454
rect 204114 529774 204734 565218
rect 204114 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 204734 529774
rect 204114 529454 204734 529538
rect 204114 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 204734 529454
rect 204114 493774 204734 529218
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 204114 457774 204734 493218
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 204114 421774 204734 457218
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 204114 385774 204734 421218
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 207834 569494 208454 604938
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 207834 533494 208454 568938
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 207834 497494 208454 532938
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 207834 461494 208454 496938
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 425494 208454 460938
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 207834 389494 208454 424938
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 207834 353494 208454 388938
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 207834 173494 208454 208938
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 220675 318612 220741 318613
rect 220675 318548 220676 318612
rect 220740 318548 220741 318612
rect 220675 318547 220741 318548
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 220678 239461 220738 318547
rect 221514 295174 222134 330618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 223435 315484 223501 315485
rect 223435 315420 223436 315484
rect 223500 315420 223501 315484
rect 223435 315419 223501 315420
rect 222699 314668 222765 314669
rect 222699 314604 222700 314668
rect 222764 314604 222765 314668
rect 222699 314603 222765 314604
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 220675 239460 220741 239461
rect 220675 239396 220676 239460
rect 220740 239396 220741 239460
rect 220675 239395 220741 239396
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 223174 222134 258618
rect 222515 239868 222581 239869
rect 222515 239804 222516 239868
rect 222580 239804 222581 239868
rect 222515 239803 222581 239804
rect 222518 236333 222578 239803
rect 222702 239733 222762 314603
rect 223067 307460 223133 307461
rect 223067 307396 223068 307460
rect 223132 307396 223133 307460
rect 223067 307395 223133 307396
rect 223070 239733 223130 307395
rect 223251 241364 223317 241365
rect 223251 241300 223252 241364
rect 223316 241300 223317 241364
rect 223251 241299 223317 241300
rect 223254 239733 223314 241299
rect 223438 240141 223498 315419
rect 225234 298894 225854 334338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 226747 317116 226813 317117
rect 226747 317052 226748 317116
rect 226812 317052 226813 317116
rect 226747 317051 226813 317052
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 224723 297668 224789 297669
rect 224723 297604 224724 297668
rect 224788 297604 224789 297668
rect 224723 297603 224789 297604
rect 223619 289780 223685 289781
rect 223619 289716 223620 289780
rect 223684 289716 223685 289780
rect 223619 289715 223685 289716
rect 223435 240140 223501 240141
rect 223435 240076 223436 240140
rect 223500 240076 223501 240140
rect 223435 240075 223501 240076
rect 222699 239732 222765 239733
rect 222699 239668 222700 239732
rect 222764 239668 222765 239732
rect 222699 239667 222765 239668
rect 223067 239732 223133 239733
rect 223067 239668 223068 239732
rect 223132 239668 223133 239732
rect 223067 239667 223133 239668
rect 223251 239732 223317 239733
rect 223251 239668 223252 239732
rect 223316 239668 223317 239732
rect 223251 239667 223317 239668
rect 222702 237557 222762 239667
rect 222699 237556 222765 237557
rect 222699 237492 222700 237556
rect 222764 237492 222765 237556
rect 222699 237491 222765 237492
rect 222515 236332 222581 236333
rect 222515 236268 222516 236332
rect 222580 236268 222581 236332
rect 222515 236267 222581 236268
rect 223438 235653 223498 240075
rect 223622 239730 223682 289715
rect 223987 289644 224053 289645
rect 223987 289580 223988 289644
rect 224052 289580 224053 289644
rect 223987 289579 224053 289580
rect 223803 241092 223869 241093
rect 223803 241028 223804 241092
rect 223868 241028 223869 241092
rect 223803 241027 223869 241028
rect 223806 240413 223866 241027
rect 223803 240412 223869 240413
rect 223803 240348 223804 240412
rect 223868 240348 223869 240412
rect 223803 240347 223869 240348
rect 223803 239732 223869 239733
rect 223803 239730 223804 239732
rect 223622 239670 223804 239730
rect 223803 239668 223804 239670
rect 223868 239668 223869 239732
rect 223803 239667 223869 239668
rect 223990 239597 224050 289579
rect 224208 255454 224528 255486
rect 224208 255218 224250 255454
rect 224486 255218 224528 255454
rect 224208 255134 224528 255218
rect 224208 254898 224250 255134
rect 224486 254898 224528 255134
rect 224208 254866 224528 254898
rect 224171 239868 224237 239869
rect 224171 239804 224172 239868
rect 224236 239804 224237 239868
rect 224171 239803 224237 239804
rect 224539 239868 224605 239869
rect 224539 239804 224540 239868
rect 224604 239804 224605 239868
rect 224539 239803 224605 239804
rect 223987 239596 224053 239597
rect 223987 239532 223988 239596
rect 224052 239532 224053 239596
rect 223987 239531 224053 239532
rect 224174 236333 224234 239803
rect 224542 238101 224602 239803
rect 224726 239733 224786 297603
rect 225234 262894 225854 298338
rect 226563 296172 226629 296173
rect 226563 296108 226564 296172
rect 226628 296108 226629 296172
rect 226563 296107 226629 296108
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 224723 239732 224789 239733
rect 224723 239668 224724 239732
rect 224788 239668 224789 239732
rect 224723 239667 224789 239668
rect 224907 239732 224973 239733
rect 224907 239668 224908 239732
rect 224972 239668 224973 239732
rect 224907 239667 224973 239668
rect 224539 238100 224605 238101
rect 224539 238036 224540 238100
rect 224604 238036 224605 238100
rect 224539 238035 224605 238036
rect 224171 236332 224237 236333
rect 224171 236268 224172 236332
rect 224236 236268 224237 236332
rect 224171 236267 224237 236268
rect 224910 236197 224970 239667
rect 224907 236196 224973 236197
rect 224907 236132 224908 236196
rect 224972 236132 224973 236196
rect 224907 236131 224973 236132
rect 223435 235652 223501 235653
rect 223435 235588 223436 235652
rect 223500 235588 223501 235652
rect 223435 235587 223501 235588
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 226894 225854 262338
rect 226195 241364 226261 241365
rect 226195 241300 226196 241364
rect 226260 241300 226261 241364
rect 226195 241299 226261 241300
rect 226011 241092 226077 241093
rect 226011 241028 226012 241092
rect 226076 241028 226077 241092
rect 226011 241027 226077 241028
rect 226014 240277 226074 241027
rect 226011 240276 226077 240277
rect 226011 240212 226012 240276
rect 226076 240212 226077 240276
rect 226011 240211 226077 240212
rect 226011 239868 226077 239869
rect 226011 239804 226012 239868
rect 226076 239804 226077 239868
rect 226011 239803 226077 239804
rect 226014 238509 226074 239803
rect 226198 239597 226258 241299
rect 226379 240004 226445 240005
rect 226379 239940 226380 240004
rect 226444 239940 226445 240004
rect 226379 239939 226445 239940
rect 226195 239596 226261 239597
rect 226195 239532 226196 239596
rect 226260 239532 226261 239596
rect 226195 239531 226261 239532
rect 226011 238508 226077 238509
rect 226011 238444 226012 238508
rect 226076 238444 226077 238508
rect 226011 238443 226077 238444
rect 226382 238237 226442 239939
rect 226566 239869 226626 296107
rect 226563 239868 226629 239869
rect 226563 239804 226564 239868
rect 226628 239804 226629 239868
rect 226563 239803 226629 239804
rect 226566 238509 226626 239803
rect 226750 239733 226810 317051
rect 228219 304332 228285 304333
rect 228219 304268 228220 304332
rect 228284 304268 228285 304332
rect 228219 304267 228285 304268
rect 227851 304196 227917 304197
rect 227851 304132 227852 304196
rect 227916 304132 227917 304196
rect 227851 304131 227917 304132
rect 227299 298756 227365 298757
rect 227299 298692 227300 298756
rect 227364 298692 227365 298756
rect 227299 298691 227365 298692
rect 226931 290732 226997 290733
rect 226931 290668 226932 290732
rect 226996 290668 226997 290732
rect 226931 290667 226997 290668
rect 226934 245670 226994 290667
rect 226934 245610 227178 245670
rect 226931 240820 226997 240821
rect 226931 240756 226932 240820
rect 226996 240756 226997 240820
rect 226931 240755 226997 240756
rect 226934 239733 226994 240755
rect 226747 239732 226813 239733
rect 226747 239668 226748 239732
rect 226812 239668 226813 239732
rect 226747 239667 226813 239668
rect 226931 239732 226997 239733
rect 226931 239668 226932 239732
rect 226996 239668 226997 239732
rect 226931 239667 226997 239668
rect 226563 238508 226629 238509
rect 226563 238444 226564 238508
rect 226628 238444 226629 238508
rect 226563 238443 226629 238444
rect 226379 238236 226445 238237
rect 226379 238172 226380 238236
rect 226444 238172 226445 238236
rect 226379 238171 226445 238172
rect 226750 238101 226810 239667
rect 227118 239597 227178 245610
rect 227302 239869 227362 298691
rect 227667 241228 227733 241229
rect 227667 241164 227668 241228
rect 227732 241164 227733 241228
rect 227667 241163 227733 241164
rect 227483 240548 227549 240549
rect 227483 240484 227484 240548
rect 227548 240484 227549 240548
rect 227483 240483 227549 240484
rect 227299 239868 227365 239869
rect 227299 239804 227300 239868
rect 227364 239804 227365 239868
rect 227299 239803 227365 239804
rect 227115 239596 227181 239597
rect 227115 239532 227116 239596
rect 227180 239532 227181 239596
rect 227115 239531 227181 239532
rect 226747 238100 226813 238101
rect 226747 238036 226748 238100
rect 226812 238036 226813 238100
rect 226747 238035 226813 238036
rect 227118 234630 227178 239531
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 226934 234570 227178 234630
rect 226934 196621 226994 234570
rect 227302 200701 227362 239803
rect 227486 239597 227546 240483
rect 227483 239596 227549 239597
rect 227483 239532 227484 239596
rect 227548 239532 227549 239596
rect 227483 239531 227549 239532
rect 227670 239461 227730 241163
rect 227854 240005 227914 304131
rect 228035 302836 228101 302837
rect 228035 302772 228036 302836
rect 228100 302772 228101 302836
rect 228035 302771 228101 302772
rect 227851 240004 227917 240005
rect 227851 239940 227852 240004
rect 227916 239940 227917 240004
rect 227851 239939 227917 239940
rect 227667 239460 227733 239461
rect 227667 239396 227668 239460
rect 227732 239396 227733 239460
rect 227667 239395 227733 239396
rect 227854 238781 227914 239939
rect 228038 239733 228098 302771
rect 228222 240141 228282 304267
rect 228954 302614 229574 338058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 594334 233294 629778
rect 232674 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 233294 594334
rect 232674 594014 233294 594098
rect 232674 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 233294 594014
rect 232674 558334 233294 593778
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522334 233294 557778
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 232674 486334 233294 521778
rect 232674 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 233294 486334
rect 232674 486014 233294 486098
rect 232674 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 233294 486014
rect 232674 450334 233294 485778
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 232674 414334 233294 449778
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 232674 378334 233294 413778
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 232674 342334 233294 377778
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232267 318884 232333 318885
rect 232267 318820 232268 318884
rect 232332 318820 232333 318884
rect 232267 318819 232333 318820
rect 232083 315756 232149 315757
rect 232083 315692 232084 315756
rect 232148 315692 232149 315756
rect 232083 315691 232149 315692
rect 230979 308684 231045 308685
rect 230979 308620 230980 308684
rect 231044 308620 231045 308684
rect 230979 308619 231045 308620
rect 230243 307596 230309 307597
rect 230243 307532 230244 307596
rect 230308 307532 230309 307596
rect 230243 307531 230309 307532
rect 230059 307324 230125 307325
rect 230059 307260 230060 307324
rect 230124 307260 230125 307324
rect 230059 307259 230125 307260
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228403 296036 228469 296037
rect 228403 295972 228404 296036
rect 228468 295972 228469 296036
rect 228403 295971 228469 295972
rect 228219 240140 228285 240141
rect 228219 240076 228220 240140
rect 228284 240076 228285 240140
rect 228219 240075 228285 240076
rect 228219 239868 228285 239869
rect 228219 239804 228220 239868
rect 228284 239866 228285 239868
rect 228406 239866 228466 295971
rect 228954 266614 229574 302058
rect 229875 294676 229941 294677
rect 229875 294612 229876 294676
rect 229940 294612 229941 294676
rect 229875 294611 229941 294612
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228587 240820 228653 240821
rect 228587 240756 228588 240820
rect 228652 240756 228653 240820
rect 228587 240755 228653 240756
rect 228284 239806 228466 239866
rect 228284 239804 228285 239806
rect 228219 239803 228285 239804
rect 228035 239732 228101 239733
rect 228035 239668 228036 239732
rect 228100 239668 228101 239732
rect 228035 239667 228101 239668
rect 227851 238780 227917 238781
rect 227851 238716 227852 238780
rect 227916 238716 227917 238780
rect 227851 238715 227917 238716
rect 227667 237964 227733 237965
rect 227667 237900 227668 237964
rect 227732 237900 227733 237964
rect 227667 237899 227733 237900
rect 227670 223549 227730 237899
rect 228406 236061 228466 239806
rect 228590 239461 228650 240755
rect 228587 239460 228653 239461
rect 228587 239396 228588 239460
rect 228652 239396 228653 239460
rect 228587 239395 228653 239396
rect 228590 238237 228650 239395
rect 228587 238236 228653 238237
rect 228587 238172 228588 238236
rect 228652 238172 228653 238236
rect 228587 238171 228653 238172
rect 228587 238100 228653 238101
rect 228587 238036 228588 238100
rect 228652 238036 228653 238100
rect 228587 238035 228653 238036
rect 228403 236060 228469 236061
rect 228403 235996 228404 236060
rect 228468 235996 228469 236060
rect 228403 235995 228469 235996
rect 227667 223548 227733 223549
rect 227667 223484 227668 223548
rect 227732 223484 227733 223548
rect 227667 223483 227733 223484
rect 228590 220421 228650 238035
rect 228954 230614 229574 266058
rect 229691 240684 229757 240685
rect 229691 240620 229692 240684
rect 229756 240620 229757 240684
rect 229691 240619 229757 240620
rect 229694 239189 229754 240619
rect 229878 239733 229938 294611
rect 230062 240413 230122 307259
rect 230059 240412 230125 240413
rect 230059 240348 230060 240412
rect 230124 240348 230125 240412
rect 230059 240347 230125 240348
rect 229875 239732 229941 239733
rect 229875 239668 229876 239732
rect 229940 239668 229941 239732
rect 229875 239667 229941 239668
rect 229691 239188 229757 239189
rect 229691 239124 229692 239188
rect 229756 239124 229757 239188
rect 229691 239123 229757 239124
rect 229875 237420 229941 237421
rect 229875 237356 229876 237420
rect 229940 237356 229941 237420
rect 229875 237355 229941 237356
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228587 220420 228653 220421
rect 228587 220356 228588 220420
rect 228652 220356 228653 220420
rect 228587 220355 228653 220356
rect 228590 213213 228650 220355
rect 228587 213212 228653 213213
rect 228587 213148 228588 213212
rect 228652 213148 228653 213212
rect 228587 213147 228653 213148
rect 227299 200700 227365 200701
rect 227299 200636 227300 200700
rect 227364 200636 227365 200700
rect 227299 200635 227365 200636
rect 226931 196620 226997 196621
rect 226931 196556 226932 196620
rect 226996 196556 226997 196620
rect 226931 196555 226997 196556
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 194614 229574 230058
rect 229878 224909 229938 237355
rect 229875 224908 229941 224909
rect 229875 224844 229876 224908
rect 229940 224844 229941 224908
rect 229875 224843 229941 224844
rect 230062 199341 230122 240347
rect 230246 238781 230306 307531
rect 230427 240412 230493 240413
rect 230427 240348 230428 240412
rect 230492 240348 230493 240412
rect 230427 240347 230493 240348
rect 230795 240412 230861 240413
rect 230795 240348 230796 240412
rect 230860 240348 230861 240412
rect 230795 240347 230861 240348
rect 230430 239733 230490 240347
rect 230611 239868 230677 239869
rect 230611 239804 230612 239868
rect 230676 239804 230677 239868
rect 230611 239803 230677 239804
rect 230427 239732 230493 239733
rect 230427 239668 230428 239732
rect 230492 239668 230493 239732
rect 230427 239667 230493 239668
rect 230243 238780 230309 238781
rect 230243 238716 230244 238780
rect 230308 238716 230309 238780
rect 230243 238715 230309 238716
rect 230246 234021 230306 238715
rect 230614 238237 230674 239803
rect 230798 239597 230858 240347
rect 230982 240277 231042 308619
rect 231531 297804 231597 297805
rect 231531 297740 231532 297804
rect 231596 297740 231597 297804
rect 231531 297739 231597 297740
rect 231163 291956 231229 291957
rect 231163 291892 231164 291956
rect 231228 291892 231229 291956
rect 231163 291891 231229 291892
rect 231166 240821 231226 291891
rect 231534 245670 231594 297739
rect 231715 297396 231781 297397
rect 231715 297332 231716 297396
rect 231780 297332 231781 297396
rect 231715 297331 231781 297332
rect 231350 245610 231594 245670
rect 231163 240820 231229 240821
rect 231163 240756 231164 240820
rect 231228 240756 231229 240820
rect 231163 240755 231229 240756
rect 230979 240276 231045 240277
rect 230979 240212 230980 240276
rect 231044 240212 231045 240276
rect 230979 240211 231045 240212
rect 230979 239732 231045 239733
rect 230979 239668 230980 239732
rect 231044 239730 231045 239732
rect 231350 239730 231410 245610
rect 231531 240004 231597 240005
rect 231531 239940 231532 240004
rect 231596 239940 231597 240004
rect 231531 239939 231597 239940
rect 231044 239670 231410 239730
rect 231044 239668 231045 239670
rect 230979 239667 231045 239668
rect 230795 239596 230861 239597
rect 230795 239532 230796 239596
rect 230860 239532 230861 239596
rect 230795 239531 230861 239532
rect 231534 238509 231594 239939
rect 231718 239597 231778 297331
rect 231899 289780 231965 289781
rect 231899 289716 231900 289780
rect 231964 289716 231965 289780
rect 231899 289715 231965 289716
rect 231902 240141 231962 289715
rect 231899 240140 231965 240141
rect 231899 240076 231900 240140
rect 231964 240076 231965 240140
rect 231899 240075 231965 240076
rect 232086 239733 232146 315691
rect 232270 239869 232330 318819
rect 232674 306334 233294 341778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 598054 237014 633498
rect 236394 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 237014 598054
rect 236394 597734 237014 597818
rect 236394 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 237014 597734
rect 236394 562054 237014 597498
rect 236394 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 237014 562054
rect 236394 561734 237014 561818
rect 236394 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 237014 561734
rect 236394 526054 237014 561498
rect 236394 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 237014 526054
rect 236394 525734 237014 525818
rect 236394 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 237014 525734
rect 236394 490054 237014 525498
rect 236394 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 237014 490054
rect 236394 489734 237014 489818
rect 236394 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 237014 489734
rect 236394 454054 237014 489498
rect 236394 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 237014 454054
rect 236394 453734 237014 453818
rect 236394 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 237014 453734
rect 236394 418054 237014 453498
rect 236394 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 237014 418054
rect 236394 417734 237014 417818
rect 236394 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 237014 417734
rect 236394 382054 237014 417498
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236394 346054 237014 381498
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 234475 310996 234541 310997
rect 234475 310932 234476 310996
rect 234540 310932 234541 310996
rect 234475 310931 234541 310932
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 270334 233294 305778
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 232451 240956 232517 240957
rect 232451 240892 232452 240956
rect 232516 240892 232517 240956
rect 232451 240891 232517 240892
rect 232267 239868 232333 239869
rect 232267 239804 232268 239868
rect 232332 239804 232333 239868
rect 232267 239803 232333 239804
rect 232083 239732 232149 239733
rect 232083 239668 232084 239732
rect 232148 239668 232149 239732
rect 232083 239667 232149 239668
rect 231715 239596 231781 239597
rect 231715 239532 231716 239596
rect 231780 239532 231781 239596
rect 231715 239531 231781 239532
rect 231899 239596 231965 239597
rect 231899 239532 231900 239596
rect 231964 239532 231965 239596
rect 231899 239531 231965 239532
rect 231902 238645 231962 239531
rect 231899 238644 231965 238645
rect 231899 238580 231900 238644
rect 231964 238580 231965 238644
rect 231899 238579 231965 238580
rect 231531 238508 231597 238509
rect 231531 238444 231532 238508
rect 231596 238444 231597 238508
rect 231531 238443 231597 238444
rect 230611 238236 230677 238237
rect 230611 238172 230612 238236
rect 230676 238172 230677 238236
rect 230611 238171 230677 238172
rect 231715 238100 231781 238101
rect 231715 238036 231716 238100
rect 231780 238036 231781 238100
rect 231715 238035 231781 238036
rect 231347 237964 231413 237965
rect 231347 237900 231348 237964
rect 231412 237900 231413 237964
rect 231347 237899 231413 237900
rect 230243 234020 230309 234021
rect 230243 233956 230244 234020
rect 230308 233956 230309 234020
rect 230243 233955 230309 233956
rect 231350 220285 231410 237899
rect 231531 237556 231597 237557
rect 231531 237492 231532 237556
rect 231596 237492 231597 237556
rect 231531 237491 231597 237492
rect 231347 220284 231413 220285
rect 231347 220220 231348 220284
rect 231412 220220 231413 220284
rect 231347 220219 231413 220220
rect 231534 220149 231594 237491
rect 231531 220148 231597 220149
rect 231531 220084 231532 220148
rect 231596 220084 231597 220148
rect 231531 220083 231597 220084
rect 231534 219450 231594 220083
rect 231166 219390 231594 219450
rect 230979 218108 231045 218109
rect 230979 218044 230980 218108
rect 231044 218044 231045 218108
rect 230979 218043 231045 218044
rect 230059 199340 230125 199341
rect 230059 199276 230060 199340
rect 230124 199276 230125 199340
rect 230059 199275 230125 199276
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 230982 182885 231042 218043
rect 231166 203557 231226 219390
rect 231718 218789 231778 238035
rect 232270 235245 232330 239803
rect 232454 239733 232514 240891
rect 232451 239732 232517 239733
rect 232451 239668 232452 239732
rect 232516 239668 232517 239732
rect 232451 239667 232517 239668
rect 232451 238508 232517 238509
rect 232451 238444 232452 238508
rect 232516 238444 232517 238508
rect 232451 238443 232517 238444
rect 232267 235244 232333 235245
rect 232267 235180 232268 235244
rect 232332 235180 232333 235244
rect 232267 235179 232333 235180
rect 232454 221917 232514 238443
rect 232674 234334 233294 269778
rect 234291 241092 234357 241093
rect 234291 241028 234292 241092
rect 234356 241028 234357 241092
rect 234291 241027 234357 241028
rect 234294 239869 234354 241027
rect 233923 239868 233989 239869
rect 233923 239804 233924 239868
rect 233988 239804 233989 239868
rect 233923 239803 233989 239804
rect 234291 239868 234357 239869
rect 234291 239804 234292 239868
rect 234356 239804 234357 239868
rect 234291 239803 234357 239804
rect 233739 239732 233805 239733
rect 233739 239668 233740 239732
rect 233804 239668 233805 239732
rect 233739 239667 233805 239668
rect 233555 239596 233621 239597
rect 233555 239532 233556 239596
rect 233620 239532 233621 239596
rect 233555 239531 233621 239532
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232451 221916 232517 221917
rect 232451 221852 232452 221916
rect 232516 221852 232517 221916
rect 232451 221851 232517 221852
rect 232454 221509 232514 221851
rect 232451 221508 232517 221509
rect 232451 221444 232452 221508
rect 232516 221444 232517 221508
rect 232451 221443 232517 221444
rect 231715 218788 231781 218789
rect 231715 218724 231716 218788
rect 231780 218724 231781 218788
rect 231715 218723 231781 218724
rect 231718 218109 231778 218723
rect 231715 218108 231781 218109
rect 231715 218044 231716 218108
rect 231780 218044 231781 218108
rect 231715 218043 231781 218044
rect 231163 203556 231229 203557
rect 231163 203492 231164 203556
rect 231228 203492 231229 203556
rect 231163 203491 231229 203492
rect 232674 198334 233294 233778
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 230979 182884 231045 182885
rect 230979 182820 230980 182884
rect 231044 182820 231045 182884
rect 230979 182819 231045 182820
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 162334 233294 197778
rect 233558 188325 233618 239531
rect 233742 227085 233802 239667
rect 233926 238645 233986 239803
rect 234478 239597 234538 310931
rect 236394 310054 237014 345498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 601774 240734 637218
rect 240114 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 240734 601774
rect 240114 601454 240734 601538
rect 240114 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 240734 601454
rect 240114 565774 240734 601218
rect 240114 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 240734 565774
rect 240114 565454 240734 565538
rect 240114 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 240734 565454
rect 240114 529774 240734 565218
rect 240114 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 240734 529774
rect 240114 529454 240734 529538
rect 240114 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 240734 529454
rect 240114 493774 240734 529218
rect 240114 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 240734 493774
rect 240114 493454 240734 493538
rect 240114 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 240734 493454
rect 240114 457774 240734 493218
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 240114 421774 240734 457218
rect 240114 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 240734 421774
rect 240114 421454 240734 421538
rect 240114 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 240734 421454
rect 240114 385774 240734 421218
rect 240114 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 240734 385774
rect 240114 385454 240734 385538
rect 240114 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 240734 385454
rect 240114 349774 240734 385218
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 240114 313774 240734 349218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 605494 244454 640938
rect 243834 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 244454 605494
rect 243834 605174 244454 605258
rect 243834 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 244454 605174
rect 243834 569494 244454 604938
rect 243834 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 244454 569494
rect 243834 569174 244454 569258
rect 243834 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 244454 569174
rect 243834 533494 244454 568938
rect 243834 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 244454 533494
rect 243834 533174 244454 533258
rect 243834 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 244454 533174
rect 243834 497494 244454 532938
rect 243834 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 244454 497494
rect 243834 497174 244454 497258
rect 243834 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 244454 497174
rect 243834 461494 244454 496938
rect 243834 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 244454 461494
rect 243834 461174 244454 461258
rect 243834 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 244454 461174
rect 243834 425494 244454 460938
rect 243834 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 244454 425494
rect 243834 425174 244454 425258
rect 243834 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 244454 425174
rect 243834 389494 244454 424938
rect 243834 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 244454 389494
rect 243834 389174 244454 389258
rect 243834 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 244454 389174
rect 243834 353494 244454 388938
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 243834 317494 244454 352938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 246803 319020 246869 319021
rect 246803 318956 246804 319020
rect 246868 318956 246869 319020
rect 246803 318955 246869 318956
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 243491 315484 243557 315485
rect 243491 315420 243492 315484
rect 243556 315420 243557 315484
rect 243491 315419 243557 315420
rect 240114 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 240734 313774
rect 240114 313454 240734 313538
rect 240114 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 240734 313454
rect 238155 312900 238221 312901
rect 238155 312836 238156 312900
rect 238220 312836 238221 312900
rect 238155 312835 238221 312836
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 235211 289780 235277 289781
rect 235211 289716 235212 289780
rect 235276 289716 235277 289780
rect 235211 289715 235277 289716
rect 235214 239869 235274 289715
rect 235395 289644 235461 289645
rect 235395 289580 235396 289644
rect 235460 289580 235461 289644
rect 235395 289579 235461 289580
rect 234659 239868 234725 239869
rect 234659 239804 234660 239868
rect 234724 239804 234725 239868
rect 234659 239803 234725 239804
rect 235211 239868 235277 239869
rect 235211 239804 235212 239868
rect 235276 239804 235277 239868
rect 235211 239803 235277 239804
rect 234475 239596 234541 239597
rect 234475 239532 234476 239596
rect 234540 239532 234541 239596
rect 234475 239531 234541 239532
rect 234662 238645 234722 239803
rect 233923 238644 233989 238645
rect 233923 238580 233924 238644
rect 233988 238580 233989 238644
rect 233923 238579 233989 238580
rect 234659 238644 234725 238645
rect 234659 238580 234660 238644
rect 234724 238580 234725 238644
rect 234659 238579 234725 238580
rect 235214 236877 235274 239803
rect 235398 239733 235458 289579
rect 236394 274054 237014 309498
rect 238158 306917 238218 312835
rect 238339 312764 238405 312765
rect 238339 312700 238340 312764
rect 238404 312700 238405 312764
rect 238339 312699 238405 312700
rect 238155 306916 238221 306917
rect 238155 306852 238156 306916
rect 238220 306852 238221 306916
rect 238155 306851 238221 306852
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236131 239868 236197 239869
rect 236131 239804 236132 239868
rect 236196 239804 236197 239868
rect 236131 239803 236197 239804
rect 235395 239732 235461 239733
rect 235395 239668 235396 239732
rect 235460 239668 235461 239732
rect 235395 239667 235461 239668
rect 236134 239461 236194 239803
rect 236131 239460 236197 239461
rect 236131 239396 236132 239460
rect 236196 239396 236197 239460
rect 236131 239395 236197 239396
rect 236394 238054 237014 273498
rect 238342 253950 238402 312699
rect 238707 312628 238773 312629
rect 238707 312564 238708 312628
rect 238772 312564 238773 312628
rect 238707 312563 238773 312564
rect 238710 312490 238770 312563
rect 238526 312430 238770 312490
rect 238526 307050 238586 312430
rect 238526 306990 238954 307050
rect 238523 306916 238589 306917
rect 238523 306852 238524 306916
rect 238588 306852 238589 306916
rect 238523 306851 238589 306852
rect 238158 253890 238402 253950
rect 237235 240140 237301 240141
rect 237235 240076 237236 240140
rect 237300 240076 237301 240140
rect 237235 240075 237301 240076
rect 237238 238101 237298 240075
rect 238158 240005 238218 253890
rect 238339 240412 238405 240413
rect 238339 240348 238340 240412
rect 238404 240348 238405 240412
rect 238339 240347 238405 240348
rect 237419 240004 237485 240005
rect 237419 239940 237420 240004
rect 237484 239940 237485 240004
rect 237419 239939 237485 239940
rect 238155 240004 238221 240005
rect 238155 239940 238156 240004
rect 238220 239940 238221 240004
rect 238155 239939 238221 239940
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 237235 238100 237301 238101
rect 237235 238036 237236 238100
rect 237300 238036 237301 238100
rect 237235 238035 237301 238036
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 235211 236876 235277 236877
rect 235211 236812 235212 236876
rect 235276 236812 235277 236876
rect 235211 236811 235277 236812
rect 234291 235380 234357 235381
rect 234291 235316 234292 235380
rect 234356 235316 234357 235380
rect 234291 235315 234357 235316
rect 233739 227084 233805 227085
rect 233739 227020 233740 227084
rect 233804 227020 233805 227084
rect 233739 227019 233805 227020
rect 233742 193901 233802 227019
rect 234294 222733 234354 235315
rect 235763 234836 235829 234837
rect 235763 234772 235764 234836
rect 235828 234772 235829 234836
rect 235763 234771 235829 234772
rect 235579 234564 235645 234565
rect 235579 234500 235580 234564
rect 235644 234500 235645 234564
rect 235579 234499 235645 234500
rect 235582 224365 235642 234499
rect 235579 224364 235645 224365
rect 235579 224300 235580 224364
rect 235644 224300 235645 224364
rect 235579 224299 235645 224300
rect 234291 222732 234357 222733
rect 234291 222668 234292 222732
rect 234356 222668 234357 222732
rect 234291 222667 234357 222668
rect 234294 219450 234354 222667
rect 233926 219390 234354 219450
rect 233926 207637 233986 219390
rect 235766 218925 235826 234771
rect 235763 218924 235829 218925
rect 235763 218860 235764 218924
rect 235828 218860 235829 218924
rect 235763 218859 235829 218860
rect 235766 218109 235826 218859
rect 235763 218108 235829 218109
rect 235763 218044 235764 218108
rect 235828 218044 235829 218108
rect 235763 218043 235829 218044
rect 233923 207636 233989 207637
rect 233923 207572 233924 207636
rect 233988 207572 233989 207636
rect 233923 207571 233989 207572
rect 236394 202054 237014 237498
rect 237422 224501 237482 239939
rect 238342 239325 238402 240347
rect 238526 239869 238586 306851
rect 238894 306373 238954 306990
rect 238891 306372 238957 306373
rect 238891 306308 238892 306372
rect 238956 306308 238957 306372
rect 238891 306307 238957 306308
rect 239259 300116 239325 300117
rect 239259 300052 239260 300116
rect 239324 300052 239325 300116
rect 239259 300051 239325 300052
rect 238891 296852 238957 296853
rect 238891 296850 238892 296852
rect 238710 296790 238892 296850
rect 238710 296581 238770 296790
rect 238891 296788 238892 296790
rect 238956 296788 238957 296852
rect 238891 296787 238957 296788
rect 238707 296580 238773 296581
rect 238707 296516 238708 296580
rect 238772 296516 238773 296580
rect 238707 296515 238773 296516
rect 238891 290324 238957 290325
rect 238891 290260 238892 290324
rect 238956 290260 238957 290324
rect 238891 290259 238957 290260
rect 238894 253950 238954 290259
rect 238710 253890 238954 253950
rect 238523 239868 238589 239869
rect 238523 239804 238524 239868
rect 238588 239804 238589 239868
rect 238523 239803 238589 239804
rect 238710 239597 238770 253890
rect 239262 248430 239322 300051
rect 240114 277774 240734 313218
rect 241283 313036 241349 313037
rect 241283 312972 241284 313036
rect 241348 312972 241349 313036
rect 241283 312971 241349 312972
rect 240915 305692 240981 305693
rect 240915 305628 240916 305692
rect 240980 305628 240981 305692
rect 240915 305627 240981 305628
rect 240114 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 240734 277774
rect 240114 277454 240734 277538
rect 240114 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 240734 277454
rect 239568 259174 239888 259206
rect 239568 258938 239610 259174
rect 239846 258938 239888 259174
rect 239568 258854 239888 258938
rect 239568 258618 239610 258854
rect 239846 258618 239888 258854
rect 239568 258586 239888 258618
rect 238894 248370 239322 248430
rect 238894 239733 238954 248370
rect 240114 241774 240734 277218
rect 239075 241772 239141 241773
rect 239075 241708 239076 241772
rect 239140 241708 239141 241772
rect 239075 241707 239141 241708
rect 239078 239869 239138 241707
rect 240114 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 240734 241774
rect 240114 241454 240734 241538
rect 240114 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 240734 241454
rect 239075 239868 239141 239869
rect 239075 239804 239076 239868
rect 239140 239804 239141 239868
rect 239075 239803 239141 239804
rect 238891 239732 238957 239733
rect 238891 239668 238892 239732
rect 238956 239668 238957 239732
rect 238891 239667 238957 239668
rect 238707 239596 238773 239597
rect 238707 239532 238708 239596
rect 238772 239532 238773 239596
rect 238707 239531 238773 239532
rect 238339 239324 238405 239325
rect 238339 239260 238340 239324
rect 238404 239260 238405 239324
rect 238339 239259 238405 239260
rect 237419 224500 237485 224501
rect 237419 224436 237420 224500
rect 237484 224436 237485 224500
rect 237419 224435 237485 224436
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 233739 193900 233805 193901
rect 233739 193836 233740 193900
rect 233804 193836 233805 193900
rect 233739 193835 233805 193836
rect 233555 188324 233621 188325
rect 233555 188260 233556 188324
rect 233620 188260 233621 188324
rect 233555 188259 233621 188260
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 166054 237014 201498
rect 238894 199477 238954 239667
rect 239078 226949 239138 239803
rect 239443 239596 239509 239597
rect 239443 239532 239444 239596
rect 239508 239532 239509 239596
rect 239443 239531 239509 239532
rect 239075 226948 239141 226949
rect 239075 226884 239076 226948
rect 239140 226884 239141 226948
rect 239075 226883 239141 226884
rect 238891 199476 238957 199477
rect 238891 199412 238892 199476
rect 238956 199412 238957 199476
rect 238891 199411 238957 199412
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 236394 130054 237014 165498
rect 239446 156637 239506 239531
rect 240114 205774 240734 241218
rect 240918 239869 240978 305627
rect 240915 239868 240981 239869
rect 240915 239804 240916 239868
rect 240980 239804 240981 239868
rect 240915 239803 240981 239804
rect 240918 237965 240978 239803
rect 241286 239597 241346 312971
rect 242203 312356 242269 312357
rect 242203 312292 242204 312356
rect 242268 312292 242269 312356
rect 242203 312291 242269 312292
rect 242019 300388 242085 300389
rect 242019 300324 242020 300388
rect 242084 300324 242085 300388
rect 242019 300323 242085 300324
rect 242022 239869 242082 300323
rect 242019 239868 242085 239869
rect 242019 239804 242020 239868
rect 242084 239804 242085 239868
rect 242019 239803 242085 239804
rect 242206 239597 242266 312291
rect 243307 312220 243373 312221
rect 243307 312156 243308 312220
rect 243372 312156 243373 312220
rect 243307 312155 243373 312156
rect 242387 291820 242453 291821
rect 242387 291756 242388 291820
rect 242452 291756 242453 291820
rect 242387 291755 242453 291756
rect 242390 239733 242450 291755
rect 243123 240004 243189 240005
rect 243123 239940 243124 240004
rect 243188 239940 243189 240004
rect 243123 239939 243189 239940
rect 242755 239868 242821 239869
rect 242755 239804 242756 239868
rect 242820 239804 242821 239868
rect 242755 239803 242821 239804
rect 242387 239732 242453 239733
rect 242387 239668 242388 239732
rect 242452 239668 242453 239732
rect 242387 239667 242453 239668
rect 241283 239596 241349 239597
rect 241283 239532 241284 239596
rect 241348 239532 241349 239596
rect 241283 239531 241349 239532
rect 242203 239596 242269 239597
rect 242203 239532 242204 239596
rect 242268 239532 242269 239596
rect 242203 239531 242269 239532
rect 241651 239188 241717 239189
rect 241651 239124 241652 239188
rect 241716 239124 241717 239188
rect 241651 239123 241717 239124
rect 240915 237964 240981 237965
rect 240915 237900 240916 237964
rect 240980 237900 240981 237964
rect 240915 237899 240981 237900
rect 241654 235925 241714 239123
rect 241651 235924 241717 235925
rect 241651 235860 241652 235924
rect 241716 235860 241717 235924
rect 241651 235859 241717 235860
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 240114 169774 240734 205218
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 239443 156636 239509 156637
rect 239443 156572 239444 156636
rect 239508 156572 239509 156636
rect 239443 156571 239509 156572
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 94054 237014 129498
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 133774 240734 169218
rect 242206 141405 242266 239531
rect 242758 239050 242818 239803
rect 242574 238990 242818 239050
rect 242387 236740 242453 236741
rect 242387 236676 242388 236740
rect 242452 236676 242453 236740
rect 242387 236675 242453 236676
rect 242390 229805 242450 236675
rect 242387 229804 242453 229805
rect 242387 229740 242388 229804
rect 242452 229740 242453 229804
rect 242387 229739 242453 229740
rect 242390 204917 242450 229739
rect 242574 227357 242634 238990
rect 242755 238644 242821 238645
rect 242755 238580 242756 238644
rect 242820 238580 242821 238644
rect 242755 238579 242821 238580
rect 242758 232661 242818 238579
rect 243126 234565 243186 239939
rect 243310 239597 243370 312155
rect 243307 239596 243373 239597
rect 243307 239532 243308 239596
rect 243372 239532 243373 239596
rect 243307 239531 243373 239532
rect 243494 239461 243554 315419
rect 243834 281494 244454 316938
rect 246435 311404 246501 311405
rect 246435 311340 246436 311404
rect 246500 311340 246501 311404
rect 246435 311339 246501 311340
rect 245515 307732 245581 307733
rect 245515 307668 245516 307732
rect 245580 307668 245581 307732
rect 245515 307667 245581 307668
rect 245331 290596 245397 290597
rect 245331 290532 245332 290596
rect 245396 290532 245397 290596
rect 245331 290531 245397 290532
rect 243834 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 244454 281494
rect 243834 281174 244454 281258
rect 243834 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 244454 281174
rect 243834 245494 244454 280938
rect 245334 249810 245394 290531
rect 243834 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 244454 245494
rect 243834 245174 244454 245258
rect 243834 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 244454 245174
rect 243491 239460 243557 239461
rect 243491 239396 243492 239460
rect 243556 239396 243557 239460
rect 243491 239395 243557 239396
rect 243307 238644 243373 238645
rect 243307 238580 243308 238644
rect 243372 238580 243373 238644
rect 243307 238579 243373 238580
rect 243123 234564 243189 234565
rect 243123 234500 243124 234564
rect 243188 234500 243189 234564
rect 243123 234499 243189 234500
rect 242755 232660 242821 232661
rect 242755 232596 242756 232660
rect 242820 232596 242821 232660
rect 242755 232595 242821 232596
rect 242571 227356 242637 227357
rect 242571 227292 242572 227356
rect 242636 227292 242637 227356
rect 242571 227291 242637 227292
rect 242387 204916 242453 204917
rect 242387 204852 242388 204916
rect 242452 204852 242453 204916
rect 242387 204851 242453 204852
rect 242574 200701 242634 227291
rect 242758 220829 242818 232595
rect 242755 220828 242821 220829
rect 242755 220764 242756 220828
rect 242820 220764 242821 220828
rect 242755 220763 242821 220764
rect 243310 214573 243370 238579
rect 243494 228309 243554 239395
rect 243491 228308 243557 228309
rect 243491 228244 243492 228308
rect 243556 228244 243557 228308
rect 243491 228243 243557 228244
rect 243307 214572 243373 214573
rect 243307 214508 243308 214572
rect 243372 214508 243373 214572
rect 243307 214507 243373 214508
rect 243834 209494 244454 244938
rect 244966 249750 245394 249810
rect 244966 239733 245026 249750
rect 244963 239732 245029 239733
rect 244963 239668 244964 239732
rect 245028 239668 245029 239732
rect 244963 239667 245029 239668
rect 244966 211853 245026 239667
rect 245518 239597 245578 307667
rect 246438 249810 246498 311339
rect 246070 249750 246498 249810
rect 246070 239733 246130 249750
rect 246619 241500 246685 241501
rect 246619 241436 246620 241500
rect 246684 241436 246685 241500
rect 246619 241435 246685 241436
rect 246251 239868 246317 239869
rect 246251 239804 246252 239868
rect 246316 239804 246317 239868
rect 246251 239803 246317 239804
rect 246067 239732 246133 239733
rect 246067 239668 246068 239732
rect 246132 239668 246133 239732
rect 246067 239667 246133 239668
rect 245515 239596 245581 239597
rect 245515 239532 245516 239596
rect 245580 239532 245581 239596
rect 245515 239531 245581 239532
rect 245147 238644 245213 238645
rect 245147 238580 245148 238644
rect 245212 238580 245213 238644
rect 245147 238579 245213 238580
rect 245331 238644 245397 238645
rect 245331 238580 245332 238644
rect 245396 238580 245397 238644
rect 245331 238579 245397 238580
rect 245150 223141 245210 238579
rect 245147 223140 245213 223141
rect 245147 223076 245148 223140
rect 245212 223076 245213 223140
rect 245147 223075 245213 223076
rect 245334 222597 245394 238579
rect 245331 222596 245397 222597
rect 245331 222532 245332 222596
rect 245396 222532 245397 222596
rect 245331 222531 245397 222532
rect 244963 211852 245029 211853
rect 244963 211788 244964 211852
rect 245028 211788 245029 211852
rect 244963 211787 245029 211788
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 242571 200700 242637 200701
rect 242571 200636 242572 200700
rect 242636 200636 242637 200700
rect 242571 200635 242637 200636
rect 243834 173494 244454 208938
rect 245334 188325 245394 222531
rect 245331 188324 245397 188325
rect 245331 188260 245332 188324
rect 245396 188260 245397 188324
rect 245331 188259 245397 188260
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 242203 141404 242269 141405
rect 242203 141340 242204 141404
rect 242268 141340 242269 141404
rect 242203 141339 242269 141340
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 240114 97774 240734 133218
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 137494 244454 172938
rect 245518 166293 245578 239531
rect 246070 192541 246130 239667
rect 246254 213213 246314 239803
rect 246622 239597 246682 241435
rect 246806 239869 246866 318955
rect 253427 315620 253493 315621
rect 253427 315556 253428 315620
rect 253492 315556 253493 315620
rect 253427 315555 253493 315556
rect 249379 311812 249445 311813
rect 249379 311748 249380 311812
rect 249444 311748 249445 311812
rect 249379 311747 249445 311748
rect 247723 311676 247789 311677
rect 247723 311612 247724 311676
rect 247788 311612 247789 311676
rect 247723 311611 247789 311612
rect 247726 249810 247786 311611
rect 248091 311268 248157 311269
rect 248091 311204 248092 311268
rect 248156 311204 248157 311268
rect 248091 311203 248157 311204
rect 247907 297532 247973 297533
rect 247907 297468 247908 297532
rect 247972 297468 247973 297532
rect 247907 297467 247973 297468
rect 247542 249750 247786 249810
rect 247542 247050 247602 249750
rect 247358 246990 247602 247050
rect 246803 239868 246869 239869
rect 246803 239804 246804 239868
rect 246868 239804 246869 239868
rect 246803 239803 246869 239804
rect 246619 239596 246685 239597
rect 246619 239532 246620 239596
rect 246684 239532 246685 239596
rect 246619 239531 246685 239532
rect 246622 231165 246682 239531
rect 247358 239461 247418 246990
rect 247539 239868 247605 239869
rect 247539 239804 247540 239868
rect 247604 239804 247605 239868
rect 247539 239803 247605 239804
rect 247355 239460 247421 239461
rect 247355 239396 247356 239460
rect 247420 239396 247421 239460
rect 247355 239395 247421 239396
rect 246803 238644 246869 238645
rect 246803 238580 246804 238644
rect 246868 238580 246869 238644
rect 246803 238579 246869 238580
rect 246619 231164 246685 231165
rect 246619 231100 246620 231164
rect 246684 231100 246685 231164
rect 246619 231099 246685 231100
rect 246806 223413 246866 238579
rect 246803 223412 246869 223413
rect 246803 223348 246804 223412
rect 246868 223348 246869 223412
rect 246803 223347 246869 223348
rect 246251 213212 246317 213213
rect 246251 213148 246252 213212
rect 246316 213148 246317 213212
rect 246251 213147 246317 213148
rect 246067 192540 246133 192541
rect 246067 192476 246068 192540
rect 246132 192476 246133 192540
rect 246067 192475 246133 192476
rect 245515 166292 245581 166293
rect 245515 166228 245516 166292
rect 245580 166228 245581 166292
rect 245515 166227 245581 166228
rect 246806 152421 246866 223347
rect 247358 186965 247418 239395
rect 247542 199341 247602 239803
rect 247910 239733 247970 297467
rect 248094 239869 248154 311203
rect 249195 311132 249261 311133
rect 249195 311068 249196 311132
rect 249260 311068 249261 311132
rect 249195 311067 249261 311068
rect 249011 290052 249077 290053
rect 249011 289988 249012 290052
rect 249076 289988 249077 290052
rect 249011 289987 249077 289988
rect 248275 240684 248341 240685
rect 248275 240620 248276 240684
rect 248340 240620 248341 240684
rect 248275 240619 248341 240620
rect 248091 239868 248157 239869
rect 248091 239804 248092 239868
rect 248156 239804 248157 239868
rect 248091 239803 248157 239804
rect 248278 239733 248338 240619
rect 249014 239869 249074 289987
rect 249011 239868 249077 239869
rect 249011 239804 249012 239868
rect 249076 239804 249077 239868
rect 249011 239803 249077 239804
rect 247907 239732 247973 239733
rect 247907 239668 247908 239732
rect 247972 239668 247973 239732
rect 247907 239667 247973 239668
rect 248275 239732 248341 239733
rect 248275 239668 248276 239732
rect 248340 239668 248341 239732
rect 248275 239667 248341 239668
rect 247723 239596 247789 239597
rect 247723 239532 247724 239596
rect 247788 239532 247789 239596
rect 247723 239531 247789 239532
rect 247726 224229 247786 239531
rect 248275 238644 248341 238645
rect 248275 238580 248276 238644
rect 248340 238580 248341 238644
rect 248275 238579 248341 238580
rect 247723 224228 247789 224229
rect 247723 224164 247724 224228
rect 247788 224164 247789 224228
rect 247723 224163 247789 224164
rect 248278 223277 248338 238579
rect 248275 223276 248341 223277
rect 248275 223212 248276 223276
rect 248340 223212 248341 223276
rect 248275 223211 248341 223212
rect 247539 199340 247605 199341
rect 247539 199276 247540 199340
rect 247604 199276 247605 199340
rect 247539 199275 247605 199276
rect 247355 186964 247421 186965
rect 247355 186900 247356 186964
rect 247420 186900 247421 186964
rect 247355 186899 247421 186900
rect 246803 152420 246869 152421
rect 246803 152356 246804 152420
rect 246868 152356 246869 152420
rect 246803 152355 246869 152356
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 101494 244454 136938
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 248278 6085 248338 223211
rect 249014 178669 249074 239803
rect 249198 239461 249258 311067
rect 249382 239597 249442 311747
rect 249563 311540 249629 311541
rect 249563 311476 249564 311540
rect 249628 311476 249629 311540
rect 249563 311475 249629 311476
rect 249566 239733 249626 311475
rect 253243 310180 253309 310181
rect 253243 310116 253244 310180
rect 253308 310116 253309 310180
rect 253243 310115 253309 310116
rect 253059 310044 253125 310045
rect 253059 309980 253060 310044
rect 253124 309980 253125 310044
rect 253059 309979 253125 309980
rect 252139 309500 252205 309501
rect 252139 309436 252140 309500
rect 252204 309436 252205 309500
rect 252139 309435 252205 309436
rect 251587 300252 251653 300253
rect 251587 300188 251588 300252
rect 251652 300188 251653 300252
rect 251587 300187 251653 300188
rect 250483 290052 250549 290053
rect 250483 289988 250484 290052
rect 250548 289988 250549 290052
rect 250483 289987 250549 289988
rect 250299 289508 250365 289509
rect 250299 289444 250300 289508
rect 250364 289444 250365 289508
rect 250299 289443 250365 289444
rect 250302 239869 250362 289443
rect 250299 239868 250365 239869
rect 250299 239804 250300 239868
rect 250364 239804 250365 239868
rect 250299 239803 250365 239804
rect 249563 239732 249629 239733
rect 249563 239668 249564 239732
rect 249628 239668 249629 239732
rect 249563 239667 249629 239668
rect 249379 239596 249445 239597
rect 249379 239532 249380 239596
rect 249444 239532 249445 239596
rect 249379 239531 249445 239532
rect 249195 239460 249261 239461
rect 249195 239396 249196 239460
rect 249260 239396 249261 239460
rect 249195 239395 249261 239396
rect 249011 178668 249077 178669
rect 249011 178604 249012 178668
rect 249076 178604 249077 178668
rect 249011 178603 249077 178604
rect 249198 167653 249258 239395
rect 249379 238644 249445 238645
rect 249379 238580 249380 238644
rect 249444 238580 249445 238644
rect 249379 238579 249445 238580
rect 249382 222869 249442 238579
rect 249566 236197 249626 239667
rect 250115 238644 250181 238645
rect 250115 238580 250116 238644
rect 250180 238580 250181 238644
rect 250115 238579 250181 238580
rect 249563 236196 249629 236197
rect 249563 236132 249564 236196
rect 249628 236132 249629 236196
rect 249563 236131 249629 236132
rect 250118 226269 250178 238579
rect 250486 237965 250546 289987
rect 250667 289780 250733 289781
rect 250667 289716 250668 289780
rect 250732 289716 250733 289780
rect 250667 289715 250733 289716
rect 250670 239733 250730 289715
rect 251590 239869 251650 300187
rect 251771 289644 251837 289645
rect 251771 289580 251772 289644
rect 251836 289580 251837 289644
rect 251771 289579 251837 289580
rect 251035 239868 251101 239869
rect 251035 239804 251036 239868
rect 251100 239804 251101 239868
rect 251035 239803 251101 239804
rect 251587 239868 251653 239869
rect 251587 239804 251588 239868
rect 251652 239804 251653 239868
rect 251587 239803 251653 239804
rect 250667 239732 250733 239733
rect 250667 239668 250668 239732
rect 250732 239668 250733 239732
rect 250667 239667 250733 239668
rect 250483 237964 250549 237965
rect 250483 237900 250484 237964
rect 250548 237900 250549 237964
rect 250483 237899 250549 237900
rect 250670 236197 250730 239667
rect 250851 239460 250917 239461
rect 250851 239396 250852 239460
rect 250916 239396 250917 239460
rect 250851 239395 250917 239396
rect 250667 236196 250733 236197
rect 250667 236132 250668 236196
rect 250732 236132 250733 236196
rect 250667 236131 250733 236132
rect 250115 226268 250181 226269
rect 250115 226204 250116 226268
rect 250180 226204 250181 226268
rect 250115 226203 250181 226204
rect 250854 223005 250914 239395
rect 250851 223004 250917 223005
rect 250851 222940 250852 223004
rect 250916 222940 250917 223004
rect 250851 222939 250917 222940
rect 249379 222868 249445 222869
rect 249379 222804 249380 222868
rect 249444 222804 249445 222868
rect 249379 222803 249445 222804
rect 249382 197981 249442 222803
rect 250854 202197 250914 222939
rect 250851 202196 250917 202197
rect 250851 202132 250852 202196
rect 250916 202132 250917 202196
rect 250851 202131 250917 202132
rect 249379 197980 249445 197981
rect 249379 197916 249380 197980
rect 249444 197916 249445 197980
rect 249379 197915 249445 197916
rect 249195 167652 249261 167653
rect 249195 167588 249196 167652
rect 249260 167588 249261 167652
rect 249195 167587 249261 167588
rect 251038 138685 251098 239803
rect 251035 138684 251101 138685
rect 251035 138620 251036 138684
rect 251100 138620 251101 138684
rect 251035 138619 251101 138620
rect 248275 6084 248341 6085
rect 248275 6020 248276 6084
rect 248340 6020 248341 6084
rect 248275 6019 248341 6020
rect 251590 3637 251650 239803
rect 251774 239597 251834 289579
rect 252142 239733 252202 309435
rect 252875 294540 252941 294541
rect 252875 294476 252876 294540
rect 252940 294476 252941 294540
rect 252875 294475 252941 294476
rect 252878 239869 252938 294475
rect 252875 239868 252941 239869
rect 252875 239804 252876 239868
rect 252940 239804 252941 239868
rect 252875 239803 252941 239804
rect 251955 239732 252021 239733
rect 251955 239668 251956 239732
rect 252020 239668 252021 239732
rect 251955 239667 252021 239668
rect 252139 239732 252205 239733
rect 252139 239668 252140 239732
rect 252204 239668 252205 239732
rect 252139 239667 252205 239668
rect 251771 239596 251837 239597
rect 251771 239532 251772 239596
rect 251836 239532 251837 239596
rect 251771 239531 251837 239532
rect 251958 221645 252018 239667
rect 251955 221644 252021 221645
rect 251955 221580 251956 221644
rect 252020 221580 252021 221644
rect 251955 221579 252021 221580
rect 251587 3636 251653 3637
rect 251587 3572 251588 3636
rect 251652 3572 251653 3636
rect 251587 3571 251653 3572
rect 252142 3501 252202 239667
rect 253062 239597 253122 309979
rect 253246 239733 253306 310115
rect 253243 239732 253309 239733
rect 253243 239668 253244 239732
rect 253308 239668 253309 239732
rect 253243 239667 253309 239668
rect 253059 239596 253125 239597
rect 253059 239594 253060 239596
rect 252878 239534 253060 239594
rect 252878 231870 252938 239534
rect 253059 239532 253060 239534
rect 253124 239532 253125 239596
rect 253059 239531 253125 239532
rect 253059 238644 253125 238645
rect 253059 238580 253060 238644
rect 253124 238580 253125 238644
rect 253059 238579 253125 238580
rect 252694 231810 252938 231870
rect 252694 6901 252754 231810
rect 253062 228717 253122 238579
rect 253059 228716 253125 228717
rect 253059 228652 253060 228716
rect 253124 228652 253125 228716
rect 253059 228651 253125 228652
rect 252691 6900 252757 6901
rect 252691 6836 252692 6900
rect 252756 6836 252757 6900
rect 252691 6835 252757 6836
rect 253246 6765 253306 239667
rect 253430 239189 253490 315555
rect 253794 291454 254414 326898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 254715 310316 254781 310317
rect 254715 310252 254716 310316
rect 254780 310252 254781 310316
rect 254715 310251 254781 310252
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253427 239188 253493 239189
rect 253427 239124 253428 239188
rect 253492 239124 253493 239188
rect 253427 239123 253493 239124
rect 253794 219454 254414 254898
rect 254718 239597 254778 310251
rect 257514 295174 258134 330618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 259315 308548 259381 308549
rect 259315 308484 259316 308548
rect 259380 308484 259381 308548
rect 259315 308483 259381 308484
rect 259131 308412 259197 308413
rect 259131 308348 259132 308412
rect 259196 308348 259197 308412
rect 259131 308347 259197 308348
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257107 290460 257173 290461
rect 257107 290396 257108 290460
rect 257172 290396 257173 290460
rect 257107 290395 257173 290396
rect 255451 290052 255517 290053
rect 255451 289988 255452 290052
rect 255516 289988 255517 290052
rect 255451 289987 255517 289988
rect 254928 255454 255248 255486
rect 254928 255218 254970 255454
rect 255206 255218 255248 255454
rect 254928 255134 255248 255218
rect 254928 254898 254970 255134
rect 255206 254898 255248 255134
rect 254928 254866 255248 254898
rect 255454 239597 255514 289987
rect 255635 289780 255701 289781
rect 255635 289716 255636 289780
rect 255700 289716 255701 289780
rect 255635 289715 255701 289716
rect 255638 239869 255698 289715
rect 255819 289644 255885 289645
rect 255819 289580 255820 289644
rect 255884 289580 255885 289644
rect 255819 289579 255885 289580
rect 255635 239868 255701 239869
rect 255635 239804 255636 239868
rect 255700 239804 255701 239868
rect 255635 239803 255701 239804
rect 255822 239597 255882 289579
rect 256187 287740 256253 287741
rect 256187 287676 256188 287740
rect 256252 287676 256253 287740
rect 256187 287675 256253 287676
rect 256190 239869 256250 287675
rect 256187 239868 256253 239869
rect 256187 239866 256188 239868
rect 256006 239806 256188 239866
rect 254715 239596 254781 239597
rect 254715 239532 254716 239596
rect 254780 239532 254781 239596
rect 254715 239531 254781 239532
rect 255451 239596 255517 239597
rect 255451 239532 255452 239596
rect 255516 239532 255517 239596
rect 255451 239531 255517 239532
rect 255819 239596 255885 239597
rect 255819 239532 255820 239596
rect 255884 239532 255885 239596
rect 255819 239531 255885 239532
rect 254718 237965 254778 239531
rect 254715 237964 254781 237965
rect 254715 237900 254716 237964
rect 254780 237900 254781 237964
rect 254715 237899 254781 237900
rect 255083 236060 255149 236061
rect 255083 235996 255084 236060
rect 255148 235996 255149 236060
rect 255083 235995 255149 235996
rect 254899 235924 254965 235925
rect 254899 235860 254900 235924
rect 254964 235860 254965 235924
rect 254899 235859 254965 235860
rect 254902 223821 254962 235859
rect 255086 225997 255146 235995
rect 255083 225996 255149 225997
rect 255083 225932 255084 225996
rect 255148 225932 255149 225996
rect 255083 225931 255149 225932
rect 254899 223820 254965 223821
rect 254899 223756 254900 223820
rect 254964 223756 254965 223820
rect 254899 223755 254965 223756
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 255086 156637 255146 225931
rect 255083 156636 255149 156637
rect 255083 156572 255084 156636
rect 255148 156572 255149 156636
rect 255083 156571 255149 156572
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253243 6764 253309 6765
rect 253243 6700 253244 6764
rect 253308 6700 253309 6764
rect 253243 6699 253309 6700
rect 252139 3500 252205 3501
rect 252139 3436 252140 3500
rect 252204 3436 252205 3500
rect 252139 3435 252205 3436
rect 253794 3454 254414 38898
rect 256006 6357 256066 239806
rect 256187 239804 256188 239806
rect 256252 239804 256253 239868
rect 256187 239803 256253 239804
rect 256923 239868 256989 239869
rect 256923 239804 256924 239868
rect 256988 239804 256989 239868
rect 256923 239803 256989 239804
rect 256739 239732 256805 239733
rect 256739 239730 256740 239732
rect 256558 239670 256740 239730
rect 256371 239596 256437 239597
rect 256371 239532 256372 239596
rect 256436 239532 256437 239596
rect 256371 239531 256437 239532
rect 256187 237964 256253 237965
rect 256187 237900 256188 237964
rect 256252 237900 256253 237964
rect 256187 237899 256253 237900
rect 256190 221509 256250 237899
rect 256187 221508 256253 221509
rect 256187 221444 256188 221508
rect 256252 221444 256253 221508
rect 256187 221443 256253 221444
rect 256190 6629 256250 221443
rect 256187 6628 256253 6629
rect 256187 6564 256188 6628
rect 256252 6564 256253 6628
rect 256187 6563 256253 6564
rect 256374 6493 256434 239531
rect 256558 232933 256618 239670
rect 256739 239668 256740 239670
rect 256804 239668 256805 239732
rect 256739 239667 256805 239668
rect 256739 239460 256805 239461
rect 256739 239396 256740 239460
rect 256804 239396 256805 239460
rect 256739 239395 256805 239396
rect 256742 237693 256802 239395
rect 256739 237692 256805 237693
rect 256739 237628 256740 237692
rect 256804 237628 256805 237692
rect 256739 237627 256805 237628
rect 256739 235244 256805 235245
rect 256739 235180 256740 235244
rect 256804 235180 256805 235244
rect 256739 235179 256805 235180
rect 256555 232932 256621 232933
rect 256555 232868 256556 232932
rect 256620 232868 256621 232932
rect 256555 232867 256621 232868
rect 256742 224093 256802 235179
rect 256739 224092 256805 224093
rect 256739 224028 256740 224092
rect 256804 224028 256805 224092
rect 256739 224027 256805 224028
rect 256742 169013 256802 224027
rect 256926 221373 256986 239803
rect 257110 239597 257170 290395
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257107 239596 257173 239597
rect 257107 239532 257108 239596
rect 257172 239532 257173 239596
rect 257107 239531 257173 239532
rect 257107 236740 257173 236741
rect 257107 236676 257108 236740
rect 257172 236676 257173 236740
rect 257107 236675 257173 236676
rect 256923 221372 256989 221373
rect 256923 221308 256924 221372
rect 256988 221308 256989 221372
rect 256923 221307 256989 221308
rect 256739 169012 256805 169013
rect 256739 168948 256740 169012
rect 256804 168948 256805 169012
rect 256739 168947 256805 168948
rect 256926 151061 256986 221307
rect 257110 218653 257170 236675
rect 257514 223174 258134 258618
rect 258763 241636 258829 241637
rect 258763 241572 258764 241636
rect 258828 241572 258829 241636
rect 258763 241571 258829 241572
rect 258766 239597 258826 241571
rect 258947 239868 259013 239869
rect 258947 239804 258948 239868
rect 259012 239804 259013 239868
rect 258947 239803 259013 239804
rect 258763 239596 258829 239597
rect 258763 239532 258764 239596
rect 258828 239532 258829 239596
rect 258763 239531 258829 239532
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257107 218652 257173 218653
rect 257107 218588 257108 218652
rect 257172 218588 257173 218652
rect 257107 218587 257173 218588
rect 256923 151060 256989 151061
rect 256923 150996 256924 151060
rect 256988 150996 256989 151060
rect 256923 150995 256989 150996
rect 257110 15877 257170 218587
rect 257514 187174 258134 222618
rect 258950 218517 259010 239803
rect 259134 239461 259194 308347
rect 259318 240005 259378 308483
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260603 290868 260669 290869
rect 260603 290804 260604 290868
rect 260668 290804 260669 290868
rect 260603 290803 260669 290804
rect 259315 240004 259381 240005
rect 259315 239940 259316 240004
rect 259380 239940 259381 240004
rect 259315 239939 259381 239940
rect 259131 239460 259197 239461
rect 259131 239396 259132 239460
rect 259196 239396 259197 239460
rect 259131 239395 259197 239396
rect 258947 218516 259013 218517
rect 258947 218452 258948 218516
rect 259012 218452 259013 218516
rect 258947 218451 259013 218452
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 258950 146981 259010 218451
rect 258947 146980 259013 146981
rect 258947 146916 258948 146980
rect 259012 146916 259013 146980
rect 258947 146915 259013 146916
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257107 15876 257173 15877
rect 257107 15812 257108 15876
rect 257172 15812 257173 15876
rect 257107 15811 257173 15812
rect 257514 7174 258134 42618
rect 259134 25533 259194 239395
rect 259131 25532 259197 25533
rect 259131 25468 259132 25532
rect 259196 25468 259197 25532
rect 259131 25467 259197 25468
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 256371 6492 256437 6493
rect 256371 6428 256372 6492
rect 256436 6428 256437 6492
rect 256371 6427 256437 6428
rect 256003 6356 256069 6357
rect 256003 6292 256004 6356
rect 256068 6292 256069 6356
rect 256003 6291 256069 6292
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 -1306 258134 6618
rect 259318 6221 259378 239939
rect 260606 239597 260666 290803
rect 261234 262894 261854 298338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 263547 291548 263613 291549
rect 263547 291484 263548 291548
rect 263612 291484 263613 291548
rect 263547 291483 263613 291484
rect 263550 287061 263610 291483
rect 263547 287060 263613 287061
rect 263547 286996 263548 287060
rect 263612 286996 263613 287060
rect 263547 286995 263613 286996
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 260971 242044 261037 242045
rect 260971 241980 260972 242044
rect 261036 241980 261037 242044
rect 260971 241979 261037 241980
rect 260787 239868 260853 239869
rect 260787 239804 260788 239868
rect 260852 239804 260853 239868
rect 260787 239803 260853 239804
rect 260603 239596 260669 239597
rect 260603 239532 260604 239596
rect 260668 239532 260669 239596
rect 260603 239531 260669 239532
rect 260235 239324 260301 239325
rect 260235 239260 260236 239324
rect 260300 239260 260301 239324
rect 260235 239259 260301 239260
rect 260051 235244 260117 235245
rect 260051 235180 260052 235244
rect 260116 235180 260117 235244
rect 260051 235179 260117 235180
rect 260054 219061 260114 235179
rect 260238 224637 260298 239259
rect 260419 237556 260485 237557
rect 260419 237492 260420 237556
rect 260484 237492 260485 237556
rect 260419 237491 260485 237492
rect 260422 228989 260482 237491
rect 260419 228988 260485 228989
rect 260419 228924 260420 228988
rect 260484 228924 260485 228988
rect 260419 228923 260485 228924
rect 260235 224636 260301 224637
rect 260235 224572 260236 224636
rect 260300 224572 260301 224636
rect 260235 224571 260301 224572
rect 260051 219060 260117 219061
rect 260051 218996 260052 219060
rect 260116 218996 260117 219060
rect 260051 218995 260117 218996
rect 260054 218109 260114 218995
rect 260051 218108 260117 218109
rect 260051 218044 260052 218108
rect 260116 218044 260117 218108
rect 260051 218043 260117 218044
rect 259315 6220 259381 6221
rect 259315 6156 259316 6220
rect 259380 6156 259381 6220
rect 259315 6155 259381 6156
rect 260606 3365 260666 239531
rect 260790 236741 260850 239803
rect 260974 239597 261034 241979
rect 260971 239596 261037 239597
rect 260971 239532 260972 239596
rect 261036 239532 261037 239596
rect 260971 239531 261037 239532
rect 260787 236740 260853 236741
rect 260787 236676 260788 236740
rect 260852 236676 260853 236740
rect 260787 236675 260853 236676
rect 261234 226894 261854 262338
rect 264954 266614 265574 302058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 268674 594334 269294 629778
rect 268674 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 269294 594334
rect 268674 594014 269294 594098
rect 268674 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 269294 594014
rect 268674 558334 269294 593778
rect 268674 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 269294 558334
rect 268674 558014 269294 558098
rect 268674 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 269294 558014
rect 268674 522334 269294 557778
rect 268674 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 269294 522334
rect 268674 522014 269294 522098
rect 268674 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 269294 522014
rect 268674 486334 269294 521778
rect 268674 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 269294 486334
rect 268674 486014 269294 486098
rect 268674 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 269294 486014
rect 268674 450334 269294 485778
rect 268674 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 269294 450334
rect 268674 450014 269294 450098
rect 268674 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 269294 450014
rect 268674 414334 269294 449778
rect 268674 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 269294 414334
rect 268674 414014 269294 414098
rect 268674 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 269294 414014
rect 268674 378334 269294 413778
rect 268674 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 269294 378334
rect 268674 378014 269294 378098
rect 268674 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 269294 378014
rect 268674 342334 269294 377778
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 268674 306334 269294 341778
rect 268674 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 269294 306334
rect 268674 306014 269294 306098
rect 268674 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 269294 306014
rect 266491 271148 266557 271149
rect 266491 271084 266492 271148
rect 266556 271084 266557 271148
rect 266491 271083 266557 271084
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 263731 258772 263797 258773
rect 263731 258708 263732 258772
rect 263796 258708 263797 258772
rect 263731 258707 263797 258708
rect 263547 244900 263613 244901
rect 263547 244836 263548 244900
rect 263612 244836 263613 244900
rect 263547 244835 263613 244836
rect 262075 239868 262141 239869
rect 262075 239804 262076 239868
rect 262140 239804 262141 239868
rect 262075 239803 262141 239804
rect 262078 239325 262138 239803
rect 263550 239733 263610 244835
rect 263734 244082 263794 258707
rect 264099 247756 264165 247757
rect 264099 247692 264100 247756
rect 264164 247692 264165 247756
rect 264099 247691 264165 247692
rect 263734 244022 263978 244082
rect 263731 242180 263797 242181
rect 263731 242116 263732 242180
rect 263796 242116 263797 242180
rect 263731 242115 263797 242116
rect 262627 239732 262693 239733
rect 262627 239668 262628 239732
rect 262692 239730 262693 239732
rect 263547 239732 263613 239733
rect 262692 239670 262874 239730
rect 262692 239668 262693 239670
rect 262627 239667 262693 239668
rect 262627 239596 262693 239597
rect 262627 239532 262628 239596
rect 262692 239532 262693 239596
rect 262627 239531 262693 239532
rect 262075 239324 262141 239325
rect 262075 239260 262076 239324
rect 262140 239260 262141 239324
rect 262075 239259 262141 239260
rect 262075 239188 262141 239189
rect 262075 239124 262076 239188
rect 262140 239124 262141 239188
rect 262075 239123 262141 239124
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 262078 224365 262138 239123
rect 262075 224364 262141 224365
rect 262075 224300 262076 224364
rect 262140 224300 262141 224364
rect 262075 224299 262141 224300
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 260603 3364 260669 3365
rect 260603 3300 260604 3364
rect 260668 3300 260669 3364
rect 260603 3299 260669 3300
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 -2266 261854 10338
rect 262630 10301 262690 239531
rect 262814 224501 262874 239670
rect 263547 239668 263548 239732
rect 263612 239668 263613 239732
rect 263547 239667 263613 239668
rect 263547 239324 263613 239325
rect 263547 239260 263548 239324
rect 263612 239322 263613 239324
rect 263734 239322 263794 242115
rect 263918 240005 263978 244022
rect 263915 240004 263981 240005
rect 263915 239940 263916 240004
rect 263980 239940 263981 240004
rect 263915 239939 263981 239940
rect 263612 239262 263794 239322
rect 263612 239260 263613 239262
rect 263547 239259 263613 239260
rect 263179 235244 263245 235245
rect 263179 235180 263180 235244
rect 263244 235180 263245 235244
rect 263179 235179 263245 235180
rect 263182 225861 263242 235179
rect 263918 231870 263978 239939
rect 264102 238237 264162 247691
rect 264467 243948 264533 243949
rect 264467 243884 264468 243948
rect 264532 243884 264533 243948
rect 264467 243883 264533 243884
rect 264283 242316 264349 242317
rect 264283 242252 264284 242316
rect 264348 242252 264349 242316
rect 264283 242251 264349 242252
rect 264286 239869 264346 242251
rect 264283 239868 264349 239869
rect 264283 239804 264284 239868
rect 264348 239804 264349 239868
rect 264283 239803 264349 239804
rect 264286 238509 264346 239803
rect 264470 239733 264530 243883
rect 264651 241908 264717 241909
rect 264651 241844 264652 241908
rect 264716 241844 264717 241908
rect 264651 241843 264717 241844
rect 264467 239732 264533 239733
rect 264467 239668 264468 239732
rect 264532 239668 264533 239732
rect 264467 239667 264533 239668
rect 264654 239189 264714 241843
rect 264651 239188 264717 239189
rect 264651 239124 264652 239188
rect 264716 239124 264717 239188
rect 264651 239123 264717 239124
rect 264283 238508 264349 238509
rect 264283 238444 264284 238508
rect 264348 238444 264349 238508
rect 264283 238443 264349 238444
rect 264099 238236 264165 238237
rect 264099 238172 264100 238236
rect 264164 238172 264165 238236
rect 264099 238171 264165 238172
rect 264467 237964 264533 237965
rect 264467 237900 264468 237964
rect 264532 237900 264533 237964
rect 264467 237899 264533 237900
rect 263734 231810 263978 231870
rect 263179 225860 263245 225861
rect 263179 225796 263180 225860
rect 263244 225796 263245 225860
rect 263179 225795 263245 225796
rect 262811 224500 262877 224501
rect 262811 224436 262812 224500
rect 262876 224436 262877 224500
rect 262811 224435 262877 224436
rect 262814 219450 262874 224435
rect 262814 219390 263058 219450
rect 262998 191045 263058 219390
rect 262995 191044 263061 191045
rect 262995 190980 262996 191044
rect 263060 190980 263061 191044
rect 262995 190979 263061 190980
rect 263182 189685 263242 225795
rect 263179 189684 263245 189685
rect 263179 189620 263180 189684
rect 263244 189620 263245 189684
rect 263179 189619 263245 189620
rect 263734 182885 263794 231810
rect 264470 221237 264530 237899
rect 264954 230614 265574 266058
rect 266123 245036 266189 245037
rect 266123 244972 266124 245036
rect 266188 244972 266189 245036
rect 266123 244971 266189 244972
rect 265939 240956 266005 240957
rect 265939 240892 265940 240956
rect 266004 240892 266005 240956
rect 265939 240891 266005 240892
rect 265942 239869 266002 240891
rect 265939 239868 266005 239869
rect 265939 239804 265940 239868
rect 266004 239804 266005 239868
rect 265939 239803 266005 239804
rect 266126 239733 266186 244971
rect 266494 240005 266554 271083
rect 268674 270334 269294 305778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 272394 598054 273014 633498
rect 272394 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 273014 598054
rect 272394 597734 273014 597818
rect 272394 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 273014 597734
rect 272394 562054 273014 597498
rect 272394 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 273014 562054
rect 272394 561734 273014 561818
rect 272394 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 273014 561734
rect 272394 526054 273014 561498
rect 272394 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 273014 526054
rect 272394 525734 273014 525818
rect 272394 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 273014 525734
rect 272394 490054 273014 525498
rect 272394 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 273014 490054
rect 272394 489734 273014 489818
rect 272394 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 273014 489734
rect 272394 454054 273014 489498
rect 272394 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 273014 454054
rect 272394 453734 273014 453818
rect 272394 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 273014 453734
rect 272394 418054 273014 453498
rect 272394 417818 272426 418054
rect 272662 417818 272746 418054
rect 272982 417818 273014 418054
rect 272394 417734 273014 417818
rect 272394 417498 272426 417734
rect 272662 417498 272746 417734
rect 272982 417498 273014 417734
rect 272394 382054 273014 417498
rect 272394 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 273014 382054
rect 272394 381734 273014 381818
rect 272394 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 273014 381734
rect 272394 346054 273014 381498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 276114 601774 276734 637218
rect 276114 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 276734 601774
rect 276114 601454 276734 601538
rect 276114 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 276734 601454
rect 276114 565774 276734 601218
rect 276114 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 276734 565774
rect 276114 565454 276734 565538
rect 276114 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 276734 565454
rect 276114 529774 276734 565218
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 276114 493774 276734 529218
rect 276114 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 276734 493774
rect 276114 493454 276734 493538
rect 276114 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 276734 493454
rect 276114 457774 276734 493218
rect 276114 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 276734 457774
rect 276114 457454 276734 457538
rect 276114 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 276734 457454
rect 276114 421774 276734 457218
rect 276114 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 276734 421774
rect 276114 421454 276734 421538
rect 276114 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 276734 421454
rect 276114 385774 276734 421218
rect 276114 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 276734 385774
rect 276114 385454 276734 385538
rect 276114 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 276734 385454
rect 275323 375596 275389 375597
rect 275323 375532 275324 375596
rect 275388 375532 275389 375596
rect 275323 375531 275389 375532
rect 275139 375460 275205 375461
rect 275139 375396 275140 375460
rect 275204 375396 275205 375460
rect 275139 375395 275205 375396
rect 272394 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 273014 346054
rect 272394 345734 273014 345818
rect 272394 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 273014 345734
rect 272394 310054 273014 345498
rect 272394 309818 272426 310054
rect 272662 309818 272746 310054
rect 272982 309818 273014 310054
rect 272394 309734 273014 309818
rect 272394 309498 272426 309734
rect 272662 309498 272746 309734
rect 272982 309498 273014 309734
rect 269619 289916 269685 289917
rect 269619 289852 269620 289916
rect 269684 289852 269685 289916
rect 269619 289851 269685 289852
rect 268674 270098 268706 270334
rect 268942 270098 269026 270334
rect 269262 270098 269294 270334
rect 268674 270014 269294 270098
rect 268674 269778 268706 270014
rect 268942 269778 269026 270014
rect 269262 269778 269294 270014
rect 267411 258908 267477 258909
rect 267411 258844 267412 258908
rect 267476 258844 267477 258908
rect 267411 258843 267477 258844
rect 266491 240004 266557 240005
rect 266491 239940 266492 240004
rect 266556 239940 266557 240004
rect 266491 239939 266557 239940
rect 267414 239869 267474 258843
rect 267595 244220 267661 244221
rect 267595 244156 267596 244220
rect 267660 244156 267661 244220
rect 267595 244155 267661 244156
rect 267598 240005 267658 244155
rect 267595 240004 267661 240005
rect 267595 239940 267596 240004
rect 267660 239940 267661 240004
rect 267595 239939 267661 239940
rect 267411 239868 267477 239869
rect 267411 239804 267412 239868
rect 267476 239804 267477 239868
rect 267411 239803 267477 239804
rect 265939 239732 266005 239733
rect 265939 239668 265940 239732
rect 266004 239668 266005 239732
rect 265939 239667 266005 239668
rect 266123 239732 266189 239733
rect 266123 239668 266124 239732
rect 266188 239668 266189 239732
rect 266123 239667 266189 239668
rect 265942 239189 266002 239667
rect 265939 239188 266005 239189
rect 265939 239124 265940 239188
rect 266004 239124 266005 239188
rect 265939 239123 266005 239124
rect 266126 231029 266186 239667
rect 267598 238373 267658 239939
rect 267595 238372 267661 238373
rect 267595 238308 267596 238372
rect 267660 238308 267661 238372
rect 267595 238307 267661 238308
rect 268674 234334 269294 269778
rect 268674 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 269294 234334
rect 268674 234014 269294 234098
rect 268674 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 269294 234014
rect 266123 231028 266189 231029
rect 266123 230964 266124 231028
rect 266188 230964 266189 231028
rect 266123 230963 266189 230964
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264467 221236 264533 221237
rect 264467 221172 264468 221236
rect 264532 221172 264533 221236
rect 264467 221171 264533 221172
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263731 182884 263797 182885
rect 263731 182820 263732 182884
rect 263796 182820 263797 182884
rect 263731 182819 263797 182820
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 262627 10300 262693 10301
rect 262627 10236 262628 10300
rect 262692 10236 262693 10300
rect 262627 10235 262693 10236
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 198334 269294 233778
rect 268674 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 269294 198334
rect 268674 198014 269294 198098
rect 268674 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 269294 198014
rect 268674 162334 269294 197778
rect 268674 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 269294 162334
rect 268674 162014 269294 162098
rect 268674 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 269294 162014
rect 268674 126334 269294 161778
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 90334 269294 125778
rect 269622 125629 269682 289851
rect 272394 274054 273014 309498
rect 275142 292093 275202 375395
rect 275326 294813 275386 375531
rect 276114 349774 276734 385218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 605494 280454 640938
rect 279834 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 280454 605494
rect 279834 605174 280454 605258
rect 279834 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 280454 605174
rect 279834 569494 280454 604938
rect 279834 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 280454 569494
rect 279834 569174 280454 569258
rect 279834 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 280454 569174
rect 279834 533494 280454 568938
rect 279834 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 280454 533494
rect 279834 533174 280454 533258
rect 279834 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 280454 533174
rect 279834 497494 280454 532938
rect 279834 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 280454 497494
rect 279834 497174 280454 497258
rect 279834 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 280454 497174
rect 279834 461494 280454 496938
rect 279834 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 280454 461494
rect 279834 461174 280454 461258
rect 279834 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 280454 461174
rect 279834 425494 280454 460938
rect 279834 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 280454 425494
rect 279834 425174 280454 425258
rect 279834 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 280454 425174
rect 279834 389494 280454 424938
rect 279834 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 280454 389494
rect 279834 389174 280454 389258
rect 279834 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 280454 389174
rect 277899 375732 277965 375733
rect 277899 375668 277900 375732
rect 277964 375668 277965 375732
rect 277899 375667 277965 375668
rect 276114 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 276734 349774
rect 276114 349454 276734 349538
rect 276114 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 276734 349454
rect 276114 313774 276734 349218
rect 276114 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 276734 313774
rect 276114 313454 276734 313538
rect 276114 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 276734 313454
rect 275323 294812 275389 294813
rect 275323 294748 275324 294812
rect 275388 294748 275389 294812
rect 275323 294747 275389 294748
rect 275139 292092 275205 292093
rect 275139 292028 275140 292092
rect 275204 292028 275205 292092
rect 275139 292027 275205 292028
rect 272394 273818 272426 274054
rect 272662 273818 272746 274054
rect 272982 273818 273014 274054
rect 272394 273734 273014 273818
rect 272394 273498 272426 273734
rect 272662 273498 272746 273734
rect 272982 273498 273014 273734
rect 272394 238054 273014 273498
rect 272394 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 273014 238054
rect 272394 237734 273014 237818
rect 272394 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 273014 237734
rect 272394 202054 273014 237498
rect 272394 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 273014 202054
rect 272394 201734 273014 201818
rect 272394 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 273014 201734
rect 272394 166054 273014 201498
rect 272394 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 273014 166054
rect 272394 165734 273014 165818
rect 272394 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 273014 165734
rect 272394 130054 273014 165498
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 269619 125628 269685 125629
rect 269619 125564 269620 125628
rect 269684 125564 269685 125628
rect 269619 125563 269685 125564
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 268674 54334 269294 89778
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 94054 273014 129498
rect 272394 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 273014 94054
rect 272394 93734 273014 93818
rect 272394 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 273014 93734
rect 272394 58054 273014 93498
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 277774 276734 313218
rect 277902 293317 277962 375667
rect 278083 374236 278149 374237
rect 278083 374172 278084 374236
rect 278148 374172 278149 374236
rect 278083 374171 278149 374172
rect 277899 293316 277965 293317
rect 277899 293252 277900 293316
rect 277964 293252 277965 293316
rect 277899 293251 277965 293252
rect 278086 293181 278146 374171
rect 279834 353494 280454 388938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 285627 371924 285693 371925
rect 285627 371860 285628 371924
rect 285692 371860 285693 371924
rect 285627 371859 285693 371860
rect 283787 369612 283853 369613
rect 283787 369548 283788 369612
rect 283852 369548 283853 369612
rect 283787 369547 283853 369548
rect 283051 369476 283117 369477
rect 283051 369412 283052 369476
rect 283116 369412 283117 369476
rect 283051 369411 283117 369412
rect 282683 369204 282749 369205
rect 282683 369140 282684 369204
rect 282748 369140 282749 369204
rect 282683 369139 282749 369140
rect 281395 360228 281461 360229
rect 281395 360164 281396 360228
rect 281460 360164 281461 360228
rect 281395 360163 281461 360164
rect 279834 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 280454 353494
rect 279834 353174 280454 353258
rect 279834 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 280454 353174
rect 279834 317494 280454 352938
rect 279834 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 280454 317494
rect 279834 317174 280454 317258
rect 279834 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 280454 317174
rect 278083 293180 278149 293181
rect 278083 293116 278084 293180
rect 278148 293116 278149 293180
rect 278083 293115 278149 293116
rect 276114 277538 276146 277774
rect 276382 277538 276466 277774
rect 276702 277538 276734 277774
rect 276114 277454 276734 277538
rect 276114 277218 276146 277454
rect 276382 277218 276466 277454
rect 276702 277218 276734 277454
rect 276114 241774 276734 277218
rect 276114 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 276734 241774
rect 276114 241454 276734 241538
rect 276114 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 276734 241454
rect 276114 205774 276734 241218
rect 276114 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 276734 205774
rect 276114 205454 276734 205538
rect 276114 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 276734 205454
rect 276114 169774 276734 205218
rect 276114 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 276734 169774
rect 276114 169454 276734 169538
rect 276114 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 276734 169454
rect 276114 133774 276734 169218
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 276114 97774 276734 133218
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 276114 61774 276734 97218
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 281494 280454 316938
rect 279834 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 280454 281494
rect 279834 281174 280454 281258
rect 279834 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 280454 281174
rect 279834 245494 280454 280938
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 279834 209494 280454 244938
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 279834 173494 280454 208938
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 279834 137494 280454 172938
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 279834 101494 280454 136938
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 279834 65494 280454 100938
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 281398 31789 281458 360163
rect 282686 289101 282746 369139
rect 283054 360210 283114 369411
rect 283790 362269 283850 369547
rect 283971 369476 284037 369477
rect 283971 369412 283972 369476
rect 284036 369412 284037 369476
rect 283971 369411 284037 369412
rect 284891 369476 284957 369477
rect 284891 369412 284892 369476
rect 284956 369412 284957 369476
rect 284891 369411 284957 369412
rect 283787 362268 283853 362269
rect 283787 362204 283788 362268
rect 283852 362204 283853 362268
rect 283787 362203 283853 362204
rect 283974 360229 284034 369411
rect 284894 367573 284954 369411
rect 285630 367845 285690 371859
rect 288019 369884 288085 369885
rect 288019 369820 288020 369884
rect 288084 369820 288085 369884
rect 288019 369819 288085 369820
rect 287283 369476 287349 369477
rect 287283 369412 287284 369476
rect 287348 369412 287349 369476
rect 287283 369411 287349 369412
rect 285627 367844 285693 367845
rect 285627 367780 285628 367844
rect 285692 367780 285693 367844
rect 285627 367779 285693 367780
rect 284891 367572 284957 367573
rect 284891 367508 284892 367572
rect 284956 367508 284957 367572
rect 284891 367507 284957 367508
rect 282870 360150 283114 360210
rect 283971 360228 284037 360229
rect 283971 360164 283972 360228
rect 284036 360164 284037 360228
rect 283971 360163 284037 360164
rect 282870 321570 282930 360150
rect 283971 321876 284037 321877
rect 283971 321812 283972 321876
rect 284036 321812 284037 321876
rect 283971 321811 284037 321812
rect 282870 321510 283114 321570
rect 283054 319293 283114 321510
rect 283419 320380 283485 320381
rect 283419 320316 283420 320380
rect 283484 320316 283485 320380
rect 283419 320315 283485 320316
rect 283787 320380 283853 320381
rect 283787 320316 283788 320380
rect 283852 320316 283853 320380
rect 283787 320315 283853 320316
rect 283235 320108 283301 320109
rect 283235 320044 283236 320108
rect 283300 320044 283301 320108
rect 283422 320106 283482 320315
rect 283422 320046 283666 320106
rect 283235 320043 283301 320044
rect 283051 319292 283117 319293
rect 283051 319228 283052 319292
rect 283116 319228 283117 319292
rect 283051 319227 283117 319228
rect 282867 318612 282933 318613
rect 282867 318548 282868 318612
rect 282932 318548 282933 318612
rect 282867 318547 282933 318548
rect 282870 318205 282930 318547
rect 282867 318204 282933 318205
rect 282867 318140 282868 318204
rect 282932 318140 282933 318204
rect 282867 318139 282933 318140
rect 283238 311910 283298 320043
rect 283419 319972 283485 319973
rect 283419 319908 283420 319972
rect 283484 319908 283485 319972
rect 283419 319907 283485 319908
rect 282870 311850 283298 311910
rect 282683 289100 282749 289101
rect 282683 289036 282684 289100
rect 282748 289036 282749 289100
rect 282683 289035 282749 289036
rect 282870 220557 282930 311850
rect 282867 220556 282933 220557
rect 282867 220492 282868 220556
rect 282932 220492 282933 220556
rect 282867 220491 282933 220492
rect 283422 220285 283482 319907
rect 283606 318341 283666 320046
rect 283603 318340 283669 318341
rect 283603 318276 283604 318340
rect 283668 318276 283669 318340
rect 283603 318275 283669 318276
rect 283790 317933 283850 320315
rect 283974 319293 284034 321811
rect 284339 320108 284405 320109
rect 284339 320044 284340 320108
rect 284404 320044 284405 320108
rect 284339 320043 284405 320044
rect 283971 319292 284037 319293
rect 283971 319228 283972 319292
rect 284036 319228 284037 319292
rect 283971 319227 284037 319228
rect 283787 317932 283853 317933
rect 283787 317868 283788 317932
rect 283852 317868 283853 317932
rect 283787 317867 283853 317868
rect 283419 220284 283485 220285
rect 283419 220220 283420 220284
rect 283484 220220 283485 220284
rect 283419 220219 283485 220220
rect 284342 219333 284402 320043
rect 284523 317660 284589 317661
rect 284523 317596 284524 317660
rect 284588 317596 284589 317660
rect 284523 317595 284589 317596
rect 284526 307189 284586 317595
rect 284523 307188 284589 307189
rect 284523 307124 284524 307188
rect 284588 307124 284589 307188
rect 284523 307123 284589 307124
rect 284894 283525 284954 367507
rect 287286 320789 287346 369411
rect 288022 367709 288082 369819
rect 288019 367708 288085 367709
rect 288019 367644 288020 367708
rect 288084 367644 288085 367708
rect 288019 367643 288085 367644
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 288019 321604 288085 321605
rect 288019 321540 288020 321604
rect 288084 321540 288085 321604
rect 288019 321539 288085 321540
rect 288022 320789 288082 321539
rect 287283 320788 287349 320789
rect 287283 320724 287284 320788
rect 287348 320724 287349 320788
rect 287283 320723 287349 320724
rect 288019 320788 288085 320789
rect 288019 320724 288020 320788
rect 288084 320724 288085 320788
rect 288019 320723 288085 320724
rect 288939 320380 289005 320381
rect 288939 320316 288940 320380
rect 289004 320316 289005 320380
rect 288939 320315 289005 320316
rect 285627 320244 285693 320245
rect 285627 320180 285628 320244
rect 285692 320180 285693 320244
rect 285627 320179 285693 320180
rect 287835 320244 287901 320245
rect 287835 320180 287836 320244
rect 287900 320180 287901 320244
rect 287835 320179 287901 320180
rect 288755 320244 288821 320245
rect 288755 320180 288756 320244
rect 288820 320180 288821 320244
rect 288755 320179 288821 320180
rect 285443 319972 285509 319973
rect 285443 319908 285444 319972
rect 285508 319908 285509 319972
rect 285443 319907 285509 319908
rect 285446 319293 285506 319907
rect 285443 319292 285509 319293
rect 285443 319228 285444 319292
rect 285508 319228 285509 319292
rect 285443 319227 285509 319228
rect 285630 317933 285690 320179
rect 285811 320108 285877 320109
rect 285811 320044 285812 320108
rect 285876 320044 285877 320108
rect 285811 320043 285877 320044
rect 286731 320108 286797 320109
rect 286731 320044 286732 320108
rect 286796 320044 286797 320108
rect 286731 320043 286797 320044
rect 287651 320108 287717 320109
rect 287651 320044 287652 320108
rect 287716 320044 287717 320108
rect 287651 320043 287717 320044
rect 285627 317932 285693 317933
rect 285627 317868 285628 317932
rect 285692 317868 285693 317932
rect 285627 317867 285693 317868
rect 285627 317524 285693 317525
rect 285627 317460 285628 317524
rect 285692 317460 285693 317524
rect 285627 317459 285693 317460
rect 284891 283524 284957 283525
rect 284891 283460 284892 283524
rect 284956 283460 284957 283524
rect 284891 283459 284957 283460
rect 285630 220693 285690 317459
rect 285814 314533 285874 320043
rect 286734 318749 286794 320043
rect 287654 319293 287714 320043
rect 287651 319292 287717 319293
rect 287651 319228 287652 319292
rect 287716 319228 287717 319292
rect 287651 319227 287717 319228
rect 286731 318748 286797 318749
rect 286731 318684 286732 318748
rect 286796 318684 286797 318748
rect 286731 318683 286797 318684
rect 287099 318748 287165 318749
rect 287099 318684 287100 318748
rect 287164 318684 287165 318748
rect 287099 318683 287165 318684
rect 285995 317660 286061 317661
rect 285995 317596 285996 317660
rect 286060 317596 286061 317660
rect 285995 317595 286061 317596
rect 285811 314532 285877 314533
rect 285811 314468 285812 314532
rect 285876 314468 285877 314532
rect 285811 314467 285877 314468
rect 285998 309909 286058 317595
rect 285995 309908 286061 309909
rect 285995 309844 285996 309908
rect 286060 309844 286061 309908
rect 285995 309843 286061 309844
rect 285627 220692 285693 220693
rect 285627 220628 285628 220692
rect 285692 220628 285693 220692
rect 285627 220627 285693 220628
rect 287102 220285 287162 318683
rect 287283 317524 287349 317525
rect 287283 317460 287284 317524
rect 287348 317460 287349 317524
rect 287283 317459 287349 317460
rect 287467 317524 287533 317525
rect 287467 317460 287468 317524
rect 287532 317460 287533 317524
rect 287467 317459 287533 317460
rect 287286 304333 287346 317459
rect 287470 309365 287530 317459
rect 287467 309364 287533 309365
rect 287467 309300 287468 309364
rect 287532 309300 287533 309364
rect 287467 309299 287533 309300
rect 287283 304332 287349 304333
rect 287283 304268 287284 304332
rect 287348 304268 287349 304332
rect 287283 304267 287349 304268
rect 287838 223549 287898 320179
rect 288019 320108 288085 320109
rect 288019 320044 288020 320108
rect 288084 320044 288085 320108
rect 288019 320043 288085 320044
rect 288203 320108 288269 320109
rect 288203 320044 288204 320108
rect 288268 320044 288269 320108
rect 288203 320043 288269 320044
rect 288571 320108 288637 320109
rect 288571 320044 288572 320108
rect 288636 320044 288637 320108
rect 288571 320043 288637 320044
rect 288022 318749 288082 320043
rect 288206 318749 288266 320043
rect 288019 318748 288085 318749
rect 288019 318684 288020 318748
rect 288084 318684 288085 318748
rect 288019 318683 288085 318684
rect 288203 318748 288269 318749
rect 288203 318684 288204 318748
rect 288268 318684 288269 318748
rect 288203 318683 288269 318684
rect 288387 317524 288453 317525
rect 288387 317460 288388 317524
rect 288452 317460 288453 317524
rect 288387 317459 288453 317460
rect 287835 223548 287901 223549
rect 287835 223484 287836 223548
rect 287900 223484 287901 223548
rect 287835 223483 287901 223484
rect 287099 220284 287165 220285
rect 287099 220220 287100 220284
rect 287164 220220 287165 220284
rect 287099 220219 287165 220220
rect 284339 219332 284405 219333
rect 284339 219268 284340 219332
rect 284404 219268 284405 219332
rect 284339 219267 284405 219268
rect 288390 219197 288450 317459
rect 288574 312085 288634 320043
rect 288758 318749 288818 320179
rect 288755 318748 288821 318749
rect 288755 318684 288756 318748
rect 288820 318684 288821 318748
rect 288755 318683 288821 318684
rect 288571 312084 288637 312085
rect 288571 312020 288572 312084
rect 288636 312020 288637 312084
rect 288571 312019 288637 312020
rect 288942 310453 289002 320315
rect 289491 320244 289557 320245
rect 289491 320180 289492 320244
rect 289556 320180 289557 320244
rect 289491 320179 289557 320180
rect 289123 320108 289189 320109
rect 289123 320044 289124 320108
rect 289188 320044 289189 320108
rect 289123 320043 289189 320044
rect 289126 314397 289186 320043
rect 289307 319972 289373 319973
rect 289307 319908 289308 319972
rect 289372 319908 289373 319972
rect 289307 319907 289373 319908
rect 289310 319293 289370 319907
rect 289307 319292 289373 319293
rect 289307 319228 289308 319292
rect 289372 319228 289373 319292
rect 289307 319227 289373 319228
rect 289494 318749 289554 320179
rect 289491 318748 289557 318749
rect 289491 318684 289492 318748
rect 289556 318684 289557 318748
rect 289491 318683 289557 318684
rect 289123 314396 289189 314397
rect 289123 314332 289124 314396
rect 289188 314332 289189 314396
rect 289123 314331 289189 314332
rect 288939 310452 289005 310453
rect 288939 310388 288940 310452
rect 289004 310388 289005 310452
rect 288939 310387 289005 310388
rect 289794 291454 290414 326898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 296483 371380 296549 371381
rect 296483 371316 296484 371380
rect 296548 371316 296549 371380
rect 296483 371315 296549 371316
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293171 321740 293237 321741
rect 293171 321676 293172 321740
rect 293236 321676 293237 321740
rect 293171 321675 293237 321676
rect 291883 320788 291949 320789
rect 291883 320724 291884 320788
rect 291948 320724 291949 320788
rect 291883 320723 291949 320724
rect 292619 320788 292685 320789
rect 292619 320724 292620 320788
rect 292684 320724 292685 320788
rect 292619 320723 292685 320724
rect 290779 320380 290845 320381
rect 290779 320316 290780 320380
rect 290844 320316 290845 320380
rect 290779 320315 290845 320316
rect 290595 320108 290661 320109
rect 290595 320044 290596 320108
rect 290660 320044 290661 320108
rect 290595 320043 290661 320044
rect 290598 319293 290658 320043
rect 290595 319292 290661 319293
rect 290595 319228 290596 319292
rect 290660 319228 290661 319292
rect 290595 319227 290661 319228
rect 290782 311910 290842 320315
rect 290963 320244 291029 320245
rect 290963 320180 290964 320244
rect 291028 320180 291029 320244
rect 290963 320179 291029 320180
rect 291331 320244 291397 320245
rect 291331 320180 291332 320244
rect 291396 320180 291397 320244
rect 291331 320179 291397 320180
rect 290966 319293 291026 320179
rect 291147 319972 291213 319973
rect 291147 319908 291148 319972
rect 291212 319908 291213 319972
rect 291147 319907 291213 319908
rect 290963 319292 291029 319293
rect 290963 319228 290964 319292
rect 291028 319228 291029 319292
rect 290963 319227 291029 319228
rect 291150 318749 291210 319907
rect 291147 318748 291213 318749
rect 291147 318684 291148 318748
rect 291212 318684 291213 318748
rect 291147 318683 291213 318684
rect 291147 318204 291213 318205
rect 291147 318140 291148 318204
rect 291212 318140 291213 318204
rect 291147 318139 291213 318140
rect 290598 311850 290842 311910
rect 290598 309773 290658 311850
rect 290595 309772 290661 309773
rect 290595 309708 290596 309772
rect 290660 309708 290661 309772
rect 290595 309707 290661 309708
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 291150 219877 291210 318139
rect 291334 317661 291394 320179
rect 291515 320108 291581 320109
rect 291515 320044 291516 320108
rect 291580 320044 291581 320108
rect 291515 320043 291581 320044
rect 291699 320108 291765 320109
rect 291699 320044 291700 320108
rect 291764 320044 291765 320108
rect 291699 320043 291765 320044
rect 291518 319293 291578 320043
rect 291515 319292 291581 319293
rect 291515 319228 291516 319292
rect 291580 319228 291581 319292
rect 291515 319227 291581 319228
rect 291702 318069 291762 320043
rect 291699 318068 291765 318069
rect 291699 318004 291700 318068
rect 291764 318004 291765 318068
rect 291699 318003 291765 318004
rect 291886 317933 291946 320723
rect 292067 320108 292133 320109
rect 292067 320044 292068 320108
rect 292132 320044 292133 320108
rect 292067 320043 292133 320044
rect 292070 318885 292130 320043
rect 292435 319972 292501 319973
rect 292435 319908 292436 319972
rect 292500 319908 292501 319972
rect 292435 319907 292501 319908
rect 292067 318884 292133 318885
rect 292067 318820 292068 318884
rect 292132 318820 292133 318884
rect 292067 318819 292133 318820
rect 292438 318205 292498 319907
rect 292622 318477 292682 320723
rect 292803 320380 292869 320381
rect 292803 320316 292804 320380
rect 292868 320316 292869 320380
rect 292803 320315 292869 320316
rect 292619 318476 292685 318477
rect 292619 318412 292620 318476
rect 292684 318412 292685 318476
rect 292619 318411 292685 318412
rect 292806 318341 292866 320315
rect 292987 320108 293053 320109
rect 292987 320044 292988 320108
rect 293052 320044 293053 320108
rect 292987 320043 293053 320044
rect 292803 318340 292869 318341
rect 292803 318276 292804 318340
rect 292868 318276 292869 318340
rect 292803 318275 292869 318276
rect 292435 318204 292501 318205
rect 292435 318140 292436 318204
rect 292500 318140 292501 318204
rect 292435 318139 292501 318140
rect 291883 317932 291949 317933
rect 291883 317868 291884 317932
rect 291948 317868 291949 317932
rect 291883 317867 291949 317868
rect 291331 317660 291397 317661
rect 291331 317596 291332 317660
rect 291396 317596 291397 317660
rect 291331 317595 291397 317596
rect 291331 317524 291397 317525
rect 291331 317460 291332 317524
rect 291396 317460 291397 317524
rect 291331 317459 291397 317460
rect 291515 317524 291581 317525
rect 291515 317460 291516 317524
rect 291580 317460 291581 317524
rect 291515 317459 291581 317460
rect 292619 317524 292685 317525
rect 292619 317460 292620 317524
rect 292684 317460 292685 317524
rect 292619 317459 292685 317460
rect 291334 297397 291394 317459
rect 291518 309637 291578 317459
rect 291515 309636 291581 309637
rect 291515 309572 291516 309636
rect 291580 309572 291581 309636
rect 291515 309571 291581 309572
rect 291331 297396 291397 297397
rect 291331 297332 291332 297396
rect 291396 297332 291397 297396
rect 291331 297331 291397 297332
rect 292622 221917 292682 317459
rect 292990 312085 293050 320043
rect 293174 319429 293234 321675
rect 293355 320244 293421 320245
rect 293355 320180 293356 320244
rect 293420 320180 293421 320244
rect 293355 320179 293421 320180
rect 293171 319428 293237 319429
rect 293171 319364 293172 319428
rect 293236 319364 293237 319428
rect 293171 319363 293237 319364
rect 293358 318885 293418 320179
rect 293355 318884 293421 318885
rect 293355 318820 293356 318884
rect 293420 318820 293421 318884
rect 293355 318819 293421 318820
rect 292987 312084 293053 312085
rect 292987 312020 292988 312084
rect 293052 312020 293053 312084
rect 292987 312019 293053 312020
rect 293514 295174 294134 330618
rect 294459 320788 294525 320789
rect 294459 320724 294460 320788
rect 294524 320724 294525 320788
rect 294459 320723 294525 320724
rect 295747 320788 295813 320789
rect 295747 320724 295748 320788
rect 295812 320724 295813 320788
rect 295747 320723 295813 320724
rect 294275 320108 294341 320109
rect 294275 320044 294276 320108
rect 294340 320044 294341 320108
rect 294275 320043 294341 320044
rect 294278 315349 294338 320043
rect 294462 318885 294522 320723
rect 294643 320244 294709 320245
rect 294643 320180 294644 320244
rect 294708 320180 294709 320244
rect 294643 320179 294709 320180
rect 294827 320244 294893 320245
rect 294827 320180 294828 320244
rect 294892 320180 294893 320244
rect 294827 320179 294893 320180
rect 294459 318884 294525 318885
rect 294459 318820 294460 318884
rect 294524 318820 294525 318884
rect 294459 318819 294525 318820
rect 294459 317660 294525 317661
rect 294459 317596 294460 317660
rect 294524 317596 294525 317660
rect 294459 317595 294525 317596
rect 294275 315348 294341 315349
rect 294275 315284 294276 315348
rect 294340 315284 294341 315348
rect 294275 315283 294341 315284
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 292619 221916 292685 221917
rect 292619 221852 292620 221916
rect 292684 221852 292685 221916
rect 292619 221851 292685 221852
rect 291147 219876 291213 219877
rect 291147 219812 291148 219876
rect 291212 219812 291213 219876
rect 291147 219811 291213 219812
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 288387 219196 288453 219197
rect 288387 219132 288388 219196
rect 288452 219132 288453 219196
rect 288387 219131 288453 219132
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 281395 31788 281461 31789
rect 281395 31724 281396 31788
rect 281460 31724 281461 31788
rect 281395 31723 281461 31724
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 187174 294134 222618
rect 294462 222053 294522 317595
rect 294646 224909 294706 320179
rect 294830 319429 294890 320179
rect 295011 320108 295077 320109
rect 295011 320044 295012 320108
rect 295076 320044 295077 320108
rect 295011 320043 295077 320044
rect 295563 320108 295629 320109
rect 295563 320044 295564 320108
rect 295628 320044 295629 320108
rect 295563 320043 295629 320044
rect 294827 319428 294893 319429
rect 294827 319364 294828 319428
rect 294892 319364 294893 319428
rect 294827 319363 294893 319364
rect 295014 318885 295074 320043
rect 295379 319972 295445 319973
rect 295379 319908 295380 319972
rect 295444 319908 295445 319972
rect 295379 319907 295445 319908
rect 295011 318884 295077 318885
rect 295011 318820 295012 318884
rect 295076 318820 295077 318884
rect 295011 318819 295077 318820
rect 294827 317932 294893 317933
rect 294827 317868 294828 317932
rect 294892 317868 294893 317932
rect 294827 317867 294893 317868
rect 294830 315077 294890 317867
rect 294827 315076 294893 315077
rect 294827 315012 294828 315076
rect 294892 315012 294893 315076
rect 294827 315011 294893 315012
rect 295382 314261 295442 319907
rect 295566 317525 295626 320043
rect 295563 317524 295629 317525
rect 295563 317460 295564 317524
rect 295628 317460 295629 317524
rect 295563 317459 295629 317460
rect 295379 314260 295445 314261
rect 295379 314196 295380 314260
rect 295444 314196 295445 314260
rect 295379 314195 295445 314196
rect 295750 307189 295810 320723
rect 295931 320108 295997 320109
rect 295931 320044 295932 320108
rect 295996 320044 295997 320108
rect 295931 320043 295997 320044
rect 295934 318885 295994 320043
rect 296486 319429 296546 371315
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 299979 369476 300045 369477
rect 299979 369412 299980 369476
rect 300044 369412 300045 369476
rect 299979 369411 300045 369412
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297035 320108 297101 320109
rect 297035 320044 297036 320108
rect 297100 320044 297101 320108
rect 297035 320043 297101 320044
rect 296851 319972 296917 319973
rect 296851 319908 296852 319972
rect 296916 319908 296917 319972
rect 296851 319907 296917 319908
rect 296483 319428 296549 319429
rect 296483 319364 296484 319428
rect 296548 319364 296549 319428
rect 296483 319363 296549 319364
rect 296854 318885 296914 319907
rect 295931 318884 295997 318885
rect 295931 318820 295932 318884
rect 295996 318820 295997 318884
rect 295931 318819 295997 318820
rect 296667 318884 296733 318885
rect 296667 318820 296668 318884
rect 296732 318820 296733 318884
rect 296667 318819 296733 318820
rect 296851 318884 296917 318885
rect 296851 318820 296852 318884
rect 296916 318820 296917 318884
rect 296851 318819 296917 318820
rect 295931 318612 295997 318613
rect 295931 318548 295932 318612
rect 295996 318548 295997 318612
rect 295931 318547 295997 318548
rect 295747 307188 295813 307189
rect 295747 307124 295748 307188
rect 295812 307124 295813 307188
rect 295747 307123 295813 307124
rect 295934 240685 295994 318547
rect 296670 314125 296730 318819
rect 296667 314124 296733 314125
rect 296667 314060 296668 314124
rect 296732 314060 296733 314124
rect 296667 314059 296733 314060
rect 297038 313989 297098 320043
rect 297035 313988 297101 313989
rect 297035 313924 297036 313988
rect 297100 313924 297101 313988
rect 297035 313923 297101 313924
rect 297234 298894 297854 334338
rect 299243 320788 299309 320789
rect 299243 320724 299244 320788
rect 299308 320724 299309 320788
rect 299243 320723 299309 320724
rect 297955 320244 298021 320245
rect 297955 320180 297956 320244
rect 298020 320180 298021 320244
rect 297955 320179 298021 320180
rect 299059 320244 299125 320245
rect 299059 320180 299060 320244
rect 299124 320180 299125 320244
rect 299059 320179 299125 320180
rect 297958 318477 298018 320179
rect 298323 320108 298389 320109
rect 298323 320044 298324 320108
rect 298388 320044 298389 320108
rect 298323 320043 298389 320044
rect 298139 318748 298205 318749
rect 298139 318684 298140 318748
rect 298204 318684 298205 318748
rect 298139 318683 298205 318684
rect 297955 318476 298021 318477
rect 297955 318412 297956 318476
rect 298020 318412 298021 318476
rect 297955 318411 298021 318412
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 295931 240684 295997 240685
rect 295931 240620 295932 240684
rect 295996 240620 295997 240684
rect 295931 240619 295997 240620
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 294643 224908 294709 224909
rect 294643 224844 294644 224908
rect 294708 224844 294709 224908
rect 294643 224843 294709 224844
rect 294459 222052 294525 222053
rect 294459 221988 294460 222052
rect 294524 221988 294525 222052
rect 294459 221987 294525 221988
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 190894 297854 226338
rect 298142 221781 298202 318683
rect 298326 307053 298386 320043
rect 299062 318749 299122 320179
rect 299246 318885 299306 320723
rect 299982 320653 300042 369411
rect 300954 338614 301574 374058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 630334 305294 665778
rect 304674 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 305294 630334
rect 304674 630014 305294 630098
rect 304674 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 305294 630014
rect 304674 594334 305294 629778
rect 304674 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 305294 594334
rect 304674 594014 305294 594098
rect 304674 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 305294 594014
rect 304674 558334 305294 593778
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 304674 522334 305294 557778
rect 304674 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 305294 522334
rect 304674 522014 305294 522098
rect 304674 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 305294 522014
rect 304674 486334 305294 521778
rect 304674 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 305294 486334
rect 304674 486014 305294 486098
rect 304674 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 305294 486014
rect 304674 450334 305294 485778
rect 304674 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 305294 450334
rect 304674 450014 305294 450098
rect 304674 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 305294 450014
rect 304674 414334 305294 449778
rect 304674 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 305294 414334
rect 304674 414014 305294 414098
rect 304674 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 305294 414014
rect 304674 378334 305294 413778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 598054 309014 633498
rect 308394 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 309014 598054
rect 308394 597734 309014 597818
rect 308394 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 309014 597734
rect 308394 562054 309014 597498
rect 308394 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 309014 562054
rect 308394 561734 309014 561818
rect 308394 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 309014 561734
rect 308394 526054 309014 561498
rect 308394 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 309014 526054
rect 308394 525734 309014 525818
rect 308394 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 309014 525734
rect 308394 490054 309014 525498
rect 308394 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 309014 490054
rect 308394 489734 309014 489818
rect 308394 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 309014 489734
rect 308394 454054 309014 489498
rect 308394 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 309014 454054
rect 308394 453734 309014 453818
rect 308394 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 309014 453734
rect 308394 418054 309014 453498
rect 308394 417818 308426 418054
rect 308662 417818 308746 418054
rect 308982 417818 309014 418054
rect 308394 417734 309014 417818
rect 308394 417498 308426 417734
rect 308662 417498 308746 417734
rect 308982 417498 309014 417734
rect 305499 386340 305565 386341
rect 305499 386276 305500 386340
rect 305564 386276 305565 386340
rect 305499 386275 305565 386276
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 302739 369476 302805 369477
rect 302739 369412 302740 369476
rect 302804 369412 302805 369476
rect 302739 369411 302805 369412
rect 303659 369476 303725 369477
rect 303659 369412 303660 369476
rect 303724 369412 303725 369476
rect 303659 369411 303725 369412
rect 302742 345030 302802 369411
rect 302742 344970 302986 345030
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 299979 320652 300045 320653
rect 299979 320588 299980 320652
rect 300044 320588 300045 320652
rect 299979 320587 300045 320588
rect 299611 320380 299677 320381
rect 299611 320316 299612 320380
rect 299676 320316 299677 320380
rect 299611 320315 299677 320316
rect 299795 320380 299861 320381
rect 299795 320316 299796 320380
rect 299860 320316 299861 320380
rect 299795 320315 299861 320316
rect 299427 320108 299493 320109
rect 299427 320044 299428 320108
rect 299492 320044 299493 320108
rect 299427 320043 299493 320044
rect 299243 318884 299309 318885
rect 299243 318820 299244 318884
rect 299308 318820 299309 318884
rect 299243 318819 299309 318820
rect 299059 318748 299125 318749
rect 299059 318684 299060 318748
rect 299124 318684 299125 318748
rect 299059 318683 299125 318684
rect 298507 317932 298573 317933
rect 298507 317868 298508 317932
rect 298572 317868 298573 317932
rect 298507 317867 298573 317868
rect 298510 312493 298570 317867
rect 299430 315893 299490 320043
rect 299614 318746 299674 320315
rect 299798 318885 299858 320315
rect 300531 320244 300597 320245
rect 300531 320180 300532 320244
rect 300596 320180 300597 320244
rect 300531 320179 300597 320180
rect 299979 320108 300045 320109
rect 299979 320044 299980 320108
rect 300044 320044 300045 320108
rect 299979 320043 300045 320044
rect 299982 319429 300042 320043
rect 299979 319428 300045 319429
rect 299979 319364 299980 319428
rect 300044 319364 300045 319428
rect 299979 319363 300045 319364
rect 300534 318885 300594 320179
rect 300715 320108 300781 320109
rect 300715 320044 300716 320108
rect 300780 320044 300781 320108
rect 300715 320043 300781 320044
rect 300718 319429 300778 320043
rect 300715 319428 300781 319429
rect 300715 319364 300716 319428
rect 300780 319364 300781 319428
rect 300715 319363 300781 319364
rect 299795 318884 299861 318885
rect 299795 318820 299796 318884
rect 299860 318820 299861 318884
rect 299795 318819 299861 318820
rect 300531 318884 300597 318885
rect 300531 318820 300532 318884
rect 300596 318820 300597 318884
rect 300531 318819 300597 318820
rect 299614 318686 299858 318746
rect 299611 317524 299677 317525
rect 299611 317460 299612 317524
rect 299676 317460 299677 317524
rect 299611 317459 299677 317460
rect 299427 315892 299493 315893
rect 299427 315828 299428 315892
rect 299492 315828 299493 315892
rect 299427 315827 299493 315828
rect 299614 315213 299674 317459
rect 299611 315212 299677 315213
rect 299611 315148 299612 315212
rect 299676 315148 299677 315212
rect 299611 315147 299677 315148
rect 298507 312492 298573 312493
rect 298507 312428 298508 312492
rect 298572 312428 298573 312492
rect 298507 312427 298573 312428
rect 298323 307052 298389 307053
rect 298323 306988 298324 307052
rect 298388 306988 298389 307052
rect 298323 306987 298389 306988
rect 299798 231301 299858 318686
rect 299979 318340 300045 318341
rect 299979 318276 299980 318340
rect 300044 318276 300045 318340
rect 299979 318275 300045 318276
rect 299982 232661 300042 318275
rect 300954 302614 301574 338058
rect 301819 320108 301885 320109
rect 301819 320044 301820 320108
rect 301884 320044 301885 320108
rect 301819 320043 301885 320044
rect 302371 320108 302437 320109
rect 302371 320044 302372 320108
rect 302436 320044 302437 320108
rect 302371 320043 302437 320044
rect 301822 319429 301882 320043
rect 301819 319428 301885 319429
rect 301819 319364 301820 319428
rect 301884 319364 301885 319428
rect 301819 319363 301885 319364
rect 302003 318748 302069 318749
rect 302003 318684 302004 318748
rect 302068 318684 302069 318748
rect 302003 318683 302069 318684
rect 301819 317524 301885 317525
rect 301819 317460 301820 317524
rect 301884 317460 301885 317524
rect 301819 317459 301885 317460
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 299979 232660 300045 232661
rect 299979 232596 299980 232660
rect 300044 232596 300045 232660
rect 299979 232595 300045 232596
rect 299795 231300 299861 231301
rect 299795 231236 299796 231300
rect 299860 231236 299861 231300
rect 299795 231235 299861 231236
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 298139 221780 298205 221781
rect 298139 221716 298140 221780
rect 298204 221716 298205 221780
rect 298139 221715 298205 221716
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 194614 301574 230058
rect 301822 222189 301882 317459
rect 302006 227629 302066 318683
rect 302374 311910 302434 320043
rect 302926 319429 302986 344970
rect 303662 321061 303722 369411
rect 304674 342334 305294 377778
rect 305502 369477 305562 386275
rect 308394 382054 309014 417498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 312114 601774 312734 637218
rect 312114 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 312734 601774
rect 312114 601454 312734 601538
rect 312114 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 312734 601454
rect 312114 565774 312734 601218
rect 312114 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 312734 565774
rect 312114 565454 312734 565538
rect 312114 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 312734 565454
rect 312114 529774 312734 565218
rect 312114 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 312734 529774
rect 312114 529454 312734 529538
rect 312114 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 312734 529454
rect 312114 493774 312734 529218
rect 312114 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 312734 493774
rect 312114 493454 312734 493538
rect 312114 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 312734 493454
rect 312114 457774 312734 493218
rect 312114 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 312734 457774
rect 312114 457454 312734 457538
rect 312114 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 312734 457454
rect 312114 421774 312734 457218
rect 312114 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 312734 421774
rect 312114 421454 312734 421538
rect 312114 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 312734 421454
rect 309179 403612 309245 403613
rect 309179 403548 309180 403612
rect 309244 403548 309245 403612
rect 309179 403547 309245 403548
rect 308394 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 309014 382054
rect 308394 381734 309014 381818
rect 308394 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 309014 381734
rect 306419 377364 306485 377365
rect 306419 377300 306420 377364
rect 306484 377300 306485 377364
rect 306419 377299 306485 377300
rect 306422 369477 306482 377299
rect 307707 374644 307773 374645
rect 307707 374580 307708 374644
rect 307772 374580 307773 374644
rect 307707 374579 307773 374580
rect 307523 372604 307589 372605
rect 307523 372540 307524 372604
rect 307588 372540 307589 372604
rect 307523 372539 307589 372540
rect 305499 369476 305565 369477
rect 305499 369412 305500 369476
rect 305564 369412 305565 369476
rect 305499 369411 305565 369412
rect 306419 369476 306485 369477
rect 306419 369412 306420 369476
rect 306484 369412 306485 369476
rect 306419 369411 306485 369412
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 303659 321060 303725 321061
rect 303659 320996 303660 321060
rect 303724 320996 303725 321060
rect 303659 320995 303725 320996
rect 303659 320244 303725 320245
rect 303659 320180 303660 320244
rect 303724 320180 303725 320244
rect 303659 320179 303725 320180
rect 302923 319428 302989 319429
rect 302923 319364 302924 319428
rect 302988 319364 302989 319428
rect 302923 319363 302989 319364
rect 303475 318340 303541 318341
rect 303475 318276 303476 318340
rect 303540 318276 303541 318340
rect 303475 318275 303541 318276
rect 302739 317932 302805 317933
rect 302739 317868 302740 317932
rect 302804 317868 302805 317932
rect 302739 317867 302805 317868
rect 302190 311850 302434 311910
rect 302003 227628 302069 227629
rect 302003 227564 302004 227628
rect 302068 227564 302069 227628
rect 302003 227563 302069 227564
rect 302190 227357 302250 311850
rect 302742 241501 302802 317867
rect 302923 317796 302989 317797
rect 302923 317732 302924 317796
rect 302988 317732 302989 317796
rect 302923 317731 302989 317732
rect 302926 307733 302986 317731
rect 302923 307732 302989 307733
rect 302923 307668 302924 307732
rect 302988 307668 302989 307732
rect 302923 307667 302989 307668
rect 302739 241500 302805 241501
rect 302739 241436 302740 241500
rect 302804 241436 302805 241500
rect 302739 241435 302805 241436
rect 302187 227356 302253 227357
rect 302187 227292 302188 227356
rect 302252 227292 302253 227356
rect 302187 227291 302253 227292
rect 301819 222188 301885 222189
rect 301819 222124 301820 222188
rect 301884 222124 301885 222188
rect 301819 222123 301885 222124
rect 303478 219197 303538 318275
rect 303475 219196 303541 219197
rect 303475 219132 303476 219196
rect 303540 219132 303541 219196
rect 303475 219131 303541 219132
rect 303662 213893 303722 320179
rect 303843 320108 303909 320109
rect 303843 320044 303844 320108
rect 303908 320044 303909 320108
rect 303843 320043 303909 320044
rect 304395 320108 304461 320109
rect 304395 320044 304396 320108
rect 304460 320044 304461 320108
rect 304395 320043 304461 320044
rect 303846 318205 303906 320043
rect 304398 319429 304458 320043
rect 304395 319428 304461 319429
rect 304395 319364 304396 319428
rect 304460 319364 304461 319428
rect 304395 319363 304461 319364
rect 304395 318748 304461 318749
rect 304395 318684 304396 318748
rect 304460 318684 304461 318748
rect 304395 318683 304461 318684
rect 303843 318204 303909 318205
rect 303843 318140 303844 318204
rect 303908 318140 303909 318204
rect 303843 318139 303909 318140
rect 303843 317660 303909 317661
rect 303843 317596 303844 317660
rect 303908 317596 303909 317660
rect 303843 317595 303909 317596
rect 303846 223141 303906 317595
rect 304211 317524 304277 317525
rect 304211 317460 304212 317524
rect 304276 317460 304277 317524
rect 304211 317459 304277 317460
rect 303843 223140 303909 223141
rect 303843 223076 303844 223140
rect 303908 223076 303909 223140
rect 303843 223075 303909 223076
rect 303659 213892 303725 213893
rect 303659 213828 303660 213892
rect 303724 213828 303725 213892
rect 303659 213827 303725 213828
rect 304214 208317 304274 317459
rect 304398 233205 304458 318683
rect 304674 306334 305294 341778
rect 305502 319293 305562 369411
rect 306422 321333 306482 369411
rect 307526 369341 307586 372539
rect 307710 369870 307770 374579
rect 307710 369810 308138 369870
rect 307523 369340 307589 369341
rect 307523 369276 307524 369340
rect 307588 369276 307589 369340
rect 307523 369275 307589 369276
rect 306419 321332 306485 321333
rect 306419 321268 306420 321332
rect 306484 321268 306485 321332
rect 306419 321267 306485 321268
rect 305683 320108 305749 320109
rect 305683 320044 305684 320108
rect 305748 320044 305749 320108
rect 305683 320043 305749 320044
rect 306051 320108 306117 320109
rect 306051 320044 306052 320108
rect 306116 320044 306117 320108
rect 306051 320043 306117 320044
rect 306235 320108 306301 320109
rect 306235 320044 306236 320108
rect 306300 320044 306301 320108
rect 306235 320043 306301 320044
rect 306603 320108 306669 320109
rect 306603 320044 306604 320108
rect 306668 320044 306669 320108
rect 306603 320043 306669 320044
rect 307155 320108 307221 320109
rect 307155 320044 307156 320108
rect 307220 320044 307221 320108
rect 307155 320043 307221 320044
rect 307339 320108 307405 320109
rect 307339 320044 307340 320108
rect 307404 320044 307405 320108
rect 307339 320043 307405 320044
rect 305499 319292 305565 319293
rect 305499 319228 305500 319292
rect 305564 319228 305565 319292
rect 305499 319227 305565 319228
rect 305686 318885 305746 320043
rect 306054 319429 306114 320043
rect 306238 319429 306298 320043
rect 306606 319429 306666 320043
rect 306971 319972 307037 319973
rect 306971 319908 306972 319972
rect 307036 319908 307037 319972
rect 306971 319907 307037 319908
rect 306974 319565 307034 319907
rect 306971 319564 307037 319565
rect 306971 319500 306972 319564
rect 307036 319500 307037 319564
rect 306971 319499 307037 319500
rect 306051 319428 306117 319429
rect 306051 319364 306052 319428
rect 306116 319364 306117 319428
rect 306051 319363 306117 319364
rect 306235 319428 306301 319429
rect 306235 319364 306236 319428
rect 306300 319364 306301 319428
rect 306235 319363 306301 319364
rect 306603 319428 306669 319429
rect 306603 319364 306604 319428
rect 306668 319364 306669 319428
rect 306603 319363 306669 319364
rect 307158 319293 307218 320043
rect 307155 319292 307221 319293
rect 307155 319228 307156 319292
rect 307220 319228 307221 319292
rect 307155 319227 307221 319228
rect 305683 318884 305749 318885
rect 305683 318820 305684 318884
rect 305748 318820 305749 318884
rect 305683 318819 305749 318820
rect 307342 318749 307402 320043
rect 307526 319565 307586 369275
rect 307710 321197 307770 369810
rect 308078 369749 308138 369810
rect 308075 369748 308141 369749
rect 308075 369684 308076 369748
rect 308140 369684 308141 369748
rect 308075 369683 308141 369684
rect 308394 346054 309014 381498
rect 309182 369870 309242 403547
rect 312114 385774 312734 421218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 605494 316454 640938
rect 315834 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 316454 605494
rect 315834 605174 316454 605258
rect 315834 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 316454 605174
rect 315834 569494 316454 604938
rect 315834 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 316454 569494
rect 315834 569174 316454 569258
rect 315834 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 316454 569174
rect 315834 533494 316454 568938
rect 315834 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 316454 533494
rect 315834 533174 316454 533258
rect 315834 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 316454 533174
rect 315834 497494 316454 532938
rect 315834 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 316454 497494
rect 315834 497174 316454 497258
rect 315834 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 316454 497174
rect 315834 461494 316454 496938
rect 315834 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 316454 461494
rect 315834 461174 316454 461258
rect 315834 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 316454 461174
rect 315834 425494 316454 460938
rect 315834 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 316454 425494
rect 315834 425174 316454 425258
rect 315834 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 316454 425174
rect 313411 389876 313477 389877
rect 313411 389812 313412 389876
rect 313476 389812 313477 389876
rect 313411 389811 313477 389812
rect 312114 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 312734 385774
rect 312114 385454 312734 385538
rect 312114 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 312734 385454
rect 309363 378724 309429 378725
rect 309363 378660 309364 378724
rect 309428 378660 309429 378724
rect 309363 378659 309429 378660
rect 309366 372605 309426 378659
rect 309363 372604 309429 372605
rect 309363 372540 309364 372604
rect 309428 372540 309429 372604
rect 309363 372539 309429 372540
rect 309182 369810 309794 369870
rect 309366 369749 309426 369810
rect 309363 369748 309429 369749
rect 309363 369684 309364 369748
rect 309428 369684 309429 369748
rect 309363 369683 309429 369684
rect 308394 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 309014 346054
rect 308394 345734 309014 345818
rect 308394 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 309014 345734
rect 307707 321196 307773 321197
rect 307707 321132 307708 321196
rect 307772 321132 307773 321196
rect 307707 321131 307773 321132
rect 307707 320380 307773 320381
rect 307707 320316 307708 320380
rect 307772 320316 307773 320380
rect 307707 320315 307773 320316
rect 307710 319565 307770 320315
rect 308075 320244 308141 320245
rect 308075 320180 308076 320244
rect 308140 320180 308141 320244
rect 308075 320179 308141 320180
rect 307891 320108 307957 320109
rect 307891 320044 307892 320108
rect 307956 320044 307957 320108
rect 307891 320043 307957 320044
rect 307523 319564 307589 319565
rect 307523 319500 307524 319564
rect 307588 319500 307589 319564
rect 307523 319499 307589 319500
rect 307707 319564 307773 319565
rect 307707 319500 307708 319564
rect 307772 319500 307773 319564
rect 307707 319499 307773 319500
rect 307339 318748 307405 318749
rect 307339 318684 307340 318748
rect 307404 318684 307405 318748
rect 307339 318683 307405 318684
rect 307894 318477 307954 320043
rect 308078 319429 308138 320179
rect 308075 319428 308141 319429
rect 308075 319364 308076 319428
rect 308140 319364 308141 319428
rect 308075 319363 308141 319364
rect 307891 318476 307957 318477
rect 307891 318412 307892 318476
rect 307956 318412 307957 318476
rect 307891 318411 307957 318412
rect 306235 317932 306301 317933
rect 306235 317868 306236 317932
rect 306300 317868 306301 317932
rect 306235 317867 306301 317868
rect 306051 317796 306117 317797
rect 306051 317732 306052 317796
rect 306116 317732 306117 317796
rect 306051 317731 306117 317732
rect 305683 317660 305749 317661
rect 305683 317596 305684 317660
rect 305748 317596 305749 317660
rect 305683 317595 305749 317596
rect 305499 317524 305565 317525
rect 305499 317460 305500 317524
rect 305564 317460 305565 317524
rect 305499 317459 305565 317460
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 304674 270334 305294 305778
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 304674 234334 305294 269778
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304395 233204 304461 233205
rect 304395 233140 304396 233204
rect 304460 233140 304461 233204
rect 304395 233139 304461 233140
rect 304211 208316 304277 208317
rect 304211 208252 304212 208316
rect 304276 208252 304277 208316
rect 304211 208251 304277 208252
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 198334 305294 233778
rect 305502 222597 305562 317459
rect 305686 290597 305746 317595
rect 305683 290596 305749 290597
rect 305683 290532 305684 290596
rect 305748 290532 305749 290596
rect 305683 290531 305749 290532
rect 306054 229261 306114 317731
rect 306051 229260 306117 229261
rect 306051 229196 306052 229260
rect 306116 229196 306117 229260
rect 306051 229195 306117 229196
rect 306238 226269 306298 317867
rect 306603 317660 306669 317661
rect 306603 317596 306604 317660
rect 306668 317596 306669 317660
rect 306603 317595 306669 317596
rect 306419 317524 306485 317525
rect 306419 317460 306420 317524
rect 306484 317460 306485 317524
rect 306419 317459 306485 317460
rect 306235 226268 306301 226269
rect 306235 226204 306236 226268
rect 306300 226204 306301 226268
rect 306235 226203 306301 226204
rect 306422 223413 306482 317459
rect 306606 297533 306666 317595
rect 308394 310054 309014 345498
rect 309547 320108 309613 320109
rect 309547 320044 309548 320108
rect 309612 320044 309613 320108
rect 309547 320043 309613 320044
rect 309550 319565 309610 320043
rect 309547 319564 309613 319565
rect 309547 319500 309548 319564
rect 309612 319500 309613 319564
rect 309547 319499 309613 319500
rect 309734 319293 309794 369810
rect 311571 369748 311637 369749
rect 311571 369684 311572 369748
rect 311636 369684 311637 369748
rect 311571 369683 311637 369684
rect 309915 369476 309981 369477
rect 309915 369412 309916 369476
rect 309980 369412 309981 369476
rect 309915 369411 309981 369412
rect 311019 369476 311085 369477
rect 311019 369412 311020 369476
rect 311084 369412 311085 369476
rect 311019 369411 311085 369412
rect 309918 325710 309978 369411
rect 310099 369340 310165 369341
rect 310099 369276 310100 369340
rect 310164 369276 310165 369340
rect 310099 369275 310165 369276
rect 310102 368661 310162 369275
rect 310099 368660 310165 368661
rect 310099 368596 310100 368660
rect 310164 368596 310165 368660
rect 310099 368595 310165 368596
rect 309918 325650 310162 325710
rect 309915 320108 309981 320109
rect 309915 320044 309916 320108
rect 309980 320044 309981 320108
rect 309915 320043 309981 320044
rect 309918 319293 309978 320043
rect 310102 319429 310162 325650
rect 310651 321196 310717 321197
rect 310651 321132 310652 321196
rect 310716 321132 310717 321196
rect 310651 321131 310717 321132
rect 310283 320244 310349 320245
rect 310283 320180 310284 320244
rect 310348 320180 310349 320244
rect 310283 320179 310349 320180
rect 310099 319428 310165 319429
rect 310099 319364 310100 319428
rect 310164 319364 310165 319428
rect 310099 319363 310165 319364
rect 309731 319292 309797 319293
rect 309731 319228 309732 319292
rect 309796 319228 309797 319292
rect 309731 319227 309797 319228
rect 309915 319292 309981 319293
rect 309915 319228 309916 319292
rect 309980 319228 309981 319292
rect 309915 319227 309981 319228
rect 310286 319021 310346 320179
rect 310467 320108 310533 320109
rect 310467 320044 310468 320108
rect 310532 320044 310533 320108
rect 310467 320043 310533 320044
rect 310283 319020 310349 319021
rect 310283 318956 310284 319020
rect 310348 318956 310349 319020
rect 310283 318955 310349 318956
rect 310099 318748 310165 318749
rect 310099 318684 310100 318748
rect 310164 318684 310165 318748
rect 310099 318683 310165 318684
rect 308394 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 309014 310054
rect 308394 309734 309014 309818
rect 308394 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 309014 309734
rect 306603 297532 306669 297533
rect 306603 297468 306604 297532
rect 306668 297468 306669 297532
rect 306603 297467 306669 297468
rect 308394 274054 309014 309498
rect 308394 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 309014 274054
rect 308394 273734 309014 273818
rect 308394 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 309014 273734
rect 308394 238054 309014 273498
rect 310102 254013 310162 318683
rect 310470 314941 310530 320043
rect 310654 319973 310714 321131
rect 310835 320244 310901 320245
rect 310835 320180 310836 320244
rect 310900 320180 310901 320244
rect 310835 320179 310901 320180
rect 310651 319972 310717 319973
rect 310651 319908 310652 319972
rect 310716 319908 310717 319972
rect 310651 319907 310717 319908
rect 310838 319293 310898 320179
rect 311022 319565 311082 369411
rect 311387 320244 311453 320245
rect 311387 320180 311388 320244
rect 311452 320180 311453 320244
rect 311387 320179 311453 320180
rect 311203 320108 311269 320109
rect 311203 320044 311204 320108
rect 311268 320044 311269 320108
rect 311203 320043 311269 320044
rect 311019 319564 311085 319565
rect 311019 319500 311020 319564
rect 311084 319500 311085 319564
rect 311019 319499 311085 319500
rect 310835 319292 310901 319293
rect 310835 319228 310836 319292
rect 310900 319228 310901 319292
rect 310835 319227 310901 319228
rect 311206 319021 311266 320043
rect 311390 319293 311450 320179
rect 311574 319565 311634 369683
rect 311755 369476 311821 369477
rect 311755 369412 311756 369476
rect 311820 369412 311821 369476
rect 311755 369411 311821 369412
rect 311571 319564 311637 319565
rect 311571 319500 311572 319564
rect 311636 319500 311637 319564
rect 311571 319499 311637 319500
rect 311758 319429 311818 369411
rect 312114 349774 312734 385218
rect 313227 380220 313293 380221
rect 313227 380156 313228 380220
rect 313292 380156 313293 380220
rect 313227 380155 313293 380156
rect 313230 369477 313290 380155
rect 313227 369476 313293 369477
rect 313227 369412 313228 369476
rect 313292 369412 313293 369476
rect 313227 369411 313293 369412
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 311755 319428 311821 319429
rect 311755 319364 311756 319428
rect 311820 319364 311821 319428
rect 311755 319363 311821 319364
rect 311387 319292 311453 319293
rect 311387 319228 311388 319292
rect 311452 319228 311453 319292
rect 311387 319227 311453 319228
rect 311203 319020 311269 319021
rect 311203 318956 311204 319020
rect 311268 318956 311269 319020
rect 311203 318955 311269 318956
rect 311755 317524 311821 317525
rect 311755 317460 311756 317524
rect 311820 317460 311821 317524
rect 311755 317459 311821 317460
rect 310467 314940 310533 314941
rect 310467 314876 310468 314940
rect 310532 314876 310533 314940
rect 310467 314875 310533 314876
rect 311019 314804 311085 314805
rect 311019 314740 311020 314804
rect 311084 314740 311085 314804
rect 311019 314739 311085 314740
rect 310099 254012 310165 254013
rect 310099 253948 310100 254012
rect 310164 253948 310165 254012
rect 310099 253947 310165 253948
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 306419 223412 306485 223413
rect 306419 223348 306420 223412
rect 306484 223348 306485 223412
rect 306419 223347 306485 223348
rect 305499 222596 305565 222597
rect 305499 222532 305500 222596
rect 305564 222532 305565 222596
rect 305499 222531 305565 222532
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 90334 305294 125778
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 202054 309014 237498
rect 311022 227221 311082 314739
rect 311758 312085 311818 317459
rect 312114 313774 312734 349218
rect 312859 320652 312925 320653
rect 312859 320588 312860 320652
rect 312924 320588 312925 320652
rect 312859 320587 312925 320588
rect 312862 318885 312922 320587
rect 313230 320517 313290 369411
rect 313414 369341 313474 389811
rect 315834 389494 316454 424938
rect 315834 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 316454 389494
rect 315834 389174 316454 389258
rect 315834 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 316454 389174
rect 314699 381580 314765 381581
rect 314699 381516 314700 381580
rect 314764 381516 314765 381580
rect 314699 381515 314765 381516
rect 314702 369477 314762 381515
rect 314699 369476 314765 369477
rect 314699 369412 314700 369476
rect 314764 369412 314765 369476
rect 314699 369411 314765 369412
rect 313411 369340 313477 369341
rect 313411 369276 313412 369340
rect 313476 369276 313477 369340
rect 313411 369275 313477 369276
rect 313414 320925 313474 369275
rect 314702 321197 314762 369411
rect 315834 353494 316454 388938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 316723 385660 316789 385661
rect 316723 385596 316724 385660
rect 316788 385596 316789 385660
rect 316723 385595 316789 385596
rect 316726 369341 316786 385595
rect 320219 369476 320285 369477
rect 320219 369412 320220 369476
rect 320284 369412 320285 369476
rect 320219 369411 320285 369412
rect 322795 369476 322861 369477
rect 322795 369412 322796 369476
rect 322860 369412 322861 369476
rect 322795 369411 322861 369412
rect 316723 369340 316789 369341
rect 316723 369276 316724 369340
rect 316788 369276 316789 369340
rect 316723 369275 316789 369276
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 314699 321196 314765 321197
rect 314699 321132 314700 321196
rect 314764 321132 314765 321196
rect 314699 321131 314765 321132
rect 313411 320924 313477 320925
rect 313411 320860 313412 320924
rect 313476 320860 313477 320924
rect 313411 320859 313477 320860
rect 313411 320652 313477 320653
rect 313411 320588 313412 320652
rect 313476 320588 313477 320652
rect 313411 320587 313477 320588
rect 313227 320516 313293 320517
rect 313227 320452 313228 320516
rect 313292 320452 313293 320516
rect 313227 320451 313293 320452
rect 313227 320380 313293 320381
rect 313227 320316 313228 320380
rect 313292 320316 313293 320380
rect 313227 320315 313293 320316
rect 313230 319021 313290 320315
rect 313414 319565 313474 320587
rect 314331 320244 314397 320245
rect 314331 320180 314332 320244
rect 314396 320180 314397 320244
rect 314331 320179 314397 320180
rect 314515 320244 314581 320245
rect 314515 320180 314516 320244
rect 314580 320180 314581 320244
rect 314515 320179 314581 320180
rect 314334 319701 314394 320179
rect 314331 319700 314397 319701
rect 314331 319636 314332 319700
rect 314396 319636 314397 319700
rect 314331 319635 314397 319636
rect 313411 319564 313477 319565
rect 313411 319500 313412 319564
rect 313476 319500 313477 319564
rect 313411 319499 313477 319500
rect 313227 319020 313293 319021
rect 313227 318956 313228 319020
rect 313292 318956 313293 319020
rect 313227 318955 313293 318956
rect 312859 318884 312925 318885
rect 312859 318820 312860 318884
rect 312924 318820 312925 318884
rect 312859 318819 312925 318820
rect 314518 318749 314578 320179
rect 314515 318748 314581 318749
rect 314515 318684 314516 318748
rect 314580 318684 314581 318748
rect 314515 318683 314581 318684
rect 314147 317796 314213 317797
rect 314147 317732 314148 317796
rect 314212 317732 314213 317796
rect 314147 317731 314213 317732
rect 313779 317524 313845 317525
rect 313779 317460 313780 317524
rect 313844 317460 313845 317524
rect 313779 317459 313845 317460
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 311755 312084 311821 312085
rect 311755 312020 311756 312084
rect 311820 312020 311821 312084
rect 311755 312019 311821 312020
rect 312114 277774 312734 313218
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 312114 241774 312734 277218
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 311019 227220 311085 227221
rect 311019 227156 311020 227220
rect 311084 227156 311085 227220
rect 311019 227155 311085 227156
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 308394 166054 309014 201498
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 308394 94054 309014 129498
rect 308394 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 309014 94054
rect 308394 93734 309014 93818
rect 308394 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 309014 93734
rect 308394 58054 309014 93498
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 205774 312734 241218
rect 313782 223005 313842 317459
rect 314150 315077 314210 317731
rect 315834 317494 316454 352938
rect 316539 320244 316605 320245
rect 316539 320180 316540 320244
rect 316604 320180 316605 320244
rect 316539 320179 316605 320180
rect 316542 319021 316602 320179
rect 316726 319429 316786 369275
rect 319299 321604 319365 321605
rect 319299 321540 319300 321604
rect 319364 321540 319365 321604
rect 319299 321539 319365 321540
rect 317459 321332 317525 321333
rect 317459 321268 317460 321332
rect 317524 321268 317525 321332
rect 317459 321267 317525 321268
rect 317462 320517 317522 321267
rect 317459 320516 317525 320517
rect 317459 320452 317460 320516
rect 317524 320452 317525 320516
rect 317459 320451 317525 320452
rect 318563 320516 318629 320517
rect 318563 320452 318564 320516
rect 318628 320452 318629 320516
rect 318563 320451 318629 320452
rect 319115 320516 319181 320517
rect 319115 320452 319116 320516
rect 319180 320452 319181 320516
rect 319115 320451 319181 320452
rect 317091 320380 317157 320381
rect 317091 320316 317092 320380
rect 317156 320316 317157 320380
rect 317091 320315 317157 320316
rect 316907 320108 316973 320109
rect 316907 320044 316908 320108
rect 316972 320044 316973 320108
rect 316907 320043 316973 320044
rect 316910 319565 316970 320043
rect 316907 319564 316973 319565
rect 316907 319500 316908 319564
rect 316972 319500 316973 319564
rect 316907 319499 316973 319500
rect 316723 319428 316789 319429
rect 316723 319364 316724 319428
rect 316788 319364 316789 319428
rect 316723 319363 316789 319364
rect 316539 319020 316605 319021
rect 316539 318956 316540 319020
rect 316604 318956 316605 319020
rect 316539 318955 316605 318956
rect 317094 318613 317154 320315
rect 318379 320108 318445 320109
rect 318379 320044 318380 320108
rect 318444 320044 318445 320108
rect 318379 320043 318445 320044
rect 318382 319429 318442 320043
rect 318379 319428 318445 319429
rect 318379 319364 318380 319428
rect 318444 319364 318445 319428
rect 318379 319363 318445 319364
rect 317091 318612 317157 318613
rect 317091 318548 317092 318612
rect 317156 318548 317157 318612
rect 317091 318547 317157 318548
rect 318011 317796 318077 317797
rect 318011 317732 318012 317796
rect 318076 317732 318077 317796
rect 318011 317731 318077 317732
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 317459 317524 317525 317525
rect 317459 317460 317460 317524
rect 317524 317460 317525 317524
rect 317459 317459 317525 317460
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 314147 315076 314213 315077
rect 314147 315012 314148 315076
rect 314212 315012 314213 315076
rect 314147 315011 314213 315012
rect 315834 281494 316454 316938
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 315834 245494 316454 280938
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 313779 223004 313845 223005
rect 313779 222940 313780 223004
rect 313844 222940 313845 223004
rect 313779 222939 313845 222940
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 312114 97774 312734 133218
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 209494 316454 244938
rect 317462 219061 317522 317459
rect 318014 286517 318074 317731
rect 318566 304061 318626 320451
rect 318747 320380 318813 320381
rect 318747 320316 318748 320380
rect 318812 320316 318813 320380
rect 318747 320315 318813 320316
rect 318750 317797 318810 320315
rect 319118 319021 319178 320451
rect 319302 320245 319362 321539
rect 319299 320244 319365 320245
rect 319299 320180 319300 320244
rect 319364 320180 319365 320244
rect 319299 320179 319365 320180
rect 319667 320244 319733 320245
rect 319667 320180 319668 320244
rect 319732 320180 319733 320244
rect 319667 320179 319733 320180
rect 319670 319429 319730 320179
rect 319667 319428 319733 319429
rect 319667 319364 319668 319428
rect 319732 319364 319733 319428
rect 319667 319363 319733 319364
rect 320222 319293 320282 369411
rect 322243 320788 322309 320789
rect 322243 320724 322244 320788
rect 322308 320724 322309 320788
rect 322243 320723 322309 320724
rect 321691 320244 321757 320245
rect 321691 320180 321692 320244
rect 321756 320180 321757 320244
rect 321691 320179 321757 320180
rect 322059 320244 322125 320245
rect 322059 320180 322060 320244
rect 322124 320180 322125 320244
rect 322059 320179 322125 320180
rect 320219 319292 320285 319293
rect 320219 319228 320220 319292
rect 320284 319228 320285 319292
rect 320219 319227 320285 319228
rect 319115 319020 319181 319021
rect 319115 318956 319116 319020
rect 319180 318956 319181 319020
rect 319115 318955 319181 318956
rect 321694 318885 321754 320179
rect 321691 318884 321757 318885
rect 321691 318820 321692 318884
rect 321756 318820 321757 318884
rect 321691 318819 321757 318820
rect 319299 317932 319365 317933
rect 319299 317868 319300 317932
rect 319364 317868 319365 317932
rect 319299 317867 319365 317868
rect 318747 317796 318813 317797
rect 318747 317732 318748 317796
rect 318812 317732 318813 317796
rect 318747 317731 318813 317732
rect 318563 304060 318629 304061
rect 318563 303996 318564 304060
rect 318628 303996 318629 304060
rect 318563 303995 318629 303996
rect 318011 286516 318077 286517
rect 318011 286452 318012 286516
rect 318076 286452 318077 286516
rect 318011 286451 318077 286452
rect 319302 224501 319362 317867
rect 322062 311949 322122 320179
rect 322246 319565 322306 320723
rect 322798 319701 322858 369411
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325371 320924 325437 320925
rect 325371 320860 325372 320924
rect 325436 320860 325437 320924
rect 325371 320859 325437 320860
rect 325374 320517 325434 320859
rect 325371 320516 325437 320517
rect 325371 320452 325372 320516
rect 325436 320452 325437 320516
rect 325371 320451 325437 320452
rect 323163 320380 323229 320381
rect 323163 320316 323164 320380
rect 323228 320316 323229 320380
rect 323163 320315 323229 320316
rect 322795 319700 322861 319701
rect 322795 319636 322796 319700
rect 322860 319636 322861 319700
rect 322795 319635 322861 319636
rect 323166 319565 323226 320315
rect 324083 320244 324149 320245
rect 324083 320180 324084 320244
rect 324148 320180 324149 320244
rect 324083 320179 324149 320180
rect 323347 320108 323413 320109
rect 323347 320044 323348 320108
rect 323412 320044 323413 320108
rect 323347 320043 323413 320044
rect 323899 320108 323965 320109
rect 323899 320044 323900 320108
rect 323964 320044 323965 320108
rect 323899 320043 323965 320044
rect 322243 319564 322309 319565
rect 322243 319500 322244 319564
rect 322308 319500 322309 319564
rect 322243 319499 322309 319500
rect 323163 319564 323229 319565
rect 323163 319500 323164 319564
rect 323228 319500 323229 319564
rect 323163 319499 323229 319500
rect 323350 319429 323410 320043
rect 323902 319429 323962 320043
rect 323347 319428 323413 319429
rect 323347 319364 323348 319428
rect 323412 319364 323413 319428
rect 323347 319363 323413 319364
rect 323899 319428 323965 319429
rect 323899 319364 323900 319428
rect 323964 319364 323965 319428
rect 323899 319363 323965 319364
rect 324086 319157 324146 320179
rect 324083 319156 324149 319157
rect 324083 319092 324084 319156
rect 324148 319092 324149 319156
rect 324083 319091 324149 319092
rect 322059 311948 322125 311949
rect 322059 311884 322060 311948
rect 322124 311884 322125 311948
rect 322059 311883 322125 311884
rect 322062 242181 322122 311883
rect 325794 291454 326414 326898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 328315 317524 328381 317525
rect 328315 317460 328316 317524
rect 328380 317460 328381 317524
rect 328315 317459 328381 317460
rect 328318 306390 328378 317459
rect 327582 306330 328378 306390
rect 327582 302293 327642 306330
rect 327579 302292 327645 302293
rect 327579 302228 327580 302292
rect 327644 302228 327645 302292
rect 327579 302227 327645 302228
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 322059 242180 322125 242181
rect 322059 242116 322060 242180
rect 322124 242116 322125 242180
rect 322059 242115 322125 242116
rect 319299 224500 319365 224501
rect 319299 224436 319300 224500
rect 319364 224436 319365 224500
rect 319299 224435 319365 224436
rect 325794 219454 326414 254898
rect 327582 243541 327642 302227
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 327579 243540 327645 243541
rect 327579 243476 327580 243540
rect 327644 243476 327645 243540
rect 327579 243475 327645 243476
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 317459 219060 317525 219061
rect 317459 218996 317460 219060
rect 317524 218996 317525 219060
rect 317459 218995 317525 218996
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 630334 341294 665778
rect 340674 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 341294 630334
rect 340674 630014 341294 630098
rect 340674 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 341294 630014
rect 340674 594334 341294 629778
rect 340674 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 341294 594334
rect 340674 594014 341294 594098
rect 340674 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 341294 594014
rect 340674 558334 341294 593778
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522334 341294 557778
rect 340674 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 341294 522334
rect 340674 522014 341294 522098
rect 340674 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 341294 522014
rect 340674 486334 341294 521778
rect 340674 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 341294 486334
rect 340674 486014 341294 486098
rect 340674 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 341294 486014
rect 340674 450334 341294 485778
rect 340674 450098 340706 450334
rect 340942 450098 341026 450334
rect 341262 450098 341294 450334
rect 340674 450014 341294 450098
rect 340674 449778 340706 450014
rect 340942 449778 341026 450014
rect 341262 449778 341294 450014
rect 340674 414334 341294 449778
rect 340674 414098 340706 414334
rect 340942 414098 341026 414334
rect 341262 414098 341294 414334
rect 340674 414014 341294 414098
rect 340674 413778 340706 414014
rect 340942 413778 341026 414014
rect 341262 413778 341294 414014
rect 340674 378334 341294 413778
rect 340674 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 341294 378334
rect 340674 378014 341294 378098
rect 340674 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 341294 378014
rect 340674 342334 341294 377778
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 306334 341294 341778
rect 340674 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 341294 306334
rect 340674 306014 341294 306098
rect 340674 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 341294 306014
rect 340674 270334 341294 305778
rect 340674 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 341294 270334
rect 340674 270014 341294 270098
rect 340674 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 341294 270014
rect 340674 234334 341294 269778
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 598054 345014 633498
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 344394 562054 345014 597498
rect 344394 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 345014 562054
rect 344394 561734 345014 561818
rect 344394 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 345014 561734
rect 344394 526054 345014 561498
rect 344394 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 345014 526054
rect 344394 525734 345014 525818
rect 344394 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 345014 525734
rect 344394 490054 345014 525498
rect 344394 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 345014 490054
rect 344394 489734 345014 489818
rect 344394 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 345014 489734
rect 344394 454054 345014 489498
rect 344394 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 345014 454054
rect 344394 453734 345014 453818
rect 344394 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 345014 453734
rect 344394 418054 345014 453498
rect 344394 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 345014 418054
rect 344394 417734 345014 417818
rect 344394 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 345014 417734
rect 344394 382054 345014 417498
rect 344394 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 345014 382054
rect 344394 381734 345014 381818
rect 344394 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 345014 381734
rect 344394 346054 345014 381498
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 344394 310054 345014 345498
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 344394 274054 345014 309498
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 344394 238054 345014 273498
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 348114 565774 348734 601218
rect 348114 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 348734 565774
rect 348114 565454 348734 565538
rect 348114 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 348734 565454
rect 348114 529774 348734 565218
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 348114 493774 348734 529218
rect 348114 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 348734 493774
rect 348114 493454 348734 493538
rect 348114 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 348734 493454
rect 348114 457774 348734 493218
rect 348114 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 348734 457774
rect 348114 457454 348734 457538
rect 348114 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 348734 457454
rect 348114 421774 348734 457218
rect 348114 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 348734 421774
rect 348114 421454 348734 421538
rect 348114 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 348734 421454
rect 348114 385774 348734 421218
rect 348114 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 348734 385774
rect 348114 385454 348734 385538
rect 348114 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 348734 385454
rect 348114 349774 348734 385218
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 348114 241774 348734 277218
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 351834 569494 352454 604938
rect 351834 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 352454 569494
rect 351834 569174 352454 569258
rect 351834 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 352454 569174
rect 351834 533494 352454 568938
rect 351834 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 352454 533494
rect 351834 533174 352454 533258
rect 351834 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 352454 533174
rect 351834 497494 352454 532938
rect 351834 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 352454 497494
rect 351834 497174 352454 497258
rect 351834 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 352454 497174
rect 351834 461494 352454 496938
rect 351834 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 352454 461494
rect 351834 461174 352454 461258
rect 351834 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 352454 461174
rect 351834 425494 352454 460938
rect 351834 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 352454 425494
rect 351834 425174 352454 425258
rect 351834 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 352454 425174
rect 351834 389494 352454 424938
rect 351834 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 352454 389494
rect 351834 389174 352454 389258
rect 351834 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 352454 389174
rect 351834 353494 352454 388938
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351834 245494 352454 280938
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 313774 420734 349218
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 133774 420734 169218
rect 420114 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 420734 133774
rect 420114 133454 420734 133538
rect 420114 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 420734 133454
rect 420114 97774 420734 133218
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 425494 424454 460938
rect 423834 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 424454 425494
rect 423834 425174 424454 425258
rect 423834 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 424454 425174
rect 423834 389494 424454 424938
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 423834 317494 424454 352938
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 423834 137494 424454 172938
rect 423834 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 424454 137494
rect 423834 137174 424454 137258
rect 423834 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 424454 137174
rect 423834 101494 424454 136938
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 306334 449294 341778
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 490054 453014 525498
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 452394 310054 453014 345498
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 493774 456734 529218
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 569494 460454 604938
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 497494 460454 532938
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 630334 485294 665778
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 486334 485294 521778
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 484674 414334 485294 449778
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 484674 378334 485294 413778
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 484674 342334 485294 377778
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 484674 306334 485294 341778
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 234334 485294 269778
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 484674 198334 485294 233778
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 634054 489014 669498
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 490054 489014 525498
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 488394 418054 489014 453498
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 488394 382054 489014 417498
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 488394 346054 489014 381498
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 488394 310054 489014 345498
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 238054 489014 273498
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 488394 202054 489014 237498
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 488394 166054 489014 201498
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 637774 492734 673218
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 601774 492734 637218
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 492114 565774 492734 601218
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 349774 492734 385218
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 492114 313774 492734 349218
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 241774 492734 277218
rect 492114 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 492734 241774
rect 492114 241454 492734 241538
rect 492114 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 492734 241454
rect 492114 205774 492734 241218
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 492114 169774 492734 205218
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 133774 492734 169218
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 492114 97774 492734 133218
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 641494 496454 676938
rect 495834 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 496454 641494
rect 495834 641174 496454 641258
rect 495834 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 496454 641174
rect 495834 605494 496454 640938
rect 495834 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 496454 605494
rect 495834 605174 496454 605258
rect 495834 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 496454 605174
rect 495834 569494 496454 604938
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 353494 496454 388938
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 495834 317494 496454 352938
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 245494 496454 280938
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 495834 209494 496454 244938
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 495834 173494 496454 208938
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 495834 137494 496454 172938
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 495834 101494 496454 136938
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 495834 65494 496454 100938
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 63866 605258 64102 605494
rect 64186 605258 64422 605494
rect 63866 604938 64102 605174
rect 64186 604938 64422 605174
rect 63866 569258 64102 569494
rect 64186 569258 64422 569494
rect 63866 568938 64102 569174
rect 64186 568938 64422 569174
rect 63866 533258 64102 533494
rect 64186 533258 64422 533494
rect 63866 532938 64102 533174
rect 64186 532938 64422 533174
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 88706 630098 88942 630334
rect 89026 630098 89262 630334
rect 88706 629778 88942 630014
rect 89026 629778 89262 630014
rect 88706 594098 88942 594334
rect 89026 594098 89262 594334
rect 88706 593778 88942 594014
rect 89026 593778 89262 594014
rect 88706 558098 88942 558334
rect 89026 558098 89262 558334
rect 88706 557778 88942 558014
rect 89026 557778 89262 558014
rect 88706 522098 88942 522334
rect 89026 522098 89262 522334
rect 88706 521778 88942 522014
rect 89026 521778 89262 522014
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 88706 234098 88942 234334
rect 89026 234098 89262 234334
rect 88706 233778 88942 234014
rect 89026 233778 89262 234014
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 88706 126098 88942 126334
rect 89026 126098 89262 126334
rect 88706 125778 88942 126014
rect 89026 125778 89262 126014
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 92426 597818 92662 598054
rect 92746 597818 92982 598054
rect 92426 597498 92662 597734
rect 92746 597498 92982 597734
rect 92426 561818 92662 562054
rect 92746 561818 92982 562054
rect 92426 561498 92662 561734
rect 92746 561498 92982 561734
rect 92426 525818 92662 526054
rect 92746 525818 92982 526054
rect 92426 525498 92662 525734
rect 92746 525498 92982 525734
rect 92426 489818 92662 490054
rect 92746 489818 92982 490054
rect 92426 489498 92662 489734
rect 92746 489498 92982 489734
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 92426 309818 92662 310054
rect 92746 309818 92982 310054
rect 92426 309498 92662 309734
rect 92746 309498 92982 309734
rect 92426 273818 92662 274054
rect 92746 273818 92982 274054
rect 92426 273498 92662 273734
rect 92746 273498 92982 273734
rect 92426 237818 92662 238054
rect 92746 237818 92982 238054
rect 92426 237498 92662 237734
rect 92746 237498 92982 237734
rect 92426 201818 92662 202054
rect 92746 201818 92982 202054
rect 92426 201498 92662 201734
rect 92746 201498 92982 201734
rect 92426 165818 92662 166054
rect 92746 165818 92982 166054
rect 92426 165498 92662 165734
rect 92746 165498 92982 165734
rect 92426 129818 92662 130054
rect 92746 129818 92982 130054
rect 92426 129498 92662 129734
rect 92746 129498 92982 129734
rect 92426 93818 92662 94054
rect 92746 93818 92982 94054
rect 92426 93498 92662 93734
rect 92746 93498 92982 93734
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 96146 601538 96382 601774
rect 96466 601538 96702 601774
rect 96146 601218 96382 601454
rect 96466 601218 96702 601454
rect 96146 565538 96382 565774
rect 96466 565538 96702 565774
rect 96146 565218 96382 565454
rect 96466 565218 96702 565454
rect 96146 529538 96382 529774
rect 96466 529538 96702 529774
rect 96146 529218 96382 529454
rect 96466 529218 96702 529454
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 96146 241538 96382 241774
rect 96466 241538 96702 241774
rect 96146 241218 96382 241454
rect 96466 241218 96702 241454
rect 96146 205538 96382 205774
rect 96466 205538 96702 205774
rect 96146 205218 96382 205454
rect 96466 205218 96702 205454
rect 96146 169538 96382 169774
rect 96466 169538 96702 169774
rect 96146 169218 96382 169454
rect 96466 169218 96702 169454
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 96146 97538 96382 97774
rect 96466 97538 96702 97774
rect 96146 97218 96382 97454
rect 96466 97218 96702 97454
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 99866 605258 100102 605494
rect 100186 605258 100422 605494
rect 99866 604938 100102 605174
rect 100186 604938 100422 605174
rect 99866 569258 100102 569494
rect 100186 569258 100422 569494
rect 99866 568938 100102 569174
rect 100186 568938 100422 569174
rect 99866 533258 100102 533494
rect 100186 533258 100422 533494
rect 99866 532938 100102 533174
rect 100186 532938 100422 533174
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 99866 281258 100102 281494
rect 100186 281258 100422 281494
rect 99866 280938 100102 281174
rect 100186 280938 100422 281174
rect 99866 245258 100102 245494
rect 100186 245258 100422 245494
rect 99866 244938 100102 245174
rect 100186 244938 100422 245174
rect 99866 209258 100102 209494
rect 100186 209258 100422 209494
rect 99866 208938 100102 209174
rect 100186 208938 100422 209174
rect 99866 173258 100102 173494
rect 100186 173258 100422 173494
rect 99866 172938 100102 173174
rect 100186 172938 100422 173174
rect 99866 137258 100102 137494
rect 100186 137258 100422 137494
rect 99866 136938 100102 137174
rect 100186 136938 100422 137174
rect 99866 101258 100102 101494
rect 100186 101258 100422 101494
rect 99866 100938 100102 101174
rect 100186 100938 100422 101174
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 124706 630098 124942 630334
rect 125026 630098 125262 630334
rect 124706 629778 124942 630014
rect 125026 629778 125262 630014
rect 124706 594098 124942 594334
rect 125026 594098 125262 594334
rect 124706 593778 124942 594014
rect 125026 593778 125262 594014
rect 124706 558098 124942 558334
rect 125026 558098 125262 558334
rect 124706 557778 124942 558014
rect 125026 557778 125262 558014
rect 124706 522098 124942 522334
rect 125026 522098 125262 522334
rect 124706 521778 124942 522014
rect 125026 521778 125262 522014
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 128426 597818 128662 598054
rect 128746 597818 128982 598054
rect 128426 597498 128662 597734
rect 128746 597498 128982 597734
rect 128426 561818 128662 562054
rect 128746 561818 128982 562054
rect 128426 561498 128662 561734
rect 128746 561498 128982 561734
rect 128426 525818 128662 526054
rect 128746 525818 128982 526054
rect 128426 525498 128662 525734
rect 128746 525498 128982 525734
rect 128426 489818 128662 490054
rect 128746 489818 128982 490054
rect 128426 489498 128662 489734
rect 128746 489498 128982 489734
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 128426 417818 128662 418054
rect 128746 417818 128982 418054
rect 128426 417498 128662 417734
rect 128746 417498 128982 417734
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 128426 129818 128662 130054
rect 128746 129818 128982 130054
rect 128426 129498 128662 129734
rect 128746 129498 128982 129734
rect 128426 93818 128662 94054
rect 128746 93818 128982 94054
rect 128426 93498 128662 93734
rect 128746 93498 128982 93734
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 132146 601538 132382 601774
rect 132466 601538 132702 601774
rect 132146 601218 132382 601454
rect 132466 601218 132702 601454
rect 132146 565538 132382 565774
rect 132466 565538 132702 565774
rect 132146 565218 132382 565454
rect 132466 565218 132702 565454
rect 132146 529538 132382 529774
rect 132466 529538 132702 529774
rect 132146 529218 132382 529454
rect 132466 529218 132702 529454
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 135866 605258 136102 605494
rect 136186 605258 136422 605494
rect 135866 604938 136102 605174
rect 136186 604938 136422 605174
rect 135866 569258 136102 569494
rect 136186 569258 136422 569494
rect 135866 568938 136102 569174
rect 136186 568938 136422 569174
rect 135866 533258 136102 533494
rect 136186 533258 136422 533494
rect 135866 532938 136102 533174
rect 136186 532938 136422 533174
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 164426 489818 164662 490054
rect 164746 489818 164982 490054
rect 164426 489498 164662 489734
rect 164746 489498 164982 489734
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 164426 417818 164662 418054
rect 164746 417818 164982 418054
rect 164426 417498 164662 417734
rect 164746 417498 164982 417734
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 171866 497258 172102 497494
rect 172186 497258 172422 497494
rect 171866 496938 172102 497174
rect 172186 496938 172422 497174
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 200426 597818 200662 598054
rect 200746 597818 200982 598054
rect 200426 597498 200662 597734
rect 200746 597498 200982 597734
rect 200426 561818 200662 562054
rect 200746 561818 200982 562054
rect 200426 561498 200662 561734
rect 200746 561498 200982 561734
rect 200426 525818 200662 526054
rect 200746 525818 200982 526054
rect 200426 525498 200662 525734
rect 200746 525498 200982 525734
rect 200426 489818 200662 490054
rect 200746 489818 200982 490054
rect 200426 489498 200662 489734
rect 200746 489498 200982 489734
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 200426 417818 200662 418054
rect 200746 417818 200982 418054
rect 200426 417498 200662 417734
rect 200746 417498 200982 417734
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 204146 601538 204382 601774
rect 204466 601538 204702 601774
rect 204146 601218 204382 601454
rect 204466 601218 204702 601454
rect 204146 565538 204382 565774
rect 204466 565538 204702 565774
rect 204146 565218 204382 565454
rect 204466 565218 204702 565454
rect 204146 529538 204382 529774
rect 204466 529538 204702 529774
rect 204146 529218 204382 529454
rect 204466 529218 204702 529454
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 224250 255218 224486 255454
rect 224250 254898 224486 255134
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 232706 594098 232942 594334
rect 233026 594098 233262 594334
rect 232706 593778 232942 594014
rect 233026 593778 233262 594014
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 232706 486098 232942 486334
rect 233026 486098 233262 486334
rect 232706 485778 232942 486014
rect 233026 485778 233262 486014
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 236426 597818 236662 598054
rect 236746 597818 236982 598054
rect 236426 597498 236662 597734
rect 236746 597498 236982 597734
rect 236426 561818 236662 562054
rect 236746 561818 236982 562054
rect 236426 561498 236662 561734
rect 236746 561498 236982 561734
rect 236426 525818 236662 526054
rect 236746 525818 236982 526054
rect 236426 525498 236662 525734
rect 236746 525498 236982 525734
rect 236426 489818 236662 490054
rect 236746 489818 236982 490054
rect 236426 489498 236662 489734
rect 236746 489498 236982 489734
rect 236426 453818 236662 454054
rect 236746 453818 236982 454054
rect 236426 453498 236662 453734
rect 236746 453498 236982 453734
rect 236426 417818 236662 418054
rect 236746 417818 236982 418054
rect 236426 417498 236662 417734
rect 236746 417498 236982 417734
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 240146 601538 240382 601774
rect 240466 601538 240702 601774
rect 240146 601218 240382 601454
rect 240466 601218 240702 601454
rect 240146 565538 240382 565774
rect 240466 565538 240702 565774
rect 240146 565218 240382 565454
rect 240466 565218 240702 565454
rect 240146 529538 240382 529774
rect 240466 529538 240702 529774
rect 240146 529218 240382 529454
rect 240466 529218 240702 529454
rect 240146 493538 240382 493774
rect 240466 493538 240702 493774
rect 240146 493218 240382 493454
rect 240466 493218 240702 493454
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 240146 421538 240382 421774
rect 240466 421538 240702 421774
rect 240146 421218 240382 421454
rect 240466 421218 240702 421454
rect 240146 385538 240382 385774
rect 240466 385538 240702 385774
rect 240146 385218 240382 385454
rect 240466 385218 240702 385454
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 243866 605258 244102 605494
rect 244186 605258 244422 605494
rect 243866 604938 244102 605174
rect 244186 604938 244422 605174
rect 243866 569258 244102 569494
rect 244186 569258 244422 569494
rect 243866 568938 244102 569174
rect 244186 568938 244422 569174
rect 243866 533258 244102 533494
rect 244186 533258 244422 533494
rect 243866 532938 244102 533174
rect 244186 532938 244422 533174
rect 243866 497258 244102 497494
rect 244186 497258 244422 497494
rect 243866 496938 244102 497174
rect 244186 496938 244422 497174
rect 243866 461258 244102 461494
rect 244186 461258 244422 461494
rect 243866 460938 244102 461174
rect 244186 460938 244422 461174
rect 243866 425258 244102 425494
rect 244186 425258 244422 425494
rect 243866 424938 244102 425174
rect 244186 424938 244422 425174
rect 243866 389258 244102 389494
rect 244186 389258 244422 389494
rect 243866 388938 244102 389174
rect 244186 388938 244422 389174
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 240146 313538 240382 313774
rect 240466 313538 240702 313774
rect 240146 313218 240382 313454
rect 240466 313218 240702 313454
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 240146 277538 240382 277774
rect 240466 277538 240702 277774
rect 240146 277218 240382 277454
rect 240466 277218 240702 277454
rect 239610 258938 239846 259174
rect 239610 258618 239846 258854
rect 240146 241538 240382 241774
rect 240466 241538 240702 241774
rect 240146 241218 240382 241454
rect 240466 241218 240702 241454
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 243866 281258 244102 281494
rect 244186 281258 244422 281494
rect 243866 280938 244102 281174
rect 244186 280938 244422 281174
rect 243866 245258 244102 245494
rect 244186 245258 244422 245494
rect 243866 244938 244102 245174
rect 244186 244938 244422 245174
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 254970 255218 255206 255454
rect 254970 254898 255206 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 268706 594098 268942 594334
rect 269026 594098 269262 594334
rect 268706 593778 268942 594014
rect 269026 593778 269262 594014
rect 268706 558098 268942 558334
rect 269026 558098 269262 558334
rect 268706 557778 268942 558014
rect 269026 557778 269262 558014
rect 268706 522098 268942 522334
rect 269026 522098 269262 522334
rect 268706 521778 268942 522014
rect 269026 521778 269262 522014
rect 268706 486098 268942 486334
rect 269026 486098 269262 486334
rect 268706 485778 268942 486014
rect 269026 485778 269262 486014
rect 268706 450098 268942 450334
rect 269026 450098 269262 450334
rect 268706 449778 268942 450014
rect 269026 449778 269262 450014
rect 268706 414098 268942 414334
rect 269026 414098 269262 414334
rect 268706 413778 268942 414014
rect 269026 413778 269262 414014
rect 268706 378098 268942 378334
rect 269026 378098 269262 378334
rect 268706 377778 268942 378014
rect 269026 377778 269262 378014
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 268706 306098 268942 306334
rect 269026 306098 269262 306334
rect 268706 305778 268942 306014
rect 269026 305778 269262 306014
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 272426 597818 272662 598054
rect 272746 597818 272982 598054
rect 272426 597498 272662 597734
rect 272746 597498 272982 597734
rect 272426 561818 272662 562054
rect 272746 561818 272982 562054
rect 272426 561498 272662 561734
rect 272746 561498 272982 561734
rect 272426 525818 272662 526054
rect 272746 525818 272982 526054
rect 272426 525498 272662 525734
rect 272746 525498 272982 525734
rect 272426 489818 272662 490054
rect 272746 489818 272982 490054
rect 272426 489498 272662 489734
rect 272746 489498 272982 489734
rect 272426 453818 272662 454054
rect 272746 453818 272982 454054
rect 272426 453498 272662 453734
rect 272746 453498 272982 453734
rect 272426 417818 272662 418054
rect 272746 417818 272982 418054
rect 272426 417498 272662 417734
rect 272746 417498 272982 417734
rect 272426 381818 272662 382054
rect 272746 381818 272982 382054
rect 272426 381498 272662 381734
rect 272746 381498 272982 381734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 276146 601538 276382 601774
rect 276466 601538 276702 601774
rect 276146 601218 276382 601454
rect 276466 601218 276702 601454
rect 276146 565538 276382 565774
rect 276466 565538 276702 565774
rect 276146 565218 276382 565454
rect 276466 565218 276702 565454
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 276146 493538 276382 493774
rect 276466 493538 276702 493774
rect 276146 493218 276382 493454
rect 276466 493218 276702 493454
rect 276146 457538 276382 457774
rect 276466 457538 276702 457774
rect 276146 457218 276382 457454
rect 276466 457218 276702 457454
rect 276146 421538 276382 421774
rect 276466 421538 276702 421774
rect 276146 421218 276382 421454
rect 276466 421218 276702 421454
rect 276146 385538 276382 385774
rect 276466 385538 276702 385774
rect 276146 385218 276382 385454
rect 276466 385218 276702 385454
rect 272426 345818 272662 346054
rect 272746 345818 272982 346054
rect 272426 345498 272662 345734
rect 272746 345498 272982 345734
rect 272426 309818 272662 310054
rect 272746 309818 272982 310054
rect 272426 309498 272662 309734
rect 272746 309498 272982 309734
rect 268706 270098 268942 270334
rect 269026 270098 269262 270334
rect 268706 269778 268942 270014
rect 269026 269778 269262 270014
rect 268706 234098 268942 234334
rect 269026 234098 269262 234334
rect 268706 233778 268942 234014
rect 269026 233778 269262 234014
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 198098 268942 198334
rect 269026 198098 269262 198334
rect 268706 197778 268942 198014
rect 269026 197778 269262 198014
rect 268706 162098 268942 162334
rect 269026 162098 269262 162334
rect 268706 161778 268942 162014
rect 269026 161778 269262 162014
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 279866 605258 280102 605494
rect 280186 605258 280422 605494
rect 279866 604938 280102 605174
rect 280186 604938 280422 605174
rect 279866 569258 280102 569494
rect 280186 569258 280422 569494
rect 279866 568938 280102 569174
rect 280186 568938 280422 569174
rect 279866 533258 280102 533494
rect 280186 533258 280422 533494
rect 279866 532938 280102 533174
rect 280186 532938 280422 533174
rect 279866 497258 280102 497494
rect 280186 497258 280422 497494
rect 279866 496938 280102 497174
rect 280186 496938 280422 497174
rect 279866 461258 280102 461494
rect 280186 461258 280422 461494
rect 279866 460938 280102 461174
rect 280186 460938 280422 461174
rect 279866 425258 280102 425494
rect 280186 425258 280422 425494
rect 279866 424938 280102 425174
rect 280186 424938 280422 425174
rect 279866 389258 280102 389494
rect 280186 389258 280422 389494
rect 279866 388938 280102 389174
rect 280186 388938 280422 389174
rect 276146 349538 276382 349774
rect 276466 349538 276702 349774
rect 276146 349218 276382 349454
rect 276466 349218 276702 349454
rect 276146 313538 276382 313774
rect 276466 313538 276702 313774
rect 276146 313218 276382 313454
rect 276466 313218 276702 313454
rect 272426 273818 272662 274054
rect 272746 273818 272982 274054
rect 272426 273498 272662 273734
rect 272746 273498 272982 273734
rect 272426 237818 272662 238054
rect 272746 237818 272982 238054
rect 272426 237498 272662 237734
rect 272746 237498 272982 237734
rect 272426 201818 272662 202054
rect 272746 201818 272982 202054
rect 272426 201498 272662 201734
rect 272746 201498 272982 201734
rect 272426 165818 272662 166054
rect 272746 165818 272982 166054
rect 272426 165498 272662 165734
rect 272746 165498 272982 165734
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 93818 272662 94054
rect 272746 93818 272982 94054
rect 272426 93498 272662 93734
rect 272746 93498 272982 93734
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 279866 353258 280102 353494
rect 280186 353258 280422 353494
rect 279866 352938 280102 353174
rect 280186 352938 280422 353174
rect 279866 317258 280102 317494
rect 280186 317258 280422 317494
rect 279866 316938 280102 317174
rect 280186 316938 280422 317174
rect 276146 277538 276382 277774
rect 276466 277538 276702 277774
rect 276146 277218 276382 277454
rect 276466 277218 276702 277454
rect 276146 241538 276382 241774
rect 276466 241538 276702 241774
rect 276146 241218 276382 241454
rect 276466 241218 276702 241454
rect 276146 205538 276382 205774
rect 276466 205538 276702 205774
rect 276146 205218 276382 205454
rect 276466 205218 276702 205454
rect 276146 169538 276382 169774
rect 276466 169538 276702 169774
rect 276146 169218 276382 169454
rect 276466 169218 276702 169454
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 281258 280102 281494
rect 280186 281258 280422 281494
rect 279866 280938 280102 281174
rect 280186 280938 280422 281174
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 304706 630098 304942 630334
rect 305026 630098 305262 630334
rect 304706 629778 304942 630014
rect 305026 629778 305262 630014
rect 304706 594098 304942 594334
rect 305026 594098 305262 594334
rect 304706 593778 304942 594014
rect 305026 593778 305262 594014
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 304706 522098 304942 522334
rect 305026 522098 305262 522334
rect 304706 521778 304942 522014
rect 305026 521778 305262 522014
rect 304706 486098 304942 486334
rect 305026 486098 305262 486334
rect 304706 485778 304942 486014
rect 305026 485778 305262 486014
rect 304706 450098 304942 450334
rect 305026 450098 305262 450334
rect 304706 449778 304942 450014
rect 305026 449778 305262 450014
rect 304706 414098 304942 414334
rect 305026 414098 305262 414334
rect 304706 413778 304942 414014
rect 305026 413778 305262 414014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 308426 597818 308662 598054
rect 308746 597818 308982 598054
rect 308426 597498 308662 597734
rect 308746 597498 308982 597734
rect 308426 561818 308662 562054
rect 308746 561818 308982 562054
rect 308426 561498 308662 561734
rect 308746 561498 308982 561734
rect 308426 525818 308662 526054
rect 308746 525818 308982 526054
rect 308426 525498 308662 525734
rect 308746 525498 308982 525734
rect 308426 489818 308662 490054
rect 308746 489818 308982 490054
rect 308426 489498 308662 489734
rect 308746 489498 308982 489734
rect 308426 453818 308662 454054
rect 308746 453818 308982 454054
rect 308426 453498 308662 453734
rect 308746 453498 308982 453734
rect 308426 417818 308662 418054
rect 308746 417818 308982 418054
rect 308426 417498 308662 417734
rect 308746 417498 308982 417734
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 312146 601538 312382 601774
rect 312466 601538 312702 601774
rect 312146 601218 312382 601454
rect 312466 601218 312702 601454
rect 312146 565538 312382 565774
rect 312466 565538 312702 565774
rect 312146 565218 312382 565454
rect 312466 565218 312702 565454
rect 312146 529538 312382 529774
rect 312466 529538 312702 529774
rect 312146 529218 312382 529454
rect 312466 529218 312702 529454
rect 312146 493538 312382 493774
rect 312466 493538 312702 493774
rect 312146 493218 312382 493454
rect 312466 493218 312702 493454
rect 312146 457538 312382 457774
rect 312466 457538 312702 457774
rect 312146 457218 312382 457454
rect 312466 457218 312702 457454
rect 312146 421538 312382 421774
rect 312466 421538 312702 421774
rect 312146 421218 312382 421454
rect 312466 421218 312702 421454
rect 308426 381818 308662 382054
rect 308746 381818 308982 382054
rect 308426 381498 308662 381734
rect 308746 381498 308982 381734
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 315866 605258 316102 605494
rect 316186 605258 316422 605494
rect 315866 604938 316102 605174
rect 316186 604938 316422 605174
rect 315866 569258 316102 569494
rect 316186 569258 316422 569494
rect 315866 568938 316102 569174
rect 316186 568938 316422 569174
rect 315866 533258 316102 533494
rect 316186 533258 316422 533494
rect 315866 532938 316102 533174
rect 316186 532938 316422 533174
rect 315866 497258 316102 497494
rect 316186 497258 316422 497494
rect 315866 496938 316102 497174
rect 316186 496938 316422 497174
rect 315866 461258 316102 461494
rect 316186 461258 316422 461494
rect 315866 460938 316102 461174
rect 316186 460938 316422 461174
rect 315866 425258 316102 425494
rect 316186 425258 316422 425494
rect 315866 424938 316102 425174
rect 316186 424938 316422 425174
rect 312146 385538 312382 385774
rect 312466 385538 312702 385774
rect 312146 385218 312382 385454
rect 312466 385218 312702 385454
rect 308426 345818 308662 346054
rect 308746 345818 308982 346054
rect 308426 345498 308662 345734
rect 308746 345498 308982 345734
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 308426 309818 308662 310054
rect 308746 309818 308982 310054
rect 308426 309498 308662 309734
rect 308746 309498 308982 309734
rect 308426 273818 308662 274054
rect 308746 273818 308982 274054
rect 308426 273498 308662 273734
rect 308746 273498 308982 273734
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 315866 389258 316102 389494
rect 316186 389258 316422 389494
rect 315866 388938 316102 389174
rect 316186 388938 316422 389174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 308426 93818 308662 94054
rect 308746 93818 308982 94054
rect 308426 93498 308662 93734
rect 308746 93498 308982 93734
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 340706 630098 340942 630334
rect 341026 630098 341262 630334
rect 340706 629778 340942 630014
rect 341026 629778 341262 630014
rect 340706 594098 340942 594334
rect 341026 594098 341262 594334
rect 340706 593778 340942 594014
rect 341026 593778 341262 594014
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 340706 522098 340942 522334
rect 341026 522098 341262 522334
rect 340706 521778 340942 522014
rect 341026 521778 341262 522014
rect 340706 486098 340942 486334
rect 341026 486098 341262 486334
rect 340706 485778 340942 486014
rect 341026 485778 341262 486014
rect 340706 450098 340942 450334
rect 341026 450098 341262 450334
rect 340706 449778 340942 450014
rect 341026 449778 341262 450014
rect 340706 414098 340942 414334
rect 341026 414098 341262 414334
rect 340706 413778 340942 414014
rect 341026 413778 341262 414014
rect 340706 378098 340942 378334
rect 341026 378098 341262 378334
rect 340706 377778 340942 378014
rect 341026 377778 341262 378014
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 340706 306098 340942 306334
rect 341026 306098 341262 306334
rect 340706 305778 340942 306014
rect 341026 305778 341262 306014
rect 340706 270098 340942 270334
rect 341026 270098 341262 270334
rect 340706 269778 340942 270014
rect 341026 269778 341262 270014
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 344426 561818 344662 562054
rect 344746 561818 344982 562054
rect 344426 561498 344662 561734
rect 344746 561498 344982 561734
rect 344426 525818 344662 526054
rect 344746 525818 344982 526054
rect 344426 525498 344662 525734
rect 344746 525498 344982 525734
rect 344426 489818 344662 490054
rect 344746 489818 344982 490054
rect 344426 489498 344662 489734
rect 344746 489498 344982 489734
rect 344426 453818 344662 454054
rect 344746 453818 344982 454054
rect 344426 453498 344662 453734
rect 344746 453498 344982 453734
rect 344426 417818 344662 418054
rect 344746 417818 344982 418054
rect 344426 417498 344662 417734
rect 344746 417498 344982 417734
rect 344426 381818 344662 382054
rect 344746 381818 344982 382054
rect 344426 381498 344662 381734
rect 344746 381498 344982 381734
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 348146 565538 348382 565774
rect 348466 565538 348702 565774
rect 348146 565218 348382 565454
rect 348466 565218 348702 565454
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 348146 493538 348382 493774
rect 348466 493538 348702 493774
rect 348146 493218 348382 493454
rect 348466 493218 348702 493454
rect 348146 457538 348382 457774
rect 348466 457538 348702 457774
rect 348146 457218 348382 457454
rect 348466 457218 348702 457454
rect 348146 421538 348382 421774
rect 348466 421538 348702 421774
rect 348146 421218 348382 421454
rect 348466 421218 348702 421454
rect 348146 385538 348382 385774
rect 348466 385538 348702 385774
rect 348146 385218 348382 385454
rect 348466 385218 348702 385454
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 351866 569258 352102 569494
rect 352186 569258 352422 569494
rect 351866 568938 352102 569174
rect 352186 568938 352422 569174
rect 351866 533258 352102 533494
rect 352186 533258 352422 533494
rect 351866 532938 352102 533174
rect 352186 532938 352422 533174
rect 351866 497258 352102 497494
rect 352186 497258 352422 497494
rect 351866 496938 352102 497174
rect 352186 496938 352422 497174
rect 351866 461258 352102 461494
rect 352186 461258 352422 461494
rect 351866 460938 352102 461174
rect 352186 460938 352422 461174
rect 351866 425258 352102 425494
rect 352186 425258 352422 425494
rect 351866 424938 352102 425174
rect 352186 424938 352422 425174
rect 351866 389258 352102 389494
rect 352186 389258 352422 389494
rect 351866 388938 352102 389174
rect 352186 388938 352422 389174
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 420146 133538 420382 133774
rect 420466 133538 420702 133774
rect 420146 133218 420382 133454
rect 420466 133218 420702 133454
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 423866 425258 424102 425494
rect 424186 425258 424422 425494
rect 423866 424938 424102 425174
rect 424186 424938 424422 425174
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 423866 137258 424102 137494
rect 424186 137258 424422 137494
rect 423866 136938 424102 137174
rect 424186 136938 424422 137174
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 492146 241538 492382 241774
rect 492466 241538 492702 241774
rect 492146 241218 492382 241454
rect 492466 241218 492702 241454
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 495866 641258 496102 641494
rect 496186 641258 496422 641494
rect 495866 640938 496102 641174
rect 496186 640938 496422 641174
rect 495866 605258 496102 605494
rect 496186 605258 496422 605494
rect 495866 604938 496102 605174
rect 496186 604938 496422 605174
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 92426 598054
rect 92662 597818 92746 598054
rect 92982 597818 128426 598054
rect 128662 597818 128746 598054
rect 128982 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 92426 597734
rect 92662 597498 92746 597734
rect 92982 597498 128426 597734
rect 128662 597498 128746 597734
rect 128982 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 88706 594334
rect 88942 594098 89026 594334
rect 89262 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 88706 594014
rect 88942 593778 89026 594014
rect 89262 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 99866 569494
rect 100102 569258 100186 569494
rect 100422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 99866 569174
rect 100102 568938 100186 569174
rect 100422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 96146 565774
rect 96382 565538 96466 565774
rect 96702 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 96146 565454
rect 96382 565218 96466 565454
rect 96702 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 92426 562054
rect 92662 561818 92746 562054
rect 92982 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 92426 561734
rect 92662 561498 92746 561734
rect 92982 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 340706 450334
rect 340942 450098 341026 450334
rect 341262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 340706 450014
rect 340942 449778 341026 450014
rect 341262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 272426 418054
rect 272662 417818 272746 418054
rect 272982 417818 308426 418054
rect 308662 417818 308746 418054
rect 308982 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 272426 417734
rect 272662 417498 272746 417734
rect 272982 417498 308426 417734
rect 308662 417498 308746 417734
rect 308982 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 340706 414334
rect 340942 414098 341026 414334
rect 341262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 340706 414014
rect 340942 413778 341026 414014
rect 341262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 272426 310054
rect 272662 309818 272746 310054
rect 272982 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 272426 309734
rect 272662 309498 272746 309734
rect 272982 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 276146 277774
rect 276382 277538 276466 277774
rect 276702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 276146 277454
rect 276382 277218 276466 277454
rect 276702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 272426 274054
rect 272662 273818 272746 274054
rect 272982 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 272426 273734
rect 272662 273498 272746 273734
rect 272982 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 268706 270334
rect 268942 270098 269026 270334
rect 269262 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 268706 270014
rect 268942 269778 269026 270014
rect 269262 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 239610 259174
rect 239846 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 239610 258854
rect 239846 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 224250 255454
rect 224486 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254970 255454
rect 255206 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 224250 255134
rect 224486 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254970 255134
rect 255206 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use macro_2to3  u_macro_2to3
timestamp 0
transform 1 0 280000 0 1 320000
box 1066 0 48890 50000
use macro_2xdrive  u_macro_2xdrive
timestamp 0
transform 1 0 220000 0 1 240000
box 1066 0 48890 50000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 255088 255336 255088 255336 0 vccd1
rlabel via4 261704 262776 261704 262776 0 vccd2
rlabel via4 269144 270216 269144 270216 0 vdda1
rlabel via4 240584 277656 240584 277656 0 vdda2
rlabel via4 236864 273936 236864 273936 0 vssa1
rlabel via4 244304 281376 244304 281376 0 vssa2
rlabel via4 257984 259056 257984 259056 0 vssd1
rlabel via4 265424 266496 265424 266496 0 vssd2
rlabel metal3 581908 6596 581908 6596 0 io_in[0]
rlabel metal2 235382 290894 235382 290894 0 io_in[10]
rlabel metal2 236433 289884 236433 289884 0 io_in[11]
rlabel metal2 237590 290928 237590 290928 0 io_in[12]
rlabel metal2 238595 289884 238595 289884 0 io_in[13]
rlabel metal2 330510 525436 330510 525436 0 io_in[14]
rlabel metal2 558946 539247 558946 539247 0 io_in[15]
rlabel metal2 241907 289884 241907 289884 0 io_in[16]
rlabel metal2 429456 703596 429456 703596 0 io_in[17]
rlabel metal2 364366 537887 364366 537887 0 io_in[18]
rlabel metal3 302565 386308 302565 386308 0 io_in[19]
rlabel metal3 581954 46308 581954 46308 0 io_in[1]
rlabel metal2 248446 371246 248446 371246 0 io_in[20]
rlabel metal2 169786 539876 169786 539876 0 io_in[21]
rlabel metal2 105110 703596 105110 703596 0 io_in[22]
rlabel metal2 40204 703596 40204 703596 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 1878 632060 1878 632060 0 io_in[25]
rlabel metal3 1878 579972 1878 579972 0 io_in[26]
rlabel metal3 1556 527884 1556 527884 0 io_in[27]
rlabel metal2 255155 289884 255155 289884 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal2 256174 290632 256174 290632 0 io_in[2]
rlabel metal3 1878 371348 1878 371348 0 io_in[30]
rlabel metal3 1878 319260 1878 319260 0 io_in[31]
rlabel metal2 232254 291006 232254 291006 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal3 1786 162860 1786 162860 0 io_in[34]
rlabel metal3 1878 110636 1878 110636 0 io_in[35]
rlabel metal3 1878 71604 1878 71604 0 io_in[36]
rlabel metal3 1878 32436 1878 32436 0 io_in[37]
rlabel metal3 583556 125732 583556 125732 0 io_in[3]
rlabel metal3 582092 165852 582092 165852 0 io_in[4]
rlabel metal2 229809 289884 229809 289884 0 io_in[5]
rlabel metal2 230966 290554 230966 290554 0 io_in[6]
rlabel metal2 232070 290928 232070 290928 0 io_in[7]
rlabel metal2 233075 289612 233075 289612 0 io_in[8]
rlabel metal2 234278 290962 234278 290962 0 io_in[9]
rlabel metal3 583556 32368 583556 32368 0 io_oeb[0]
rlabel metal2 235750 292254 235750 292254 0 io_oeb[10]
rlabel metal2 236755 289884 236755 289884 0 io_oeb[11]
rlabel metal2 237859 289884 237859 289884 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal1 526838 699686 526838 699686 0 io_oeb[15]
rlabel metal2 462346 546696 462346 546696 0 io_oeb[16]
rlabel metal2 243379 289884 243379 289884 0 io_oeb[17]
rlabel metal1 331890 703018 331890 703018 0 io_oeb[18]
rlabel metal1 267030 697578 267030 697578 0 io_oeb[19]
rlabel metal2 580198 73049 580198 73049 0 io_oeb[1]
rlabel metal2 306544 383640 306544 383640 0 io_oeb[20]
rlabel metal2 137172 703596 137172 703596 0 io_oeb[21]
rlabel metal1 72404 703018 72404 703018 0 io_oeb[22]
rlabel metal2 309258 386045 309258 386045 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal1 251712 293046 251712 293046 0 io_oeb[25]
rlabel metal1 252954 293046 252954 293046 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1740 449548 1740 449548 0 io_oeb[28]
rlabel metal2 256871 289748 256871 289748 0 io_oeb[29]
rlabel metal2 231150 334169 231150 334169 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 1878 241060 1878 241060 0 io_oeb[32]
rlabel metal3 1924 188836 1924 188836 0 io_oeb[33]
rlabel metal3 1602 136748 1602 136748 0 io_oeb[34]
rlabel metal3 1740 84660 1740 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal1 578634 193154 578634 193154 0 io_oeb[4]
rlabel metal2 230131 289884 230131 289884 0 io_oeb[5]
rlabel metal2 231235 289884 231235 289884 0 io_oeb[6]
rlabel metal2 232339 289884 232339 289884 0 io_oeb[7]
rlabel metal2 233443 289884 233443 289884 0 io_oeb[8]
rlabel metal2 579922 431103 579922 431103 0 io_oeb[9]
rlabel metal2 580198 20213 580198 20213 0 io_out[0]
rlabel metal2 236118 291642 236118 291642 0 io_out[10]
rlabel metal2 237123 289884 237123 289884 0 io_out[11]
rlabel metal2 238326 291200 238326 291200 0 io_out[12]
rlabel metal2 580198 630751 580198 630751 0 io_out[13]
rlabel metal2 580198 683553 580198 683553 0 io_out[14]
rlabel metal2 542386 548189 542386 548189 0 io_out[15]
rlabel metal2 242742 292339 242742 292339 0 io_out[16]
rlabel metal2 403650 549202 403650 549202 0 io_out[17]
rlabel metal2 348818 701940 348818 701940 0 io_out[18]
rlabel metal1 294446 700298 294446 700298 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 219006 701260 219006 701260 0 io_out[20]
rlabel metal1 154698 700094 154698 700094 0 io_out[21]
rlabel metal1 89792 699686 89792 699686 0 io_out[22]
rlabel metal1 250056 293046 250056 293046 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1786 566916 1786 566916 0 io_out[26]
rlabel metal2 254787 289884 254787 289884 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 1602 410516 1602 410516 0 io_out[29]
rlabel metal2 579646 100079 579646 100079 0 io_out[2]
rlabel metal3 1878 358428 1878 358428 0 io_out[30]
rlabel metal3 1786 306204 1786 306204 0 io_out[31]
rlabel metal3 1878 254116 1878 254116 0 io_out[32]
rlabel metal3 1924 201892 1924 201892 0 io_out[33]
rlabel metal3 1878 149804 1878 149804 0 io_out[34]
rlabel metal3 1878 97580 1878 97580 0 io_out[35]
rlabel metal3 1694 58548 1694 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel metal3 581954 139332 581954 139332 0 io_out[3]
rlabel metal1 578634 179350 578634 179350 0 io_out[4]
rlabel metal3 582046 219028 582046 219028 0 io_out[5]
rlabel metal2 231702 291710 231702 291710 0 io_out[6]
rlabel metal2 232707 289884 232707 289884 0 io_out[7]
rlabel metal2 233910 291744 233910 291744 0 io_out[8]
rlabel metal2 235014 291030 235014 291030 0 io_out[9]
rlabel metal2 125757 340 125757 340 0 la_data_in[0]
rlabel metal2 480562 2234 480562 2234 0 la_data_in[100]
rlabel metal2 483552 16560 483552 16560 0 la_data_in[101]
rlabel metal2 487409 340 487409 340 0 la_data_in[102]
rlabel metal2 328394 231472 328394 231472 0 la_data_in[103]
rlabel metal1 413540 236810 413540 236810 0 la_data_in[104]
rlabel metal2 498226 1911 498226 1911 0 la_data_in[105]
rlabel metal2 332718 219062 332718 219062 0 la_data_in[106]
rlabel metal2 505402 1962 505402 1962 0 la_data_in[107]
rlabel metal2 508898 1911 508898 1911 0 la_data_in[108]
rlabel metal2 512249 340 512249 340 0 la_data_in[109]
rlabel metal2 161322 2064 161322 2064 0 la_data_in[10]
rlabel metal2 331522 233087 331522 233087 0 la_data_in[110]
rlabel metal2 329774 212126 329774 212126 0 la_data_in[111]
rlabel metal2 523066 1843 523066 1843 0 la_data_in[112]
rlabel metal2 526417 340 526417 340 0 la_data_in[113]
rlabel metal2 527850 16864 527850 16864 0 la_data_in[114]
rlabel metal2 336674 234192 336674 234192 0 la_data_in[115]
rlabel metal2 334834 230044 334834 230044 0 la_data_in[116]
rlabel metal2 540822 2132 540822 2132 0 la_data_in[117]
rlabel metal2 334834 223108 334834 223108 0 la_data_in[118]
rlabel metal2 334006 237014 334006 237014 0 la_data_in[119]
rlabel metal2 164910 2098 164910 2098 0 la_data_in[11]
rlabel metal2 331522 235552 331522 235552 0 la_data_in[120]
rlabel metal1 429732 236742 429732 236742 0 la_data_in[121]
rlabel metal2 558072 16560 558072 16560 0 la_data_in[122]
rlabel metal2 562074 1894 562074 1894 0 la_data_in[123]
rlabel metal2 565662 1826 565662 1826 0 la_data_in[124]
rlabel metal2 568921 340 568921 340 0 la_data_in[125]
rlabel metal2 565110 110364 565110 110364 0 la_data_in[126]
rlabel metal2 328394 216240 328394 216240 0 la_data_in[127]
rlabel metal2 168406 959 168406 959 0 la_data_in[12]
rlabel metal2 171994 2166 171994 2166 0 la_data_in[13]
rlabel metal2 175398 16560 175398 16560 0 la_data_in[14]
rlabel metal2 178841 340 178841 340 0 la_data_in[15]
rlabel metal2 182383 340 182383 340 0 la_data_in[16]
rlabel metal1 213210 3536 213210 3536 0 la_data_in[17]
rlabel metal2 191130 117912 191130 117912 0 la_data_in[18]
rlabel metal2 193246 891 193246 891 0 la_data_in[19]
rlabel metal2 210450 121822 210450 121822 0 la_data_in[1]
rlabel metal2 196420 16560 196420 16560 0 la_data_in[20]
rlabel metal2 200238 16560 200238 16560 0 la_data_in[21]
rlabel metal2 203681 340 203681 340 0 la_data_in[22]
rlabel metal2 213394 278324 213394 278324 0 la_data_in[23]
rlabel metal1 294722 311134 294722 311134 0 la_data_in[24]
rlabel metal2 214222 16560 214222 16560 0 la_data_in[25]
rlabel metal2 218086 117188 218086 117188 0 la_data_in[26]
rlabel metal2 221345 340 221345 340 0 la_data_in[27]
rlabel metal1 232346 216138 232346 216138 0 la_data_in[28]
rlabel metal2 228521 340 228521 340 0 la_data_in[29]
rlabel metal2 132756 16560 132756 16560 0 la_data_in[2]
rlabel metal2 232063 340 232063 340 0 la_data_in[30]
rlabel metal2 235842 1911 235842 1911 0 la_data_in[31]
rlabel metal2 239062 16560 239062 16560 0 la_data_in[32]
rlabel metal2 242926 1894 242926 1894 0 la_data_in[33]
rlabel metal2 246185 340 246185 340 0 la_data_in[34]
rlabel metal2 250010 2234 250010 2234 0 la_data_in[35]
rlabel metal2 253506 2030 253506 2030 0 la_data_in[36]
rlabel metal2 257094 2166 257094 2166 0 la_data_in[37]
rlabel metal2 260682 2200 260682 2200 0 la_data_in[38]
rlabel metal2 264178 1860 264178 1860 0 la_data_in[39]
rlabel metal2 136482 1860 136482 1860 0 la_data_in[3]
rlabel metal2 267766 1928 267766 1928 0 la_data_in[40]
rlabel metal2 271071 340 271071 340 0 la_data_in[41]
rlabel metal2 274850 1996 274850 1996 0 la_data_in[42]
rlabel metal2 275954 119646 275954 119646 0 la_data_in[43]
rlabel metal2 281743 340 281743 340 0 la_data_in[44]
rlabel metal1 273056 3570 273056 3570 0 la_data_in[45]
rlabel metal2 289018 2166 289018 2166 0 la_data_in[46]
rlabel metal1 274942 233818 274942 233818 0 la_data_in[47]
rlabel metal2 296102 1962 296102 1962 0 la_data_in[48]
rlabel metal1 296355 3434 296355 3434 0 la_data_in[49]
rlabel metal2 139833 340 139833 340 0 la_data_in[4]
rlabel metal2 302726 16560 302726 16560 0 la_data_in[50]
rlabel metal2 306774 1996 306774 1996 0 la_data_in[51]
rlabel metal2 310033 340 310033 340 0 la_data_in[52]
rlabel metal2 313858 1928 313858 1928 0 la_data_in[53]
rlabel metal2 313950 118796 313950 118796 0 la_data_in[54]
rlabel metal2 307602 231370 307602 231370 0 la_data_in[55]
rlabel metal2 303738 232458 303738 232458 0 la_data_in[56]
rlabel metal2 328026 1911 328026 1911 0 la_data_in[57]
rlabel metal2 331614 2166 331614 2166 0 la_data_in[58]
rlabel metal2 334873 340 334873 340 0 la_data_in[59]
rlabel metal2 143566 117120 143566 117120 0 la_data_in[5]
rlabel metal2 305302 225420 305302 225420 0 la_data_in[60]
rlabel metal1 331660 223482 331660 223482 0 la_data_in[61]
rlabel metal2 345545 340 345545 340 0 la_data_in[62]
rlabel metal2 349278 108212 349278 108212 0 la_data_in[63]
rlabel metal2 352866 1690 352866 1690 0 la_data_in[64]
rlabel metal2 310454 232832 310454 232832 0 la_data_in[65]
rlabel metal2 359713 340 359713 340 0 la_data_in[66]
rlabel metal2 339434 221850 339434 221850 0 la_data_in[67]
rlabel metal2 367034 2200 367034 2200 0 la_data_in[68]
rlabel metal2 370385 340 370385 340 0 la_data_in[69]
rlabel metal2 146740 16560 146740 16560 0 la_data_in[6]
rlabel metal2 311282 230010 311282 230010 0 la_data_in[70]
rlabel metal2 334190 227392 334190 227392 0 la_data_in[71]
rlabel metal2 322966 223210 322966 223210 0 la_data_in[72]
rlabel metal2 328394 214948 328394 214948 0 la_data_in[73]
rlabel metal2 388286 2030 388286 2030 0 la_data_in[74]
rlabel metal2 391874 1860 391874 1860 0 la_data_in[75]
rlabel via3 303485 219164 303485 219164 0 la_data_in[76]
rlabel metal2 320758 213588 320758 213588 0 la_data_in[77]
rlabel metal1 383640 3842 383640 3842 0 la_data_in[78]
rlabel metal2 405904 16560 405904 16560 0 la_data_in[79]
rlabel metal2 150558 16560 150558 16560 0 la_data_in[7]
rlabel metal2 409630 1724 409630 1724 0 la_data_in[80]
rlabel metal2 313306 221714 313306 221714 0 la_data_in[81]
rlabel metal1 296194 217974 296194 217974 0 la_data_in[82]
rlabel metal2 338054 210800 338054 210800 0 la_data_in[83]
rlabel metal2 423798 1826 423798 1826 0 la_data_in[84]
rlabel metal2 427057 340 427057 340 0 la_data_in[85]
rlabel metal2 430744 16560 430744 16560 0 la_data_in[86]
rlabel metal2 425730 106624 425730 106624 0 la_data_in[87]
rlabel metal2 437966 1860 437966 1860 0 la_data_in[88]
rlabel metal3 316020 229772 316020 229772 0 la_data_in[89]
rlabel metal2 154238 1690 154238 1690 0 la_data_in[8]
rlabel metal2 445050 1860 445050 1860 0 la_data_in[90]
rlabel metal2 448638 1690 448638 1690 0 la_data_in[91]
rlabel metal2 334098 214948 334098 214948 0 la_data_in[92]
rlabel metal2 307694 213520 307694 213520 0 la_data_in[93]
rlabel metal2 458712 16560 458712 16560 0 la_data_in[94]
rlabel metal2 462569 340 462569 340 0 la_data_in[95]
rlabel metal2 466065 340 466065 340 0 la_data_in[96]
rlabel metal2 469890 1860 469890 1860 0 la_data_in[97]
rlabel metal2 473478 1690 473478 1690 0 la_data_in[98]
rlabel metal2 320114 210698 320114 210698 0 la_data_in[99]
rlabel metal2 157596 16560 157596 16560 0 la_data_in[9]
rlabel metal1 179814 157998 179814 157998 0 la_data_out[0]
rlabel metal2 481758 3627 481758 3627 0 la_data_out[100]
rlabel metal2 485254 1996 485254 1996 0 la_data_out[101]
rlabel metal2 488704 16560 488704 16560 0 la_data_out[102]
rlabel metal1 320850 245718 320850 245718 0 la_data_out[103]
rlabel metal2 329038 229080 329038 229080 0 la_data_out[104]
rlabel metal1 320850 271830 320850 271830 0 la_data_out[105]
rlabel metal2 503010 1911 503010 1911 0 la_data_out[106]
rlabel metal2 506506 125790 506506 125790 0 la_data_out[107]
rlabel metal2 508530 158015 508530 158015 0 la_data_out[108]
rlabel metal2 513590 1622 513590 1622 0 la_data_out[109]
rlabel metal2 162281 340 162281 340 0 la_data_out[10]
rlabel metal1 327750 3536 327750 3536 0 la_data_out[110]
rlabel metal3 329038 231812 329038 231812 0 la_data_out[111]
rlabel metal2 524071 340 524071 340 0 la_data_out[112]
rlabel metal2 527850 1928 527850 1928 0 la_data_out[113]
rlabel metal2 531346 2030 531346 2030 0 la_data_out[114]
rlabel metal2 534697 340 534697 340 0 la_data_out[115]
rlabel metal2 538331 340 538331 340 0 la_data_out[116]
rlabel metal2 541512 16560 541512 16560 0 la_data_out[117]
rlabel metal2 545514 1724 545514 1724 0 la_data_out[118]
rlabel metal2 548865 340 548865 340 0 la_data_out[119]
rlabel metal2 235382 208735 235382 208735 0 la_data_out[11]
rlabel metal2 552690 1996 552690 1996 0 la_data_out[120]
rlabel metal2 556186 1962 556186 1962 0 la_data_out[121]
rlabel metal2 559537 340 559537 340 0 la_data_out[122]
rlabel metal2 563171 340 563171 340 0 la_data_out[123]
rlabel metal2 315606 273921 315606 273921 0 la_data_out[124]
rlabel metal2 570170 16560 570170 16560 0 la_data_out[125]
rlabel metal3 296585 271116 296585 271116 0 la_data_out[126]
rlabel metal2 577438 2098 577438 2098 0 la_data_out[127]
rlabel metal2 169602 1860 169602 1860 0 la_data_out[12]
rlabel metal2 172953 340 172953 340 0 la_data_out[13]
rlabel metal2 176686 3627 176686 3627 0 la_data_out[14]
rlabel metal2 179860 16560 179860 16560 0 la_data_out[15]
rlabel metal2 183678 16560 183678 16560 0 la_data_out[16]
rlabel metal2 187121 340 187121 340 0 la_data_out[17]
rlabel metal2 190663 340 190663 340 0 la_data_out[18]
rlabel metal2 194442 1860 194442 1860 0 la_data_out[19]
rlabel metal2 130180 16560 130180 16560 0 la_data_out[1]
rlabel metal2 197662 16560 197662 16560 0 la_data_out[20]
rlabel metal2 201526 3627 201526 3627 0 la_data_out[21]
rlabel metal2 204700 16560 204700 16560 0 la_data_out[22]
rlabel metal2 208518 16560 208518 16560 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215694 1928 215694 1928 0 la_data_out[25]
rlabel metal2 219282 1911 219282 1911 0 la_data_out[26]
rlabel metal2 222502 16560 222502 16560 0 la_data_out[27]
rlabel metal2 234002 105570 234002 105570 0 la_data_out[28]
rlabel metal2 229862 1894 229862 1894 0 la_data_out[29]
rlabel metal2 134037 340 134037 340 0 la_data_out[2]
rlabel metal2 233358 16560 233358 16560 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal2 240343 340 240343 340 0 la_data_out[32]
rlabel metal2 244122 1928 244122 1928 0 la_data_out[33]
rlabel metal2 247342 16560 247342 16560 0 la_data_out[34]
rlabel metal2 251206 1860 251206 1860 0 la_data_out[35]
rlabel metal2 254702 1860 254702 1860 0 la_data_out[36]
rlabel metal2 258198 16560 258198 16560 0 la_data_out[37]
rlabel metal2 261786 1996 261786 1996 0 la_data_out[38]
rlabel metal2 265374 2064 265374 2064 0 la_data_out[39]
rlabel metal2 137441 340 137441 340 0 la_data_out[3]
rlabel metal2 268633 340 268633 340 0 la_data_out[40]
rlabel metal2 272458 1928 272458 1928 0 la_data_out[41]
rlabel metal2 276046 1928 276046 1928 0 la_data_out[42]
rlabel metal2 279305 340 279305 340 0 la_data_out[43]
rlabel metal2 283038 16560 283038 16560 0 la_data_out[44]
rlabel metal1 294722 307394 294722 307394 0 la_data_out[45]
rlabel metal2 290214 1928 290214 1928 0 la_data_out[46]
rlabel metal2 293473 340 293473 340 0 la_data_out[47]
rlabel metal2 298034 230758 298034 230758 0 la_data_out[48]
rlabel metal2 300794 1894 300794 1894 0 la_data_out[49]
rlabel metal2 141036 16560 141036 16560 0 la_data_out[4]
rlabel metal2 304145 340 304145 340 0 la_data_out[50]
rlabel metal2 253322 231523 253322 231523 0 la_data_out[51]
rlabel metal2 311466 1911 311466 1911 0 la_data_out[52]
rlabel metal2 315054 1758 315054 1758 0 la_data_out[53]
rlabel metal2 315146 229080 315146 229080 0 la_data_out[54]
rlabel metal2 321862 16560 321862 16560 0 la_data_out[55]
rlabel metal2 325634 1928 325634 1928 0 la_data_out[56]
rlabel metal2 329222 1894 329222 1894 0 la_data_out[57]
rlabel metal2 307602 236878 307602 236878 0 la_data_out[58]
rlabel metal1 330280 226338 330280 226338 0 la_data_out[59]
rlabel metal1 291272 310454 291272 310454 0 la_data_out[5]
rlabel metal1 330464 4046 330464 4046 0 la_data_out[60]
rlabel metal1 331660 226338 331660 226338 0 la_data_out[61]
rlabel metal2 346702 16560 346702 16560 0 la_data_out[62]
rlabel metal2 350474 1860 350474 1860 0 la_data_out[63]
rlabel metal2 354062 2200 354062 2200 0 la_data_out[64]
rlabel metal1 338054 4046 338054 4046 0 la_data_out[65]
rlabel metal2 361146 1622 361146 1622 0 la_data_out[66]
rlabel metal2 364504 16560 364504 16560 0 la_data_out[67]
rlabel metal2 367993 340 367993 340 0 la_data_out[68]
rlabel metal2 371489 340 371489 340 0 la_data_out[69]
rlabel metal2 148113 340 148113 340 0 la_data_out[6]
rlabel metal2 375314 1860 375314 1860 0 la_data_out[70]
rlabel metal2 378665 340 378665 340 0 la_data_out[71]
rlabel metal1 312478 293998 312478 293998 0 la_data_out[72]
rlabel metal2 385986 1911 385986 1911 0 la_data_out[73]
rlabel metal2 312846 242097 312846 242097 0 la_data_out[74]
rlabel metal2 392833 340 392833 340 0 la_data_out[75]
rlabel metal2 396329 340 396329 340 0 la_data_out[76]
rlabel metal2 314318 237184 314318 237184 0 la_data_out[77]
rlabel metal1 313904 259386 313904 259386 0 la_data_out[78]
rlabel metal2 407238 1775 407238 1775 0 la_data_out[79]
rlabel metal2 151846 108892 151846 108892 0 la_data_out[7]
rlabel metal2 289386 268124 289386 268124 0 la_data_out[80]
rlabel metal1 364090 311134 364090 311134 0 la_data_out[81]
rlabel metal1 314456 308414 314456 308414 0 la_data_out[82]
rlabel metal1 314732 253946 314732 253946 0 la_data_out[83]
rlabel metal2 424994 1860 424994 1860 0 la_data_out[84]
rlabel metal2 428168 16560 428168 16560 0 la_data_out[85]
rlabel metal2 280968 310284 280968 310284 0 la_data_out[86]
rlabel metal3 310017 253980 310017 253980 0 la_data_out[87]
rlabel metal1 289984 224434 289984 224434 0 la_data_out[88]
rlabel metal2 442152 16560 442152 16560 0 la_data_out[89]
rlabel metal2 155434 2030 155434 2030 0 la_data_out[8]
rlabel metal2 446009 340 446009 340 0 la_data_out[90]
rlabel metal2 449834 2574 449834 2574 0 la_data_out[91]
rlabel metal2 329682 301512 329682 301512 0 la_data_out[92]
rlabel metal2 456918 1775 456918 1775 0 la_data_out[93]
rlabel metal2 460414 3424 460414 3424 0 la_data_out[94]
rlabel metal2 463864 16560 463864 16560 0 la_data_out[95]
rlabel metal2 466992 16560 466992 16560 0 la_data_out[96]
rlabel metal1 326807 291890 326807 291890 0 la_data_out[97]
rlabel metal3 335340 236776 335340 236776 0 la_data_out[98]
rlabel metal2 478170 1911 478170 1911 0 la_data_out[99]
rlabel metal2 158838 16560 158838 16560 0 la_data_out[9]
rlabel metal1 127604 11798 127604 11798 0 la_oenb[0]
rlabel metal2 482625 340 482625 340 0 la_oenb[100]
rlabel metal2 486450 1843 486450 1843 0 la_oenb[101]
rlabel metal1 296010 238782 296010 238782 0 la_oenb[102]
rlabel metal2 493297 340 493297 340 0 la_oenb[103]
rlabel metal1 291042 224706 291042 224706 0 la_oenb[104]
rlabel metal2 500618 1911 500618 1911 0 la_oenb[105]
rlabel metal2 503969 340 503969 340 0 la_oenb[106]
rlabel metal2 507465 340 507465 340 0 la_oenb[107]
rlabel metal1 416300 252586 416300 252586 0 la_oenb[108]
rlabel metal3 388953 191012 388953 191012 0 la_oenb[109]
rlabel metal1 292008 307530 292008 307530 0 la_oenb[10]
rlabel metal1 304152 307122 304152 307122 0 la_oenb[110]
rlabel metal2 521771 340 521771 340 0 la_oenb[111]
rlabel metal2 525458 1792 525458 1792 0 la_oenb[112]
rlabel metal2 528809 340 528809 340 0 la_oenb[113]
rlabel metal2 532542 1690 532542 1690 0 la_oenb[114]
rlabel metal3 264569 221204 264569 221204 0 la_oenb[115]
rlabel metal2 539626 3627 539626 3627 0 la_oenb[116]
rlabel metal2 542977 340 542977 340 0 la_oenb[117]
rlabel metal2 546611 340 546611 340 0 la_oenb[118]
rlabel metal2 547170 109276 547170 109276 0 la_oenb[119]
rlabel metal2 235566 217464 235566 217464 0 la_oenb[11]
rlabel metal2 324898 205224 324898 205224 0 la_oenb[120]
rlabel metal2 557382 1928 557382 1928 0 la_oenb[121]
rlabel metal2 560878 1928 560878 1928 0 la_oenb[122]
rlabel metal2 564466 3627 564466 3627 0 la_oenb[123]
rlabel metal2 563730 89964 563730 89964 0 la_oenb[124]
rlabel metal3 297298 272476 297298 272476 0 la_oenb[125]
rlabel metal2 575138 1911 575138 1911 0 la_oenb[126]
rlabel metal2 578450 16560 578450 16560 0 la_oenb[127]
rlabel metal3 235681 289612 235681 289612 0 la_oenb[12]
rlabel metal2 174103 340 174103 340 0 la_oenb[13]
rlabel metal1 177284 11798 177284 11798 0 la_oenb[14]
rlabel metal2 236118 221238 236118 221238 0 la_oenb[15]
rlabel metal2 184966 118803 184966 118803 0 la_oenb[16]
rlabel metal2 237222 219606 237222 219606 0 la_oenb[17]
rlabel metal2 191958 16560 191958 16560 0 la_oenb[18]
rlabel metal2 195401 340 195401 340 0 la_oenb[19]
rlabel metal4 232484 221680 232484 221680 0 la_oenb[1]
rlabel metal2 199134 2234 199134 2234 0 la_oenb[20]
rlabel metal3 238372 306884 238372 306884 0 la_oenb[21]
rlabel metal1 238004 233886 238004 233886 0 la_oenb[22]
rlabel metal2 209806 3627 209806 3627 0 la_oenb[23]
rlabel metal2 213394 1911 213394 1911 0 la_oenb[24]
rlabel metal2 216798 16560 216798 16560 0 la_oenb[25]
rlabel metal2 220241 340 220241 340 0 la_oenb[26]
rlabel metal2 223974 1724 223974 1724 0 la_oenb[27]
rlabel metal2 238694 293488 238694 293488 0 la_oenb[28]
rlabel metal2 231058 3627 231058 3627 0 la_oenb[29]
rlabel metal2 135286 2030 135286 2030 0 la_oenb[2]
rlabel metal3 270365 305660 270365 305660 0 la_oenb[30]
rlabel metal2 237905 340 237905 340 0 la_oenb[31]
rlabel metal2 241638 16560 241638 16560 0 la_oenb[32]
rlabel metal2 245226 1911 245226 1911 0 la_oenb[33]
rlabel metal2 248814 1792 248814 1792 0 la_oenb[34]
rlabel metal2 252402 1911 252402 1911 0 la_oenb[35]
rlabel metal2 255622 16560 255622 16560 0 la_oenb[36]
rlabel metal2 259486 1911 259486 1911 0 la_oenb[37]
rlabel metal2 262745 340 262745 340 0 la_oenb[38]
rlabel metal1 243708 234022 243708 234022 0 la_oenb[39]
rlabel metal2 138874 1911 138874 1911 0 la_oenb[3]
rlabel metal2 270066 1911 270066 1911 0 la_oenb[40]
rlabel metal2 273463 340 273463 340 0 la_oenb[41]
rlabel metal2 277150 1724 277150 1724 0 la_oenb[42]
rlabel metal2 281198 214200 281198 214200 0 la_oenb[43]
rlabel metal2 284326 231132 284326 231132 0 la_oenb[44]
rlabel metal2 287822 1894 287822 1894 0 la_oenb[45]
rlabel metal2 291410 1894 291410 1894 0 la_oenb[46]
rlabel metal2 294446 16560 294446 16560 0 la_oenb[47]
rlabel metal2 298303 340 298303 340 0 la_oenb[48]
rlabel metal2 301990 1928 301990 1928 0 la_oenb[49]
rlabel metal4 233956 213512 233956 213512 0 la_oenb[4]
rlabel metal3 275655 213180 275655 213180 0 la_oenb[50]
rlabel metal2 309074 1928 309074 1928 0 la_oenb[51]
rlabel metal2 312662 1962 312662 1962 0 la_oenb[52]
rlabel metal3 281497 152388 281497 152388 0 la_oenb[53]
rlabel metal2 307694 210732 307694 210732 0 la_oenb[54]
rlabel metal2 323143 340 323143 340 0 la_oenb[55]
rlabel metal2 326830 1860 326830 1860 0 la_oenb[56]
rlabel metal2 330142 16560 330142 16560 0 la_oenb[57]
rlabel metal2 333914 3203 333914 3203 0 la_oenb[58]
rlabel metal2 337265 340 337265 340 0 la_oenb[59]
rlabel metal2 145721 340 145721 340 0 la_oenb[5]
rlabel metal3 279059 311780 279059 311780 0 la_oenb[60]
rlabel metal3 279795 311508 279795 311508 0 la_oenb[61]
rlabel metal2 347944 16560 347944 16560 0 la_oenb[62]
rlabel metal2 351433 340 351433 340 0 la_oenb[63]
rlabel metal3 280485 222972 280485 222972 0 la_oenb[64]
rlabel metal1 280324 311406 280324 311406 0 la_oenb[65]
rlabel metal1 281152 311202 281152 311202 0 la_oenb[66]
rlabel metal2 365838 69503 365838 69503 0 la_oenb[67]
rlabel metal2 369426 4648 369426 4648 0 la_oenb[68]
rlabel metal2 372922 2132 372922 2132 0 la_oenb[69]
rlabel metal2 233910 116935 233910 116935 0 la_oenb[6]
rlabel metal2 376510 2098 376510 2098 0 la_oenb[70]
rlabel metal2 380006 1979 380006 1979 0 la_oenb[71]
rlabel metal3 282463 309468 282463 309468 0 la_oenb[72]
rlabel metal2 386945 340 386945 340 0 la_oenb[73]
rlabel metal2 390678 1095 390678 1095 0 la_oenb[74]
rlabel metal2 394266 3390 394266 3390 0 la_oenb[75]
rlabel metal2 397762 3356 397762 3356 0 la_oenb[76]
rlabel metal3 283705 310012 283705 310012 0 la_oenb[77]
rlabel metal2 404846 3543 404846 3543 0 la_oenb[78]
rlabel metal1 313858 269042 313858 269042 0 la_oenb[79]
rlabel metal2 153042 1860 153042 1860 0 la_oenb[7]
rlabel via2 313306 222955 313306 222955 0 la_oenb[80]
rlabel metal2 255162 223431 255162 223431 0 la_oenb[81]
rlabel metal1 282440 309502 282440 309502 0 la_oenb[82]
rlabel metal2 422602 7402 422602 7402 0 la_oenb[83]
rlabel metal2 426190 3475 426190 3475 0 la_oenb[84]
rlabel metal3 256013 290020 256013 290020 0 la_oenb[85]
rlabel metal3 255967 289748 255967 289748 0 la_oenb[86]
rlabel metal3 256243 289612 256243 289612 0 la_oenb[87]
rlabel metal3 286327 287708 286327 287708 0 la_oenb[88]
rlabel metal2 443617 340 443617 340 0 la_oenb[89]
rlabel metal2 156393 340 156393 340 0 la_oenb[8]
rlabel metal4 256772 196520 256772 196520 0 la_oenb[90]
rlabel metal4 256956 186184 256956 186184 0 la_oenb[91]
rlabel metal3 287385 290428 287385 290428 0 la_oenb[92]
rlabel metal3 271101 218620 271101 218620 0 la_oenb[93]
rlabel metal2 461610 3254 461610 3254 0 la_oenb[94]
rlabel metal2 465198 3271 465198 3271 0 la_oenb[95]
rlabel metal2 468457 340 468457 340 0 la_oenb[96]
rlabel metal3 272757 218484 272757 218484 0 la_oenb[97]
rlabel metal3 289547 308380 289547 308380 0 la_oenb[98]
rlabel metal1 290398 219130 290398 219130 0 la_oenb[99]
rlabel metal2 160126 1996 160126 1996 0 la_oenb[9]
rlabel metal2 1702 1962 1702 1962 0 wb_rst_i
rlabel metal2 2898 2166 2898 2166 0 wbs_ack_o
rlabel metal2 21390 102816 21390 102816 0 wbs_adr_i[0]
rlabel metal2 47649 340 47649 340 0 wbs_adr_i[10]
rlabel metal2 51237 340 51237 340 0 wbs_adr_i[11]
rlabel metal2 54970 1911 54970 1911 0 wbs_adr_i[12]
rlabel metal2 58236 16560 58236 16560 0 wbs_adr_i[13]
rlabel metal2 62054 2098 62054 2098 0 wbs_adr_i[14]
rlabel metal2 65313 340 65313 340 0 wbs_adr_i[15]
rlabel metal2 287178 309281 287178 309281 0 wbs_adr_i[16]
rlabel metal2 213670 274924 213670 274924 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 12183 340 12183 340 0 wbs_adr_i[1]
rlabel metal2 83076 16560 83076 16560 0 wbs_adr_i[20]
rlabel metal2 214682 273190 214682 273190 0 wbs_adr_i[21]
rlabel metal2 213578 273479 213578 273479 0 wbs_adr_i[22]
rlabel metal2 93978 3627 93978 3627 0 wbs_adr_i[23]
rlabel metal2 97474 1911 97474 1911 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 104321 340 104321 340 0 wbs_adr_i[26]
rlabel metal1 254886 309842 254886 309842 0 wbs_adr_i[27]
rlabel metal2 214866 269824 214866 269824 0 wbs_adr_i[28]
rlabel metal2 114993 340 114993 340 0 wbs_adr_i[29]
rlabel metal2 17066 1690 17066 1690 0 wbs_adr_i[2]
rlabel metal2 231610 217566 231610 217566 0 wbs_adr_i[30]
rlabel metal2 122314 1911 122314 1911 0 wbs_adr_i[31]
rlabel metal2 21850 1928 21850 1928 0 wbs_adr_i[3]
rlabel metal2 26397 340 26397 340 0 wbs_adr_i[4]
rlabel metal1 126546 213214 126546 213214 0 wbs_adr_i[5]
rlabel metal2 215050 276148 215050 276148 0 wbs_adr_i[6]
rlabel metal2 37023 340 37023 340 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 210726 234872 210726 234872 0 wbs_adr_i[9]
rlabel metal2 3857 340 3857 340 0 wbs_cyc_i
rlabel metal2 8556 16560 8556 16560 0 wbs_dat_i[0]
rlabel metal2 48990 1928 48990 1928 0 wbs_dat_i[10]
rlabel metal2 55890 107848 55890 107848 0 wbs_dat_i[11]
rlabel metal2 56074 1911 56074 1911 0 wbs_dat_i[12]
rlabel metal2 59662 1962 59662 1962 0 wbs_dat_i[13]
rlabel metal2 63250 1911 63250 1911 0 wbs_dat_i[14]
rlabel metal3 146625 196588 146625 196588 0 wbs_dat_i[15]
rlabel metal2 70097 340 70097 340 0 wbs_dat_i[16]
rlabel metal2 75210 99688 75210 99688 0 wbs_dat_i[17]
rlabel metal2 77418 1826 77418 1826 0 wbs_dat_i[18]
rlabel metal2 80500 16560 80500 16560 0 wbs_dat_i[19]
rlabel metal2 13570 1928 13570 1928 0 wbs_dat_i[1]
rlabel metal1 227838 233240 227838 233240 0 wbs_dat_i[20]
rlabel metal1 229724 222122 229724 222122 0 wbs_dat_i[21]
rlabel metal2 230230 216818 230230 216818 0 wbs_dat_i[22]
rlabel metal2 94937 340 94937 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102212 16560 102212 16560 0 wbs_dat_i[25]
rlabel metal4 231196 211472 231196 211472 0 wbs_dat_i[26]
rlabel metal1 231058 228106 231058 228106 0 wbs_dat_i[27]
rlabel metal2 112601 340 112601 340 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18117 340 18117 340 0 wbs_dat_i[2]
rlabel metal3 231380 218076 231380 218076 0 wbs_dat_i[30]
rlabel metal2 152490 119425 152490 119425 0 wbs_dat_i[31]
rlabel metal2 22809 340 22809 340 0 wbs_dat_i[3]
rlabel metal2 27738 1792 27738 1792 0 wbs_dat_i[4]
rlabel metal2 214774 271864 214774 271864 0 wbs_dat_i[5]
rlabel metal2 212014 271796 212014 271796 0 wbs_dat_i[6]
rlabel metal2 38410 1928 38410 1928 0 wbs_dat_i[7]
rlabel metal2 41906 2030 41906 2030 0 wbs_dat_i[8]
rlabel metal2 45494 2234 45494 2234 0 wbs_dat_i[9]
rlabel metal2 9837 340 9837 340 0 wbs_dat_o[0]
rlabel metal2 212290 278392 212290 278392 0 wbs_dat_o[10]
rlabel metal2 53774 1962 53774 1962 0 wbs_dat_o[11]
rlabel metal2 57270 1996 57270 1996 0 wbs_dat_o[12]
rlabel metal2 60812 16560 60812 16560 0 wbs_dat_o[13]
rlabel metal2 64354 1758 64354 1758 0 wbs_dat_o[14]
rlabel metal2 67797 340 67797 340 0 wbs_dat_o[15]
rlabel metal2 71530 1911 71530 1911 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78614 2574 78614 2574 0 wbs_dat_o[18]
rlabel metal2 81873 340 81873 340 0 wbs_dat_o[19]
rlabel metal2 14766 1962 14766 1962 0 wbs_dat_o[1]
rlabel metal3 232507 289748 232507 289748 0 wbs_dat_o[20]
rlabel metal2 89194 1860 89194 1860 0 wbs_dat_o[21]
rlabel metal2 212474 235654 212474 235654 0 wbs_dat_o[22]
rlabel metal2 96278 1996 96278 1996 0 wbs_dat_o[23]
rlabel metal2 99406 16899 99406 16899 0 wbs_dat_o[24]
rlabel metal1 230092 233818 230092 233818 0 wbs_dat_o[25]
rlabel metal2 106713 340 106713 340 0 wbs_dat_o[26]
rlabel metal2 110538 5328 110538 5328 0 wbs_dat_o[27]
rlabel metal2 114034 1860 114034 1860 0 wbs_dat_o[28]
rlabel metal2 117622 3254 117622 3254 0 wbs_dat_o[29]
rlabel metal2 19458 3627 19458 3627 0 wbs_dat_o[2]
rlabel metal2 121118 1996 121118 1996 0 wbs_dat_o[30]
rlabel metal2 124706 1758 124706 1758 0 wbs_dat_o[31]
rlabel metal2 23506 17579 23506 17579 0 wbs_dat_o[3]
rlabel metal2 213394 129778 213394 129778 0 wbs_dat_o[4]
rlabel metal2 32193 340 32193 340 0 wbs_dat_o[5]
rlabel metal2 36018 82610 36018 82610 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 42957 340 42957 340 0 wbs_dat_o[8]
rlabel metal2 175950 119510 175950 119510 0 wbs_dat_o[9]
rlabel metal2 11178 45346 11178 45346 0 wbs_sel_i[0]
rlabel metal2 15962 1911 15962 1911 0 wbs_sel_i[1]
rlabel metal2 20463 340 20463 340 0 wbs_sel_i[2]
rlabel metal2 25346 6722 25346 6722 0 wbs_sel_i[3]
rlabel metal2 4738 16560 4738 16560 0 wbs_stb_i
rlabel metal2 6486 1894 6486 1894 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
