magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 5792 263 6326 535
<< pwell >>
rect 459 2661 545 2677
rect 459 2654 885 2661
rect 72 2240 885 2654
rect 459 861 885 2240
rect 459 10 920 861
<< mvnmos >>
rect 98 2475 398 2575
rect 98 2319 398 2419
rect 594 682 894 782
rect 594 526 894 626
rect 594 245 894 345
rect 594 89 894 189
<< mvpmos >>
rect 5911 329 6031 469
rect 6087 329 6207 469
<< mvnnmos >>
rect 659 1863 859 2043
rect 659 1627 859 1807
rect 659 1270 859 1450
rect 659 1034 859 1214
<< nmoslvt >>
rect 659 2552 859 2582
rect 659 2466 859 2496
rect 659 2380 859 2410
rect 659 2294 859 2324
<< ndiff >>
rect 659 2627 859 2635
rect 659 2593 671 2627
rect 705 2593 739 2627
rect 773 2593 807 2627
rect 841 2593 859 2627
rect 659 2582 859 2593
rect 659 2541 859 2552
rect 659 2507 671 2541
rect 705 2507 739 2541
rect 773 2507 807 2541
rect 841 2507 859 2541
rect 659 2496 859 2507
rect 659 2455 859 2466
rect 659 2421 671 2455
rect 705 2421 739 2455
rect 773 2421 807 2455
rect 841 2421 859 2455
rect 659 2410 859 2421
rect 659 2369 859 2380
rect 659 2335 671 2369
rect 705 2335 739 2369
rect 773 2335 807 2369
rect 841 2335 859 2369
rect 659 2324 859 2335
rect 659 2283 859 2294
rect 659 2249 671 2283
rect 705 2249 739 2283
rect 773 2249 807 2283
rect 841 2249 859 2283
rect 659 2241 859 2249
<< mvndiff >>
rect 98 2620 398 2628
rect 98 2586 148 2620
rect 182 2586 216 2620
rect 250 2586 284 2620
rect 318 2586 352 2620
rect 386 2586 398 2620
rect 98 2575 398 2586
rect 98 2464 398 2475
rect 98 2430 148 2464
rect 182 2430 216 2464
rect 250 2430 284 2464
rect 318 2430 352 2464
rect 386 2430 398 2464
rect 98 2419 398 2430
rect 98 2308 398 2319
rect 98 2274 148 2308
rect 182 2274 216 2308
rect 250 2274 284 2308
rect 318 2274 352 2308
rect 386 2274 398 2308
rect 98 2266 398 2274
rect 659 2088 859 2096
rect 659 2054 671 2088
rect 705 2054 739 2088
rect 773 2054 807 2088
rect 841 2054 859 2088
rect 659 2043 859 2054
rect 659 1852 859 1863
rect 659 1818 671 1852
rect 705 1818 739 1852
rect 773 1818 807 1852
rect 841 1818 859 1852
rect 659 1807 859 1818
rect 659 1616 859 1627
rect 659 1582 671 1616
rect 705 1582 739 1616
rect 773 1582 807 1616
rect 841 1582 859 1616
rect 659 1574 859 1582
rect 659 1495 859 1503
rect 659 1461 677 1495
rect 711 1461 745 1495
rect 779 1461 813 1495
rect 847 1461 859 1495
rect 659 1450 859 1461
rect 659 1259 859 1270
rect 659 1225 677 1259
rect 711 1225 745 1259
rect 779 1225 813 1259
rect 847 1225 859 1259
rect 659 1214 859 1225
rect 659 1023 859 1034
rect 659 989 677 1023
rect 711 989 745 1023
rect 779 989 813 1023
rect 847 989 859 1023
rect 659 981 859 989
rect 594 827 894 835
rect 594 793 606 827
rect 640 793 674 827
rect 708 793 742 827
rect 776 793 810 827
rect 844 793 894 827
rect 594 782 894 793
rect 594 671 894 682
rect 594 637 606 671
rect 640 637 674 671
rect 708 637 742 671
rect 776 637 810 671
rect 844 637 894 671
rect 594 626 894 637
rect 594 515 894 526
rect 594 481 606 515
rect 640 481 674 515
rect 708 481 742 515
rect 776 481 810 515
rect 844 481 894 515
rect 594 473 894 481
rect 594 390 894 398
rect 594 356 606 390
rect 640 356 674 390
rect 708 356 742 390
rect 776 356 810 390
rect 844 356 894 390
rect 594 345 894 356
rect 594 234 894 245
rect 594 200 606 234
rect 640 200 674 234
rect 708 200 742 234
rect 776 200 810 234
rect 844 200 894 234
rect 594 189 894 200
rect 594 78 894 89
rect 594 44 606 78
rect 640 44 674 78
rect 708 44 742 78
rect 776 44 810 78
rect 844 44 894 78
rect 594 36 894 44
<< mvpdiff >>
rect 5858 457 5911 469
rect 5858 423 5866 457
rect 5900 423 5911 457
rect 5858 389 5911 423
rect 5858 355 5866 389
rect 5900 355 5911 389
rect 5858 329 5911 355
rect 6031 457 6087 469
rect 6031 423 6042 457
rect 6076 423 6087 457
rect 6031 389 6087 423
rect 6031 355 6042 389
rect 6076 355 6087 389
rect 6031 329 6087 355
rect 6207 457 6260 469
rect 6207 423 6218 457
rect 6252 423 6260 457
rect 6207 389 6260 423
rect 6207 355 6218 389
rect 6252 355 6260 389
rect 6207 329 6260 355
<< ndiffc >>
rect 671 2593 705 2627
rect 739 2593 773 2627
rect 807 2593 841 2627
rect 671 2507 705 2541
rect 739 2507 773 2541
rect 807 2507 841 2541
rect 671 2421 705 2455
rect 739 2421 773 2455
rect 807 2421 841 2455
rect 671 2335 705 2369
rect 739 2335 773 2369
rect 807 2335 841 2369
rect 671 2249 705 2283
rect 739 2249 773 2283
rect 807 2249 841 2283
<< mvndiffc >>
rect 148 2586 182 2620
rect 216 2586 250 2620
rect 284 2586 318 2620
rect 352 2586 386 2620
rect 148 2430 182 2464
rect 216 2430 250 2464
rect 284 2430 318 2464
rect 352 2430 386 2464
rect 148 2274 182 2308
rect 216 2274 250 2308
rect 284 2274 318 2308
rect 352 2274 386 2308
rect 671 2054 705 2088
rect 739 2054 773 2088
rect 807 2054 841 2088
rect 671 1818 705 1852
rect 739 1818 773 1852
rect 807 1818 841 1852
rect 671 1582 705 1616
rect 739 1582 773 1616
rect 807 1582 841 1616
rect 677 1461 711 1495
rect 745 1461 779 1495
rect 813 1461 847 1495
rect 677 1225 711 1259
rect 745 1225 779 1259
rect 813 1225 847 1259
rect 677 989 711 1023
rect 745 989 779 1023
rect 813 989 847 1023
rect 606 793 640 827
rect 674 793 708 827
rect 742 793 776 827
rect 810 793 844 827
rect 606 637 640 671
rect 674 637 708 671
rect 742 637 776 671
rect 810 637 844 671
rect 606 481 640 515
rect 674 481 708 515
rect 742 481 776 515
rect 810 481 844 515
rect 606 356 640 390
rect 674 356 708 390
rect 742 356 776 390
rect 810 356 844 390
rect 606 200 640 234
rect 674 200 708 234
rect 742 200 776 234
rect 810 200 844 234
rect 606 44 640 78
rect 674 44 708 78
rect 742 44 776 78
rect 810 44 844 78
<< mvpdiffc >>
rect 5866 423 5900 457
rect 5866 355 5900 389
rect 6042 423 6076 457
rect 6042 355 6076 389
rect 6218 423 6252 457
rect 6218 355 6252 389
<< psubdiff >>
rect 485 2627 519 2651
rect 485 2559 519 2593
rect 485 2491 519 2525
rect 485 2423 519 2457
rect 485 2355 519 2389
rect 485 2287 519 2321
rect 485 2219 519 2253
rect 485 2151 519 2185
rect 485 2083 519 2117
rect 485 2015 519 2049
rect 485 1947 519 1981
rect 485 1879 519 1913
rect 485 1811 519 1845
rect 485 1743 519 1777
rect 485 1675 519 1709
rect 485 1607 519 1641
rect 485 1539 519 1573
rect 485 1471 519 1505
rect 485 1403 519 1437
rect 485 1335 519 1369
rect 485 1267 519 1301
rect 485 1198 519 1233
rect 485 1129 519 1164
rect 485 1060 519 1095
rect 485 991 519 1026
rect 485 922 519 957
rect 485 853 519 888
rect 485 784 519 819
rect 485 715 519 750
rect 485 646 519 681
rect 485 577 519 612
rect 485 508 519 543
rect 485 439 519 474
rect 485 370 519 405
rect 485 301 519 336
rect 485 232 519 267
rect 485 163 519 198
rect 485 94 519 129
rect 485 36 519 60
<< psubdiffcont >>
rect 485 2593 519 2627
rect 485 2525 519 2559
rect 485 2457 519 2491
rect 485 2389 519 2423
rect 485 2321 519 2355
rect 485 2253 519 2287
rect 485 2185 519 2219
rect 485 2117 519 2151
rect 485 2049 519 2083
rect 485 1981 519 2015
rect 485 1913 519 1947
rect 485 1845 519 1879
rect 485 1777 519 1811
rect 485 1709 519 1743
rect 485 1641 519 1675
rect 485 1573 519 1607
rect 485 1505 519 1539
rect 485 1437 519 1471
rect 485 1369 519 1403
rect 485 1301 519 1335
rect 485 1233 519 1267
rect 485 1164 519 1198
rect 485 1095 519 1129
rect 485 1026 519 1060
rect 485 957 519 991
rect 485 888 519 922
rect 485 819 519 853
rect 485 750 519 784
rect 485 681 519 715
rect 485 612 519 646
rect 485 543 519 577
rect 485 474 519 508
rect 485 405 519 439
rect 485 336 519 370
rect 485 267 519 301
rect 485 198 519 232
rect 485 129 519 163
rect 485 60 519 94
<< poly >>
rect 0 2559 98 2575
rect 0 2525 16 2559
rect 50 2525 98 2559
rect 0 2475 98 2525
rect 398 2475 430 2575
rect 891 2584 957 2600
rect 891 2582 907 2584
rect 627 2552 659 2582
rect 859 2552 907 2582
rect 891 2550 907 2552
rect 941 2550 957 2584
rect 891 2516 957 2550
rect 891 2496 907 2516
rect 0 2464 66 2475
rect 0 2430 16 2464
rect 50 2430 66 2464
rect 0 2419 66 2430
rect 627 2466 659 2496
rect 859 2482 907 2496
rect 941 2482 957 2516
rect 859 2466 957 2482
rect 0 2369 98 2419
rect 0 2335 16 2369
rect 50 2335 98 2369
rect 0 2319 98 2335
rect 398 2319 430 2419
rect 627 2380 659 2410
rect 859 2394 957 2410
rect 859 2380 907 2394
rect 891 2360 907 2380
rect 941 2360 957 2394
rect 891 2326 957 2360
rect 891 2324 907 2326
rect 627 2294 659 2324
rect 859 2294 907 2324
rect 891 2292 907 2294
rect 941 2292 957 2326
rect 891 2276 957 2292
rect 627 1863 659 2043
rect 859 2027 957 2043
rect 859 1993 907 2027
rect 941 1993 957 2027
rect 859 1954 957 1993
rect 859 1920 907 1954
rect 941 1920 957 1954
rect 859 1881 957 1920
rect 859 1863 907 1881
rect 891 1847 907 1863
rect 941 1847 957 1881
rect 891 1808 957 1847
rect 891 1807 907 1808
rect 627 1627 659 1807
rect 859 1774 907 1807
rect 941 1774 957 1808
rect 859 1735 957 1774
rect 859 1701 907 1735
rect 941 1701 957 1735
rect 859 1662 957 1701
rect 859 1628 907 1662
rect 941 1628 957 1662
rect 859 1627 957 1628
rect 891 1589 957 1627
rect 891 1555 907 1589
rect 941 1555 957 1589
rect 891 1516 957 1555
rect 891 1482 907 1516
rect 941 1482 957 1516
rect 891 1450 957 1482
rect 627 1270 659 1450
rect 859 1444 957 1450
rect 859 1410 907 1444
rect 941 1410 957 1444
rect 859 1372 957 1410
rect 859 1338 907 1372
rect 941 1338 957 1372
rect 859 1300 957 1338
rect 859 1270 907 1300
rect 891 1266 907 1270
rect 941 1266 957 1300
rect 891 1228 957 1266
rect 891 1214 907 1228
rect 627 1034 659 1214
rect 859 1194 907 1214
rect 941 1194 957 1228
rect 859 1156 957 1194
rect 859 1122 907 1156
rect 941 1122 957 1156
rect 859 1084 957 1122
rect 859 1050 907 1084
rect 941 1050 957 1084
rect 859 1034 957 1050
rect 562 682 594 782
rect 894 766 992 782
rect 894 732 942 766
rect 976 732 992 766
rect 894 682 992 732
rect 926 671 992 682
rect 926 637 942 671
rect 976 637 992 671
rect 926 626 992 637
rect 562 526 594 626
rect 894 576 992 626
rect 894 542 942 576
rect 976 542 992 576
rect 894 526 992 542
rect 5890 551 6031 567
rect 5890 517 5906 551
rect 5940 517 5981 551
rect 6015 517 6031 551
rect 5890 501 6031 517
rect 5911 469 6031 501
rect 6087 551 6228 567
rect 6087 517 6103 551
rect 6137 517 6178 551
rect 6212 517 6228 551
rect 6087 501 6228 517
rect 6087 469 6207 501
rect 562 245 594 345
rect 894 329 992 345
rect 894 295 942 329
rect 976 295 992 329
rect 5911 297 6031 329
rect 6087 297 6207 329
rect 894 245 992 295
rect 926 234 992 245
rect 926 200 942 234
rect 976 200 992 234
rect 926 189 992 200
rect 562 89 594 189
rect 894 139 992 189
rect 894 105 942 139
rect 976 105 992 139
rect 894 89 992 105
<< polycont >>
rect 16 2525 50 2559
rect 907 2550 941 2584
rect 16 2430 50 2464
rect 907 2482 941 2516
rect 16 2335 50 2369
rect 907 2360 941 2394
rect 907 2292 941 2326
rect 907 1993 941 2027
rect 907 1920 941 1954
rect 907 1847 941 1881
rect 907 1774 941 1808
rect 907 1701 941 1735
rect 907 1628 941 1662
rect 907 1555 941 1589
rect 907 1482 941 1516
rect 907 1410 941 1444
rect 907 1338 941 1372
rect 907 1266 941 1300
rect 907 1194 941 1228
rect 907 1122 941 1156
rect 907 1050 941 1084
rect 942 732 976 766
rect 942 637 976 671
rect 942 542 976 576
rect 5906 517 5940 551
rect 5981 517 6015 551
rect 6103 517 6137 551
rect 6178 517 6212 551
rect 942 295 976 329
rect 942 200 976 234
rect 942 105 976 139
<< locali >>
rect 133 2627 857 2651
rect 133 2620 485 2627
rect 132 2586 148 2620
rect 182 2586 216 2620
rect 250 2586 284 2620
rect 318 2586 352 2620
rect 386 2593 485 2620
rect 519 2593 671 2627
rect 705 2593 739 2627
rect 773 2593 807 2627
rect 841 2593 857 2627
rect 386 2586 402 2593
rect 16 2563 50 2575
rect 16 2464 50 2525
rect 485 2559 519 2593
rect 907 2588 941 2600
rect 907 2584 913 2588
rect 941 2550 947 2554
rect 485 2491 519 2525
rect 655 2507 667 2541
rect 705 2507 739 2541
rect 773 2507 807 2541
rect 841 2507 857 2541
rect 907 2516 947 2550
rect 941 2512 947 2516
rect 132 2430 148 2464
rect 182 2430 216 2464
rect 250 2430 284 2464
rect 335 2430 352 2464
rect 907 2478 913 2482
rect 519 2457 857 2467
rect 907 2466 941 2478
rect 485 2455 857 2457
rect 16 2369 50 2430
rect 16 2319 50 2331
rect 485 2423 671 2455
rect 519 2421 671 2423
rect 705 2421 739 2455
rect 773 2421 807 2455
rect 841 2421 857 2455
rect 519 2409 857 2421
rect 485 2357 519 2389
rect 907 2398 941 2410
rect 907 2394 913 2398
rect 793 2369 831 2372
rect 485 2355 489 2357
rect 655 2335 671 2369
rect 705 2335 739 2369
rect 793 2338 807 2369
rect 941 2360 947 2364
rect 773 2335 807 2338
rect 841 2335 857 2338
rect 519 2321 523 2323
rect 132 2274 148 2308
rect 182 2274 216 2308
rect 250 2274 284 2308
rect 318 2274 352 2308
rect 386 2294 402 2308
rect 485 2294 523 2321
rect 907 2326 947 2360
rect 941 2322 947 2326
rect 386 2287 857 2294
rect 386 2274 485 2287
rect 519 2284 857 2287
rect 132 2253 485 2274
rect 523 2283 857 2284
rect 132 2250 489 2253
rect 523 2250 671 2283
rect 132 2249 671 2250
rect 705 2249 739 2283
rect 773 2249 807 2283
rect 841 2249 857 2283
rect 907 2288 913 2292
rect 907 2276 941 2288
rect 132 2236 857 2249
rect 485 2219 523 2236
rect 519 2211 523 2219
rect 485 2177 489 2185
rect 485 2151 523 2177
rect 519 2138 523 2151
rect 485 2104 489 2117
rect 485 2083 523 2104
rect 519 2065 523 2083
rect 655 2054 671 2088
rect 705 2054 739 2088
rect 779 2086 807 2088
rect 773 2054 807 2086
rect 841 2054 857 2088
rect 485 2031 489 2049
rect 485 2015 523 2031
rect 519 1992 523 2015
rect 745 2048 779 2054
rect 907 2031 941 2043
rect 907 2027 913 2031
rect 485 1958 489 1981
rect 485 1947 523 1958
rect 519 1919 523 1947
rect 485 1885 489 1913
rect 941 1993 947 1997
rect 907 1958 947 1993
rect 907 1954 913 1958
rect 941 1920 947 1924
rect 485 1879 523 1885
rect 519 1846 523 1879
rect 485 1812 489 1845
rect 655 1818 671 1852
rect 705 1818 739 1852
rect 773 1818 807 1852
rect 841 1818 871 1852
rect 485 1811 523 1812
rect 519 1777 523 1811
rect 837 1814 871 1818
rect 907 1885 947 1920
rect 907 1881 913 1885
rect 941 1847 947 1851
rect 907 1812 947 1847
rect 907 1808 913 1812
rect 485 1773 523 1777
rect 485 1743 489 1773
rect 519 1709 523 1739
rect 485 1700 523 1709
rect 485 1675 489 1700
rect 941 1774 947 1778
rect 907 1739 947 1774
rect 907 1735 913 1739
rect 941 1701 947 1705
rect 519 1641 523 1666
rect 485 1627 523 1641
rect 485 1607 489 1627
rect 745 1616 779 1636
rect 907 1666 947 1701
rect 907 1662 913 1666
rect 941 1628 947 1632
rect 519 1573 523 1593
rect 655 1582 671 1616
rect 705 1582 739 1616
rect 773 1598 807 1616
rect 779 1582 807 1598
rect 841 1582 857 1616
rect 907 1593 947 1628
rect 907 1589 913 1593
rect 485 1554 523 1573
rect 485 1539 489 1554
rect 941 1555 947 1559
rect 907 1520 947 1555
rect 519 1505 523 1520
rect 485 1481 523 1505
rect 485 1471 489 1481
rect 661 1461 677 1495
rect 711 1461 745 1495
rect 779 1461 813 1495
rect 847 1461 871 1486
rect 519 1437 523 1447
rect 485 1408 523 1437
rect 837 1448 871 1461
rect 907 1516 913 1520
rect 941 1482 947 1486
rect 907 1447 947 1482
rect 907 1444 913 1447
rect 485 1403 489 1408
rect 519 1369 523 1374
rect 485 1335 523 1369
rect 485 1267 523 1301
rect 941 1410 947 1413
rect 907 1374 947 1410
rect 907 1372 913 1374
rect 941 1338 947 1340
rect 907 1301 947 1338
rect 907 1300 913 1301
rect 519 1262 523 1267
rect 663 1259 697 1260
rect 941 1266 947 1267
rect 485 1228 489 1233
rect 485 1198 523 1228
rect 661 1225 677 1259
rect 711 1225 745 1259
rect 779 1225 813 1259
rect 847 1225 863 1259
rect 907 1228 947 1266
rect 519 1189 523 1198
rect 663 1222 697 1225
rect 485 1155 489 1164
rect 485 1129 523 1155
rect 519 1116 523 1129
rect 485 1082 489 1095
rect 907 1156 947 1194
rect 941 1154 947 1156
rect 907 1120 913 1122
rect 485 1060 523 1082
rect 519 1043 523 1060
rect 485 1009 489 1026
rect 837 1023 871 1052
rect 907 1084 947 1120
rect 941 1080 947 1084
rect 907 1046 913 1050
rect 907 1034 941 1046
rect 485 991 523 1009
rect 519 970 523 991
rect 661 989 677 1023
rect 711 989 745 1023
rect 779 989 813 1023
rect 847 1014 871 1023
rect 485 936 489 957
rect 485 922 523 936
rect 519 897 523 922
rect 485 863 489 888
rect 485 853 523 863
rect 519 824 523 853
rect 485 790 489 819
rect 485 784 523 790
rect 519 751 523 784
rect 585 827 619 828
rect 585 793 606 827
rect 640 793 674 827
rect 708 793 742 827
rect 776 793 810 827
rect 844 793 860 827
rect 585 790 619 793
rect 942 770 976 782
rect 942 766 960 770
rect 485 717 489 750
rect 485 715 523 717
rect 519 681 523 715
rect 976 732 994 736
rect 485 678 523 681
rect 485 646 489 678
rect 745 671 779 673
rect 942 671 994 732
rect 519 612 523 644
rect 590 637 606 671
rect 640 637 674 671
rect 708 637 742 671
rect 776 637 810 671
rect 844 637 860 671
rect 485 605 523 612
rect 485 577 489 605
rect 745 635 779 637
rect 519 543 523 571
rect 942 576 994 637
rect 976 572 994 576
rect 485 532 523 543
rect 485 508 489 532
rect 519 474 523 498
rect 485 459 523 474
rect 485 439 489 459
rect 5937 551 5985 557
rect 942 538 960 542
rect 942 526 976 538
rect 5890 523 5903 551
rect 5890 517 5906 523
rect 5940 517 5981 551
rect 6019 523 6031 551
rect 6015 517 6031 523
rect 6087 517 6103 551
rect 6137 550 6178 551
rect 6149 517 6178 550
rect 6212 517 6228 551
rect 585 515 619 517
rect 585 481 606 515
rect 640 481 674 515
rect 708 481 742 515
rect 776 481 810 515
rect 844 481 860 515
rect 585 479 619 481
rect 6115 478 6149 516
rect 5866 461 5900 473
rect 519 405 523 425
rect 485 386 523 405
rect 662 390 696 392
rect 485 370 489 386
rect 590 356 606 390
rect 640 356 674 390
rect 708 356 742 390
rect 776 356 810 390
rect 844 356 860 390
rect 5866 389 5900 423
rect 519 336 523 352
rect 485 313 523 336
rect 662 354 696 356
rect 942 333 976 345
rect 5866 339 5900 351
rect 6042 457 6076 473
rect 6218 461 6252 473
rect 6042 389 6076 423
rect 6042 339 6076 355
rect 6218 389 6252 423
rect 6218 339 6252 351
rect 942 329 960 333
rect 485 301 489 313
rect 519 267 523 279
rect 976 295 994 299
rect 485 239 523 267
rect 485 232 489 239
rect 837 234 871 236
rect 519 198 523 205
rect 590 200 606 234
rect 640 200 674 234
rect 708 200 742 234
rect 776 200 810 234
rect 844 200 871 234
rect 485 165 523 198
rect 485 163 489 165
rect 837 198 871 200
rect 942 234 994 295
rect 942 139 994 200
rect 976 135 994 139
rect 519 129 523 131
rect 485 94 523 129
rect 519 91 523 94
rect 662 78 696 99
rect 942 101 960 105
rect 942 89 976 101
rect 485 57 489 60
rect 485 36 519 57
rect 590 44 606 78
rect 640 61 674 78
rect 640 44 662 61
rect 708 44 742 78
rect 776 44 810 78
rect 844 44 860 78
<< viali >>
rect 16 2559 50 2563
rect 16 2529 50 2559
rect 913 2584 947 2588
rect 913 2554 941 2584
rect 941 2554 947 2584
rect 667 2507 671 2541
rect 671 2507 701 2541
rect 739 2507 773 2541
rect 16 2430 50 2464
rect 301 2430 318 2464
rect 318 2430 335 2464
rect 373 2430 386 2464
rect 386 2430 407 2464
rect 913 2482 941 2512
rect 941 2482 947 2512
rect 913 2478 947 2482
rect 16 2335 50 2365
rect 16 2331 50 2335
rect 913 2394 947 2398
rect 759 2369 793 2372
rect 831 2369 865 2372
rect 489 2355 523 2357
rect 489 2323 519 2355
rect 519 2323 523 2355
rect 759 2338 773 2369
rect 773 2338 793 2369
rect 831 2338 841 2369
rect 841 2338 865 2369
rect 913 2364 941 2394
rect 941 2364 947 2394
rect 489 2253 519 2284
rect 519 2253 523 2284
rect 489 2250 523 2253
rect 913 2292 941 2322
rect 941 2292 947 2322
rect 913 2288 947 2292
rect 489 2185 519 2211
rect 519 2185 523 2211
rect 489 2177 523 2185
rect 489 2117 519 2138
rect 519 2117 523 2138
rect 489 2104 523 2117
rect 745 2088 779 2120
rect 489 2049 519 2065
rect 519 2049 523 2065
rect 745 2086 773 2088
rect 773 2086 779 2088
rect 489 2031 523 2049
rect 745 2014 779 2048
rect 913 2027 947 2031
rect 489 1981 519 1992
rect 519 1981 523 1992
rect 489 1958 523 1981
rect 489 1913 519 1919
rect 519 1913 523 1919
rect 489 1885 523 1913
rect 913 1997 941 2027
rect 941 1997 947 2027
rect 913 1954 947 1958
rect 913 1924 941 1954
rect 941 1924 947 1954
rect 837 1852 871 1886
rect 489 1845 519 1846
rect 519 1845 523 1846
rect 489 1812 523 1845
rect 837 1780 871 1814
rect 913 1881 947 1885
rect 913 1851 941 1881
rect 941 1851 947 1881
rect 913 1808 947 1812
rect 489 1743 523 1773
rect 489 1739 519 1743
rect 519 1739 523 1743
rect 489 1675 523 1700
rect 489 1666 519 1675
rect 519 1666 523 1675
rect 913 1778 941 1808
rect 941 1778 947 1808
rect 913 1735 947 1739
rect 913 1705 941 1735
rect 941 1705 947 1735
rect 489 1607 523 1627
rect 745 1636 779 1670
rect 913 1662 947 1666
rect 913 1632 941 1662
rect 941 1632 947 1662
rect 489 1593 519 1607
rect 519 1593 523 1607
rect 745 1582 773 1598
rect 773 1582 779 1598
rect 913 1589 947 1593
rect 745 1564 779 1582
rect 489 1539 523 1554
rect 489 1520 519 1539
rect 519 1520 523 1539
rect 913 1559 941 1589
rect 941 1559 947 1589
rect 837 1495 871 1520
rect 489 1471 523 1481
rect 489 1447 519 1471
rect 519 1447 523 1471
rect 837 1486 847 1495
rect 847 1486 871 1495
rect 837 1414 871 1448
rect 913 1516 947 1520
rect 913 1486 941 1516
rect 941 1486 947 1516
rect 913 1444 947 1447
rect 489 1403 523 1408
rect 489 1374 519 1403
rect 519 1374 523 1403
rect 489 1301 519 1335
rect 519 1301 523 1335
rect 913 1413 941 1444
rect 941 1413 947 1444
rect 913 1372 947 1374
rect 913 1340 941 1372
rect 941 1340 947 1372
rect 913 1300 947 1301
rect 489 1233 519 1262
rect 519 1233 523 1262
rect 663 1260 697 1294
rect 913 1267 941 1300
rect 941 1267 947 1300
rect 489 1228 523 1233
rect 489 1164 519 1189
rect 519 1164 523 1189
rect 663 1188 697 1222
rect 913 1194 941 1228
rect 941 1194 947 1228
rect 489 1155 523 1164
rect 489 1095 519 1116
rect 519 1095 523 1116
rect 489 1082 523 1095
rect 913 1122 941 1154
rect 941 1122 947 1154
rect 913 1120 947 1122
rect 489 1026 519 1043
rect 519 1026 523 1043
rect 489 1009 523 1026
rect 837 1052 871 1086
rect 913 1050 941 1080
rect 941 1050 947 1080
rect 913 1046 947 1050
rect 837 989 847 1014
rect 847 989 871 1014
rect 837 980 871 989
rect 489 957 519 970
rect 519 957 523 970
rect 489 936 523 957
rect 489 888 519 897
rect 519 888 523 897
rect 489 863 523 888
rect 489 819 519 824
rect 519 819 523 824
rect 489 790 523 819
rect 585 828 619 862
rect 585 756 619 790
rect 960 766 994 770
rect 489 750 519 751
rect 519 750 523 751
rect 489 717 523 750
rect 960 736 976 766
rect 976 736 994 766
rect 489 646 523 678
rect 745 673 779 707
rect 489 644 519 646
rect 519 644 523 646
rect 960 637 976 671
rect 976 637 994 671
rect 489 577 523 605
rect 745 601 779 635
rect 489 571 519 577
rect 519 571 523 577
rect 489 508 523 532
rect 489 498 519 508
rect 519 498 523 508
rect 489 439 523 459
rect 585 517 619 551
rect 960 542 976 572
rect 976 542 994 572
rect 5903 551 5937 557
rect 5985 551 6019 557
rect 960 538 994 542
rect 5903 523 5906 551
rect 5906 523 5937 551
rect 5985 523 6015 551
rect 6015 523 6019 551
rect 6115 517 6137 550
rect 6137 517 6149 550
rect 6115 516 6149 517
rect 585 445 619 479
rect 5866 457 5900 461
rect 489 425 519 439
rect 519 425 523 439
rect 5866 427 5900 457
rect 662 392 696 426
rect 489 370 523 386
rect 489 352 519 370
rect 519 352 523 370
rect 662 320 696 354
rect 5866 355 5900 385
rect 5866 351 5900 355
rect 6115 444 6149 478
rect 6218 457 6252 461
rect 6218 427 6252 457
rect 6218 355 6252 385
rect 6218 351 6252 355
rect 960 329 994 333
rect 489 301 523 313
rect 489 279 519 301
rect 519 279 523 301
rect 960 299 976 329
rect 976 299 994 329
rect 489 232 523 239
rect 837 236 871 270
rect 489 205 519 232
rect 519 205 523 232
rect 489 163 523 165
rect 837 164 871 198
rect 960 200 976 234
rect 976 200 994 234
rect 489 131 519 163
rect 519 131 523 163
rect 489 60 519 91
rect 519 60 523 91
rect 662 99 696 133
rect 960 105 976 135
rect 976 105 994 135
rect 960 101 994 105
rect 489 57 523 60
rect 662 44 674 61
rect 674 44 696 61
rect 662 27 696 44
<< metal1 >>
rect 907 2588 953 2600
rect 10 2563 56 2575
rect 10 2529 16 2563
rect 50 2529 56 2563
rect 907 2554 913 2588
rect 947 2554 953 2588
rect 10 2464 56 2529
rect 655 2541 785 2547
rect 655 2507 667 2541
rect 701 2507 739 2541
rect 773 2507 785 2541
rect 655 2501 785 2507
rect 907 2512 953 2554
rect 10 2430 16 2464
rect 50 2430 56 2464
rect 10 2365 56 2430
rect 289 2464 625 2470
rect 289 2430 301 2464
rect 335 2430 373 2464
rect 407 2430 625 2464
rect 289 2424 625 2430
tri 554 2399 579 2424 ne
rect 10 2331 16 2365
rect 50 2331 56 2365
rect 10 2319 56 2331
rect 483 2357 529 2369
rect 483 2323 489 2357
rect 523 2323 529 2357
rect 483 2284 529 2323
rect 483 2250 489 2284
rect 523 2250 529 2284
rect 483 2211 529 2250
rect 483 2177 489 2211
rect 523 2177 529 2211
rect 483 2138 529 2177
rect 483 2104 489 2138
rect 523 2104 529 2138
rect 483 2065 529 2104
rect 483 2031 489 2065
rect 523 2031 529 2065
rect 483 1992 529 2031
rect 483 1958 489 1992
rect 523 1958 529 1992
rect 483 1919 529 1958
rect 483 1885 489 1919
rect 523 1885 529 1919
rect 483 1846 529 1885
rect 483 1812 489 1846
rect 523 1812 529 1846
rect 483 1773 529 1812
rect 483 1739 489 1773
rect 523 1739 529 1773
rect 483 1700 529 1739
rect 483 1666 489 1700
rect 523 1666 529 1700
rect 483 1627 529 1666
rect 483 1593 489 1627
rect 523 1593 529 1627
rect 483 1554 529 1593
rect 483 1520 489 1554
rect 523 1520 529 1554
rect 483 1481 529 1520
rect 483 1447 489 1481
rect 523 1447 529 1481
rect 483 1408 529 1447
rect 483 1374 489 1408
rect 523 1374 529 1408
rect 483 1335 529 1374
rect 483 1301 489 1335
rect 523 1301 529 1335
rect 483 1262 529 1301
rect 483 1228 489 1262
rect 523 1228 529 1262
rect 483 1189 529 1228
rect 483 1155 489 1189
rect 523 1155 529 1189
rect 483 1116 529 1155
rect 483 1082 489 1116
rect 523 1082 529 1116
rect 483 1043 529 1082
rect 579 1077 625 2424
rect 657 1294 703 2501
rect 907 2478 913 2512
rect 947 2478 953 2512
rect 907 2466 953 2478
rect 907 2398 953 2410
rect 747 2372 877 2378
rect 747 2338 759 2372
rect 793 2338 831 2372
rect 865 2338 877 2372
rect 747 2332 877 2338
rect 657 1260 663 1294
rect 697 1260 703 1294
rect 657 1222 703 1260
rect 657 1188 663 1222
rect 697 1188 703 1222
rect 657 1176 703 1188
rect 739 2120 785 2132
rect 739 2086 745 2120
rect 779 2086 785 2120
rect 739 2048 785 2086
rect 739 2014 745 2048
rect 779 2014 785 2048
rect 739 1670 785 2014
rect 831 1886 877 2332
rect 907 2364 913 2398
rect 947 2364 953 2398
rect 907 2322 953 2364
rect 907 2288 913 2322
rect 947 2288 953 2322
rect 907 2276 953 2288
rect 831 1852 837 1886
rect 871 1852 877 1886
rect 831 1814 877 1852
rect 831 1780 837 1814
rect 871 1780 877 1814
rect 831 1768 877 1780
rect 907 2031 953 2043
rect 907 1997 913 2031
rect 947 1997 953 2031
rect 907 1958 953 1997
rect 907 1924 913 1958
rect 947 1924 953 1958
rect 907 1885 953 1924
rect 907 1851 913 1885
rect 947 1851 953 1885
rect 907 1812 953 1851
rect 907 1778 913 1812
rect 947 1778 953 1812
rect 739 1636 745 1670
rect 779 1636 785 1670
rect 739 1598 785 1636
rect 739 1564 745 1598
rect 779 1564 785 1598
rect 483 1009 489 1043
rect 523 1009 529 1043
rect 483 970 529 1009
rect 483 936 489 970
rect 523 936 529 970
rect 573 1071 625 1077
rect 573 1007 625 1019
rect 573 949 625 955
rect 483 897 529 936
rect 483 863 489 897
rect 523 863 529 897
rect 483 824 529 863
rect 483 790 489 824
rect 523 790 529 824
rect 483 751 529 790
rect 483 717 489 751
rect 523 717 529 751
rect 483 678 529 717
rect 483 644 489 678
rect 523 644 529 678
rect 483 605 529 644
rect 483 571 489 605
rect 523 571 529 605
rect 483 532 529 571
rect 483 498 489 532
rect 523 498 529 532
rect 483 459 529 498
rect 483 425 489 459
rect 523 425 529 459
rect 483 386 529 425
rect 483 352 489 386
rect 523 352 529 386
rect 483 313 529 352
rect 483 279 489 313
rect 523 279 529 313
rect 483 239 529 279
rect 483 205 489 239
rect 523 205 529 239
rect 483 165 529 205
rect 483 131 489 165
rect 523 131 529 165
rect 579 862 625 949
rect 579 828 585 862
rect 619 828 625 862
rect 579 790 625 828
rect 579 756 585 790
rect 619 756 625 790
rect 579 551 625 756
rect 579 517 585 551
rect 619 517 625 551
rect 579 479 625 517
rect 579 445 585 479
rect 619 445 625 479
rect 579 136 625 445
rect 656 1014 702 1083
rect 656 1008 708 1014
rect 656 944 708 956
rect 656 886 708 892
rect 656 426 702 886
rect 739 707 785 1564
rect 907 1739 953 1778
rect 907 1705 913 1739
rect 947 1705 953 1739
rect 907 1666 953 1705
rect 907 1632 913 1666
rect 947 1632 953 1666
rect 907 1593 953 1632
rect 907 1559 913 1593
rect 947 1559 953 1593
rect 739 673 745 707
rect 779 673 785 707
rect 739 635 785 673
rect 739 601 745 635
rect 779 601 785 635
rect 739 589 785 601
rect 831 1520 877 1532
rect 831 1486 837 1520
rect 871 1486 877 1520
rect 831 1448 877 1486
rect 831 1414 837 1448
rect 871 1414 877 1448
rect 831 1086 877 1414
rect 831 1052 837 1086
rect 871 1052 877 1086
rect 831 1014 877 1052
rect 907 1520 953 1559
rect 907 1486 913 1520
rect 947 1486 953 1520
rect 907 1447 953 1486
rect 907 1413 913 1447
rect 947 1413 953 1447
rect 907 1374 953 1413
rect 907 1340 913 1374
rect 947 1340 953 1374
rect 907 1301 953 1340
rect 907 1267 913 1301
rect 947 1267 953 1301
rect 907 1228 953 1267
rect 907 1194 913 1228
rect 947 1194 953 1228
rect 907 1154 953 1194
rect 907 1120 913 1154
rect 947 1120 953 1154
rect 907 1080 953 1120
rect 907 1046 913 1080
rect 947 1046 953 1080
rect 907 1034 953 1046
rect 831 980 837 1014
rect 871 980 877 1014
rect 656 392 662 426
rect 696 392 702 426
rect 656 354 702 392
rect 656 320 662 354
rect 696 320 702 354
rect 483 91 529 131
rect 483 57 489 91
rect 523 57 529 91
rect 483 45 529 57
rect 656 133 702 320
rect 831 270 877 980
rect 5734 906 5740 958
rect 5792 906 5804 958
rect 5856 906 5862 958
tri 5777 885 5798 906 ne
rect 5798 885 5841 906
tri 5841 885 5862 906 nw
rect 5912 906 5918 958
rect 5970 906 5982 958
rect 6034 906 6040 958
rect 6163 906 6169 958
rect 6221 906 6233 958
rect 6285 906 6291 958
tri 5912 885 5933 906 ne
rect 5933 885 5976 906
tri 5976 885 5997 906 nw
tri 6188 885 6209 906 ne
rect 6209 885 6258 906
tri 5798 882 5801 885 ne
rect 831 236 837 270
rect 871 236 877 270
rect 831 198 877 236
rect 831 164 837 198
rect 871 164 877 198
rect 831 152 877 164
rect 954 770 1000 782
rect 954 736 960 770
rect 994 736 1000 770
rect 954 671 1000 736
rect 954 637 960 671
rect 994 637 1000 671
rect 954 572 1000 637
rect 954 538 960 572
rect 994 538 1000 572
rect 954 333 1000 538
rect 5801 478 5841 885
tri 5933 882 5936 885 ne
tri 5914 563 5936 585 se
rect 5936 563 5976 885
tri 6209 882 6212 885 ne
tri 5976 563 5998 585 sw
rect 5891 557 6031 563
rect 5891 523 5903 557
rect 5937 523 5985 557
rect 6019 523 6031 557
rect 5891 517 6031 523
rect 6109 550 6155 562
rect 6109 516 6115 550
rect 6149 516 6155 550
tri 6101 492 6109 500 se
rect 6109 492 6155 516
tri 5841 478 5855 492 sw
tri 6087 478 6101 492 se
rect 6101 478 6155 492
rect 5801 473 5855 478
tri 5855 473 5860 478 sw
tri 6082 473 6087 478 se
rect 6087 473 6115 478
rect 5801 461 6115 473
rect 5801 427 5866 461
rect 5900 444 6115 461
rect 6149 473 6155 478
rect 6149 444 6156 473
rect 5900 432 6156 444
rect 6212 461 6258 885
tri 6258 883 6281 906 nw
rect 5900 427 5927 432
tri 5927 427 5932 432 nw
rect 6212 427 6218 461
rect 6252 427 6258 461
rect 5801 385 5906 427
tri 5906 406 5927 427 nw
rect 5801 351 5866 385
rect 5900 351 5906 385
rect 5801 339 5906 351
rect 6212 385 6258 427
rect 6212 351 6218 385
rect 6252 351 6258 385
rect 6212 339 6258 351
rect 954 299 960 333
rect 994 299 1000 333
rect 954 234 1000 299
rect 954 200 960 234
rect 994 200 1000 234
rect 656 99 662 133
rect 696 99 702 133
rect 656 61 702 99
rect 954 135 1000 200
rect 954 101 960 135
rect 994 101 1000 135
rect 954 89 1000 101
rect 656 27 662 61
rect 696 27 702 61
rect 656 15 702 27
<< via1 >>
rect 573 1019 625 1071
rect 573 955 625 1007
rect 656 956 708 1008
rect 656 892 708 944
rect 5740 906 5792 958
rect 5804 906 5856 958
rect 5918 906 5970 958
rect 5982 906 6034 958
rect 6169 906 6221 958
rect 6233 906 6285 958
<< metal2 >>
rect 573 1071 4987 1077
rect 625 1050 4987 1071
tri 4987 1050 5014 1077 sw
rect 625 1043 6186 1050
rect 573 1007 625 1019
tri 4946 1014 4975 1043 ne
rect 4975 1014 6186 1043
tri 6186 1014 6222 1050 sw
rect 573 949 625 955
rect 656 1008 4918 1014
rect 708 994 4918 1008
tri 4918 994 4938 1014 sw
tri 4975 994 4995 1014 ne
rect 4995 994 6222 1014
rect 708 982 4938 994
tri 2026 962 2046 982 ne
rect 2046 962 2174 982
tri 2174 962 2194 982 nw
tri 4861 962 4881 982 ne
rect 4881 962 4938 982
tri 4938 962 4970 994 sw
tri 5889 971 5912 994 ne
rect 5912 963 6222 994
tri 6222 963 6273 1014 sw
tri 4881 958 4885 962 ne
rect 4885 958 5862 962
rect 656 944 708 956
tri 4885 925 4918 958 ne
rect 4918 925 5740 958
tri 4918 906 4937 925 ne
rect 4937 906 5740 925
rect 5792 906 5804 958
rect 5856 906 5862 958
rect 5912 958 6291 963
rect 5912 906 5918 958
rect 5970 906 5982 958
rect 6034 906 6169 958
rect 6221 906 6233 958
rect 6285 906 6291 958
rect 656 886 708 892
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1666464484
transform 0 -1 859 1 0 1034
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1666464484
transform 0 1 659 1 0 1627
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808502  sky130_fd_pr__nfet_01v8__example_55959141808502_0
timestamp 1666464484
transform 0 1 659 1 0 2294
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_0
timestamp 1666464484
transform 0 -1 398 -1 0 2575
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_1
timestamp 1666464484
transform 0 1 594 1 0 526
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_2
timestamp 1666464484
transform 0 1 594 1 0 89
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808500  sky130_fd_pr__pfet_01v8__example_55959141808500_0
timestamp 1666464484
transform -1 0 6207 0 -1 469
box -1 0 297 1
<< labels >>
flabel comment s 964 998 964 998 0 FreeSans 400 0 0 0 NET248
flabel comment s 924 2347 924 2347 0 FreeSans 400 90 0 0 IN_H
<< properties >>
string GDS_END 29636908
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29617420
<< end >>
