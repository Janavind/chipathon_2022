magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 7 21 1309 203
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 177
rect 277 47 307 177
rect 361 47 391 177
rect 445 47 475 177
rect 529 47 559 177
rect 613 47 643 177
rect 697 47 727 177
rect 781 47 811 177
rect 865 47 895 177
rect 949 47 979 177
rect 1033 47 1063 177
rect 1117 47 1147 177
rect 1201 47 1231 177
<< scpmoshvt >>
rect 89 297 119 497
rect 173 297 203 497
rect 257 297 287 497
rect 341 297 371 497
rect 425 297 455 497
rect 613 297 643 497
rect 697 297 727 497
rect 781 297 811 497
rect 865 297 895 497
rect 949 297 979 497
rect 1033 297 1063 497
rect 1117 297 1147 497
rect 1201 297 1231 497
<< ndiff >>
rect 33 163 89 177
rect 33 129 45 163
rect 79 129 89 163
rect 33 95 89 129
rect 33 61 45 95
rect 79 61 89 95
rect 33 47 89 61
rect 119 163 171 177
rect 119 129 129 163
rect 163 129 171 163
rect 119 95 171 129
rect 119 61 129 95
rect 163 61 171 95
rect 119 47 171 61
rect 225 95 277 177
rect 225 61 233 95
rect 267 61 277 95
rect 225 47 277 61
rect 307 163 361 177
rect 307 129 317 163
rect 351 129 361 163
rect 307 47 361 129
rect 391 95 445 177
rect 391 61 401 95
rect 435 61 445 95
rect 391 47 445 61
rect 475 163 529 177
rect 475 129 485 163
rect 519 129 529 163
rect 475 47 529 129
rect 559 163 613 177
rect 559 129 569 163
rect 603 129 613 163
rect 559 95 613 129
rect 559 61 569 95
rect 603 61 613 95
rect 559 47 613 61
rect 643 95 697 177
rect 643 61 653 95
rect 687 61 697 95
rect 643 47 697 61
rect 727 163 781 177
rect 727 129 737 163
rect 771 129 781 163
rect 727 95 781 129
rect 727 61 737 95
rect 771 61 781 95
rect 727 47 781 61
rect 811 95 865 177
rect 811 61 821 95
rect 855 61 865 95
rect 811 47 865 61
rect 895 163 949 177
rect 895 129 905 163
rect 939 129 949 163
rect 895 95 949 129
rect 895 61 905 95
rect 939 61 949 95
rect 895 47 949 61
rect 979 95 1033 177
rect 979 61 989 95
rect 1023 61 1033 95
rect 979 47 1033 61
rect 1063 163 1117 177
rect 1063 129 1073 163
rect 1107 129 1117 163
rect 1063 95 1117 129
rect 1063 61 1073 95
rect 1107 61 1117 95
rect 1063 47 1117 61
rect 1147 95 1201 177
rect 1147 61 1157 95
rect 1191 61 1201 95
rect 1147 47 1201 61
rect 1231 163 1283 177
rect 1231 129 1241 163
rect 1275 129 1283 163
rect 1231 95 1283 129
rect 1231 61 1241 95
rect 1275 61 1283 95
rect 1231 47 1283 61
<< pdiff >>
rect 33 477 89 497
rect 33 443 45 477
rect 79 443 89 477
rect 33 409 89 443
rect 33 375 45 409
rect 79 375 89 409
rect 33 341 89 375
rect 33 307 45 341
rect 79 307 89 341
rect 33 297 89 307
rect 119 477 173 497
rect 119 443 129 477
rect 163 443 173 477
rect 119 409 173 443
rect 119 375 129 409
rect 163 375 173 409
rect 119 297 173 375
rect 203 477 257 497
rect 203 443 213 477
rect 247 443 257 477
rect 203 409 257 443
rect 203 375 213 409
rect 247 375 257 409
rect 203 341 257 375
rect 203 307 213 341
rect 247 307 257 341
rect 203 297 257 307
rect 287 477 341 497
rect 287 443 297 477
rect 331 443 341 477
rect 287 409 341 443
rect 287 375 297 409
rect 331 375 341 409
rect 287 297 341 375
rect 371 477 425 497
rect 371 443 381 477
rect 415 443 425 477
rect 371 409 425 443
rect 371 375 381 409
rect 415 375 425 409
rect 371 341 425 375
rect 371 307 381 341
rect 415 307 425 341
rect 371 297 425 307
rect 455 477 507 497
rect 455 443 465 477
rect 499 443 507 477
rect 455 409 507 443
rect 455 375 465 409
rect 499 375 507 409
rect 455 297 507 375
rect 561 477 613 497
rect 561 443 569 477
rect 603 443 613 477
rect 561 409 613 443
rect 561 375 569 409
rect 603 375 613 409
rect 561 297 613 375
rect 643 409 697 497
rect 643 375 653 409
rect 687 375 697 409
rect 643 341 697 375
rect 643 307 653 341
rect 687 307 697 341
rect 643 297 697 307
rect 727 477 781 497
rect 727 443 737 477
rect 771 443 781 477
rect 727 409 781 443
rect 727 375 737 409
rect 771 375 781 409
rect 727 297 781 375
rect 811 409 865 497
rect 811 375 821 409
rect 855 375 865 409
rect 811 341 865 375
rect 811 307 821 341
rect 855 307 865 341
rect 811 297 865 307
rect 895 477 949 497
rect 895 443 905 477
rect 939 443 949 477
rect 895 409 949 443
rect 895 375 905 409
rect 939 375 949 409
rect 895 341 949 375
rect 895 307 905 341
rect 939 307 949 341
rect 895 297 949 307
rect 979 477 1033 497
rect 979 443 989 477
rect 1023 443 1033 477
rect 979 409 1033 443
rect 979 375 989 409
rect 1023 375 1033 409
rect 979 297 1033 375
rect 1063 477 1117 497
rect 1063 443 1073 477
rect 1107 443 1117 477
rect 1063 409 1117 443
rect 1063 375 1073 409
rect 1107 375 1117 409
rect 1063 341 1117 375
rect 1063 307 1073 341
rect 1107 307 1117 341
rect 1063 297 1117 307
rect 1147 477 1201 497
rect 1147 443 1157 477
rect 1191 443 1201 477
rect 1147 409 1201 443
rect 1147 375 1157 409
rect 1191 375 1201 409
rect 1147 297 1201 375
rect 1231 477 1287 497
rect 1231 443 1241 477
rect 1275 443 1287 477
rect 1231 409 1287 443
rect 1231 375 1241 409
rect 1275 375 1287 409
rect 1231 341 1287 375
rect 1231 307 1241 341
rect 1275 307 1287 341
rect 1231 297 1287 307
<< ndiffc >>
rect 45 129 79 163
rect 45 61 79 95
rect 129 129 163 163
rect 129 61 163 95
rect 233 61 267 95
rect 317 129 351 163
rect 401 61 435 95
rect 485 129 519 163
rect 569 129 603 163
rect 569 61 603 95
rect 653 61 687 95
rect 737 129 771 163
rect 737 61 771 95
rect 821 61 855 95
rect 905 129 939 163
rect 905 61 939 95
rect 989 61 1023 95
rect 1073 129 1107 163
rect 1073 61 1107 95
rect 1157 61 1191 95
rect 1241 129 1275 163
rect 1241 61 1275 95
<< pdiffc >>
rect 45 443 79 477
rect 45 375 79 409
rect 45 307 79 341
rect 129 443 163 477
rect 129 375 163 409
rect 213 443 247 477
rect 213 375 247 409
rect 213 307 247 341
rect 297 443 331 477
rect 297 375 331 409
rect 381 443 415 477
rect 381 375 415 409
rect 381 307 415 341
rect 465 443 499 477
rect 465 375 499 409
rect 569 443 603 477
rect 569 375 603 409
rect 653 375 687 409
rect 653 307 687 341
rect 737 443 771 477
rect 737 375 771 409
rect 821 375 855 409
rect 821 307 855 341
rect 905 443 939 477
rect 905 375 939 409
rect 905 307 939 341
rect 989 443 1023 477
rect 989 375 1023 409
rect 1073 443 1107 477
rect 1073 375 1107 409
rect 1073 307 1107 341
rect 1157 443 1191 477
rect 1157 375 1191 409
rect 1241 443 1275 477
rect 1241 375 1275 409
rect 1241 307 1275 341
<< poly >>
rect 89 497 119 523
rect 173 497 203 523
rect 257 497 287 523
rect 341 497 371 523
rect 425 497 455 523
rect 613 497 643 523
rect 697 497 727 523
rect 781 497 811 523
rect 865 497 895 523
rect 949 497 979 523
rect 1033 497 1063 523
rect 1117 497 1147 523
rect 1201 497 1231 523
rect 89 265 119 297
rect 42 249 119 265
rect 42 215 61 249
rect 95 215 119 249
rect 42 199 119 215
rect 173 265 203 297
rect 257 265 287 297
rect 341 265 371 297
rect 425 265 455 297
rect 613 265 643 297
rect 697 265 727 297
rect 781 265 811 297
rect 865 265 895 297
rect 173 249 559 265
rect 173 215 189 249
rect 223 215 257 249
rect 291 215 325 249
rect 359 215 393 249
rect 427 215 559 249
rect 173 199 559 215
rect 89 177 119 199
rect 277 177 307 199
rect 361 177 391 199
rect 445 177 475 199
rect 529 177 559 199
rect 613 249 895 265
rect 613 215 629 249
rect 663 215 697 249
rect 731 215 765 249
rect 799 215 833 249
rect 867 215 895 249
rect 613 199 895 215
rect 613 177 643 199
rect 697 177 727 199
rect 781 177 811 199
rect 865 177 895 199
rect 949 265 979 297
rect 1033 265 1063 297
rect 1117 265 1147 297
rect 1201 265 1231 297
rect 949 249 1231 265
rect 949 215 959 249
rect 993 215 1027 249
rect 1061 215 1095 249
rect 1129 215 1163 249
rect 1197 215 1231 249
rect 949 199 1231 215
rect 949 177 979 199
rect 1033 177 1063 199
rect 1117 177 1147 199
rect 1201 177 1231 199
rect 89 21 119 47
rect 277 21 307 47
rect 361 21 391 47
rect 445 21 475 47
rect 529 21 559 47
rect 613 21 643 47
rect 697 21 727 47
rect 781 21 811 47
rect 865 21 895 47
rect 949 21 979 47
rect 1033 21 1063 47
rect 1117 21 1147 47
rect 1201 21 1231 47
<< polycont >>
rect 61 215 95 249
rect 189 215 223 249
rect 257 215 291 249
rect 325 215 359 249
rect 393 215 427 249
rect 629 215 663 249
rect 697 215 731 249
rect 765 215 799 249
rect 833 215 867 249
rect 959 215 993 249
rect 1027 215 1061 249
rect 1095 215 1129 249
rect 1163 215 1197 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 29 477 95 487
rect 29 443 45 477
rect 79 443 95 477
rect 29 409 95 443
rect 29 375 45 409
rect 79 375 95 409
rect 29 341 95 375
rect 129 477 171 527
rect 163 443 171 477
rect 129 409 171 443
rect 163 375 171 409
rect 129 359 171 375
rect 213 477 255 493
rect 247 443 255 477
rect 213 409 255 443
rect 247 375 255 409
rect 29 307 45 341
rect 79 325 95 341
rect 213 341 255 375
rect 289 477 339 527
rect 289 443 297 477
rect 331 443 339 477
rect 289 409 339 443
rect 289 375 297 409
rect 331 375 339 409
rect 289 359 339 375
rect 373 477 423 493
rect 373 443 381 477
rect 415 443 423 477
rect 373 409 423 443
rect 373 375 381 409
rect 415 375 423 409
rect 79 307 179 325
rect 29 291 179 307
rect 247 325 255 341
rect 373 341 423 375
rect 457 477 507 527
rect 457 443 465 477
rect 499 443 507 477
rect 457 409 507 443
rect 457 375 465 409
rect 499 375 507 409
rect 457 359 507 375
rect 555 477 947 493
rect 555 443 569 477
rect 603 459 737 477
rect 603 443 611 459
rect 555 409 611 443
rect 729 443 737 459
rect 771 459 905 477
rect 771 443 779 459
rect 555 375 569 409
rect 603 375 611 409
rect 555 359 611 375
rect 645 409 695 425
rect 645 375 653 409
rect 687 375 695 409
rect 373 325 381 341
rect 247 307 381 325
rect 415 325 423 341
rect 645 341 695 375
rect 729 409 779 443
rect 897 443 905 459
rect 939 443 947 477
rect 729 375 737 409
rect 771 375 779 409
rect 729 359 779 375
rect 813 409 863 425
rect 813 375 821 409
rect 855 375 863 409
rect 645 325 653 341
rect 415 307 653 325
rect 687 325 695 341
rect 813 341 863 375
rect 813 325 821 341
rect 687 307 821 325
rect 855 307 863 341
rect 213 291 863 307
rect 897 409 947 443
rect 897 375 905 409
rect 939 375 947 409
rect 897 341 947 375
rect 981 477 1031 527
rect 981 443 989 477
rect 1023 443 1031 477
rect 981 409 1031 443
rect 981 375 989 409
rect 1023 375 1031 409
rect 981 359 1031 375
rect 1065 477 1115 493
rect 1065 443 1073 477
rect 1107 443 1115 477
rect 1065 409 1115 443
rect 1065 375 1073 409
rect 1107 375 1115 409
rect 897 307 905 341
rect 939 325 947 341
rect 1065 341 1115 375
rect 1149 477 1199 527
rect 1149 443 1157 477
rect 1191 443 1199 477
rect 1149 409 1199 443
rect 1149 375 1157 409
rect 1191 375 1199 409
rect 1149 359 1199 375
rect 1233 477 1283 493
rect 1233 443 1241 477
rect 1275 443 1283 477
rect 1233 409 1283 443
rect 1233 375 1241 409
rect 1275 375 1283 409
rect 1065 325 1073 341
rect 939 307 1073 325
rect 1107 325 1115 341
rect 1233 341 1283 375
rect 1233 325 1241 341
rect 1107 307 1241 325
rect 1275 307 1283 341
rect 897 291 1283 307
rect 145 257 179 291
rect 489 289 863 291
rect 17 249 111 257
rect 17 215 61 249
rect 95 215 111 249
rect 145 249 455 257
rect 145 215 189 249
rect 223 215 257 249
rect 291 215 325 249
rect 359 215 393 249
rect 427 215 455 249
rect 489 215 579 289
rect 1317 257 1362 491
rect 613 249 895 255
rect 613 215 629 249
rect 663 215 697 249
rect 731 215 765 249
rect 799 215 833 249
rect 867 215 895 249
rect 929 249 1362 257
rect 929 215 959 249
rect 993 215 1027 249
rect 1061 215 1095 249
rect 1129 215 1163 249
rect 1197 215 1362 249
rect 145 179 179 215
rect 45 163 79 179
rect 45 95 79 129
rect 45 17 79 61
rect 113 163 179 179
rect 489 163 535 215
rect 113 129 129 163
rect 163 129 179 163
rect 284 129 317 163
rect 351 129 485 163
rect 519 129 535 163
rect 569 163 1291 181
rect 603 145 737 163
rect 603 129 619 145
rect 113 95 179 129
rect 569 95 619 129
rect 721 129 737 145
rect 771 145 905 163
rect 771 129 787 145
rect 113 61 129 95
rect 163 61 179 95
rect 216 61 233 95
rect 267 61 401 95
rect 435 61 569 95
rect 603 61 619 95
rect 653 95 687 111
rect 113 58 179 61
rect 653 17 687 61
rect 721 95 787 129
rect 889 129 905 145
rect 939 145 1073 163
rect 939 129 955 145
rect 721 61 737 95
rect 771 61 787 95
rect 721 51 787 61
rect 821 95 855 111
rect 821 17 855 61
rect 889 95 955 129
rect 1057 129 1073 145
rect 1107 145 1241 163
rect 1107 129 1123 145
rect 889 61 905 95
rect 939 61 955 95
rect 889 51 955 61
rect 989 95 1023 111
rect 989 17 1023 61
rect 1057 95 1123 129
rect 1225 129 1241 145
rect 1275 129 1291 163
rect 1057 61 1073 95
rect 1107 61 1123 95
rect 1057 51 1123 61
rect 1157 95 1191 111
rect 1157 17 1191 61
rect 1225 95 1291 129
rect 1225 61 1241 95
rect 1275 61 1291 95
rect 1225 51 1291 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 489 289 523 323 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o21bai_4
rlabel metal1 s 0 -48 1380 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 1352826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1342018
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 6.900 2.720 
<< end >>
