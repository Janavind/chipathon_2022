magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< pwell >>
rect 10 10 634 392
<< nmoslvt >>
rect 92 36 122 366
rect 178 36 208 366
rect 264 36 294 366
rect 350 36 380 366
rect 436 36 466 366
rect 522 36 552 366
<< ndiff >>
rect 36 329 92 366
rect 36 295 47 329
rect 81 295 92 329
rect 36 257 92 295
rect 36 223 47 257
rect 81 223 92 257
rect 36 185 92 223
rect 36 151 47 185
rect 81 151 92 185
rect 36 113 92 151
rect 36 79 47 113
rect 81 79 92 113
rect 36 36 92 79
rect 122 329 178 366
rect 122 295 133 329
rect 167 295 178 329
rect 122 257 178 295
rect 122 223 133 257
rect 167 223 178 257
rect 122 185 178 223
rect 122 151 133 185
rect 167 151 178 185
rect 122 113 178 151
rect 122 79 133 113
rect 167 79 178 113
rect 122 36 178 79
rect 208 329 264 366
rect 208 295 219 329
rect 253 295 264 329
rect 208 257 264 295
rect 208 223 219 257
rect 253 223 264 257
rect 208 185 264 223
rect 208 151 219 185
rect 253 151 264 185
rect 208 113 264 151
rect 208 79 219 113
rect 253 79 264 113
rect 208 36 264 79
rect 294 329 350 366
rect 294 295 305 329
rect 339 295 350 329
rect 294 257 350 295
rect 294 223 305 257
rect 339 223 350 257
rect 294 185 350 223
rect 294 151 305 185
rect 339 151 350 185
rect 294 113 350 151
rect 294 79 305 113
rect 339 79 350 113
rect 294 36 350 79
rect 380 329 436 366
rect 380 295 391 329
rect 425 295 436 329
rect 380 257 436 295
rect 380 223 391 257
rect 425 223 436 257
rect 380 185 436 223
rect 380 151 391 185
rect 425 151 436 185
rect 380 113 436 151
rect 380 79 391 113
rect 425 79 436 113
rect 380 36 436 79
rect 466 329 522 366
rect 466 295 477 329
rect 511 295 522 329
rect 466 257 522 295
rect 466 223 477 257
rect 511 223 522 257
rect 466 185 522 223
rect 466 151 477 185
rect 511 151 522 185
rect 466 113 522 151
rect 466 79 477 113
rect 511 79 522 113
rect 466 36 522 79
rect 552 329 608 366
rect 552 295 563 329
rect 597 295 608 329
rect 552 257 608 295
rect 552 223 563 257
rect 597 223 608 257
rect 552 185 608 223
rect 552 151 563 185
rect 597 151 608 185
rect 552 113 608 151
rect 552 79 563 113
rect 597 79 608 113
rect 552 36 608 79
<< ndiffc >>
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 305 295 339 329
rect 305 223 339 257
rect 305 151 339 185
rect 305 79 339 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
rect 477 295 511 329
rect 477 223 511 257
rect 477 151 511 185
rect 477 79 511 113
rect 563 295 597 329
rect 563 223 597 257
rect 563 151 597 185
rect 563 79 597 113
<< poly >>
rect 92 447 552 463
rect 92 413 135 447
rect 169 413 203 447
rect 237 413 271 447
rect 305 413 339 447
rect 373 413 407 447
rect 441 413 475 447
rect 509 413 552 447
rect 92 392 552 413
rect 92 366 122 392
rect 178 366 208 392
rect 264 366 294 392
rect 350 366 380 392
rect 436 366 466 392
rect 522 366 552 392
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
<< polycont >>
rect 135 413 169 447
rect 203 413 237 447
rect 271 413 305 447
rect 339 413 373 447
rect 407 413 441 447
rect 475 413 509 447
<< locali >>
rect 119 447 525 463
rect 119 413 125 447
rect 169 413 197 447
rect 237 413 269 447
rect 305 413 339 447
rect 375 413 407 447
rect 447 413 475 447
rect 519 413 525 447
rect 119 397 525 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 329 167 357
rect 133 257 167 295
rect 133 185 167 223
rect 133 113 167 151
rect 133 51 167 79
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
rect 305 329 339 357
rect 305 257 339 295
rect 305 185 339 223
rect 305 113 339 151
rect 305 51 339 79
rect 391 329 425 357
rect 391 257 425 295
rect 391 185 425 223
rect 391 113 425 151
rect 391 51 425 79
rect 477 329 511 357
rect 477 257 511 295
rect 477 185 511 223
rect 477 113 511 151
rect 477 51 511 79
rect 563 329 597 357
rect 563 257 597 295
rect 563 185 597 223
rect 563 113 597 151
rect 563 51 597 79
<< viali >>
rect 125 413 135 447
rect 135 413 159 447
rect 197 413 203 447
rect 203 413 231 447
rect 269 413 271 447
rect 271 413 303 447
rect 341 413 373 447
rect 373 413 375 447
rect 413 413 441 447
rect 441 413 447 447
rect 485 413 509 447
rect 509 413 519 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 305 295 339 329
rect 305 223 339 257
rect 305 151 339 185
rect 305 79 339 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
rect 477 295 511 329
rect 477 223 511 257
rect 477 151 511 185
rect 477 79 511 113
rect 563 295 597 329
rect 563 223 597 257
rect 563 151 597 185
rect 563 79 597 113
<< metal1 >>
rect 113 447 531 459
rect 113 413 125 447
rect 159 413 197 447
rect 231 413 269 447
rect 303 413 341 447
rect 375 413 413 447
rect 447 413 485 447
rect 519 413 531 447
rect 113 401 531 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 124 338 176 357
rect 124 274 176 286
rect 124 185 176 222
rect 124 151 133 185
rect 167 151 176 185
rect 124 113 176 151
rect 124 79 133 113
rect 167 79 176 113
rect 124 51 176 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 296 338 348 357
rect 296 274 348 286
rect 296 185 348 222
rect 296 151 305 185
rect 339 151 348 185
rect 296 113 348 151
rect 296 79 305 113
rect 339 79 348 113
rect 296 51 348 79
rect 385 329 431 357
rect 385 295 391 329
rect 425 295 431 329
rect 385 257 431 295
rect 385 223 391 257
rect 425 223 431 257
rect 385 185 431 223
rect 385 151 391 185
rect 425 151 431 185
rect 385 113 431 151
rect 385 79 391 113
rect 425 79 431 113
rect 385 -29 431 79
rect 468 338 520 357
rect 468 274 520 286
rect 468 185 520 222
rect 468 151 477 185
rect 511 151 520 185
rect 468 113 520 151
rect 468 79 477 113
rect 511 79 520 113
rect 468 51 520 79
rect 557 329 603 357
rect 557 295 563 329
rect 597 295 603 329
rect 557 257 603 295
rect 557 223 563 257
rect 597 223 603 257
rect 557 185 603 223
rect 557 151 563 185
rect 597 151 603 185
rect 557 113 603 151
rect 557 79 563 113
rect 597 79 603 113
rect 557 -29 603 79
rect 41 -89 603 -29
<< via1 >>
rect 124 329 176 338
rect 124 295 133 329
rect 133 295 167 329
rect 167 295 176 329
rect 124 286 176 295
rect 124 257 176 274
rect 124 223 133 257
rect 133 223 167 257
rect 167 223 176 257
rect 124 222 176 223
rect 296 329 348 338
rect 296 295 305 329
rect 305 295 339 329
rect 339 295 348 329
rect 296 286 348 295
rect 296 257 348 274
rect 296 223 305 257
rect 305 223 339 257
rect 339 223 348 257
rect 296 222 348 223
rect 468 329 520 338
rect 468 295 477 329
rect 477 295 511 329
rect 511 295 520 329
rect 468 286 520 295
rect 468 257 520 274
rect 468 223 477 257
rect 477 223 511 257
rect 511 223 520 257
rect 468 222 520 223
<< metal2 >>
rect 117 348 183 357
rect 117 292 122 348
rect 178 292 183 348
rect 117 286 124 292
rect 176 286 183 292
rect 117 274 183 286
rect 117 268 124 274
rect 176 268 183 274
rect 117 212 122 268
rect 178 212 183 268
rect 117 203 183 212
rect 289 348 355 357
rect 289 292 294 348
rect 350 292 355 348
rect 289 286 296 292
rect 348 286 355 292
rect 289 274 355 286
rect 289 268 296 274
rect 348 268 355 274
rect 289 212 294 268
rect 350 212 355 268
rect 289 203 355 212
rect 461 348 527 357
rect 461 292 466 348
rect 522 292 527 348
rect 461 286 468 292
rect 520 286 527 292
rect 461 274 527 286
rect 461 268 468 274
rect 520 268 527 274
rect 461 212 466 268
rect 522 212 527 268
rect 461 203 527 212
<< via2 >>
rect 122 338 178 348
rect 122 292 124 338
rect 124 292 176 338
rect 176 292 178 338
rect 122 222 124 268
rect 124 222 176 268
rect 176 222 178 268
rect 122 212 178 222
rect 294 338 350 348
rect 294 292 296 338
rect 296 292 348 338
rect 348 292 350 338
rect 294 222 296 268
rect 296 222 348 268
rect 348 222 350 268
rect 294 212 350 222
rect 466 338 522 348
rect 466 292 468 338
rect 468 292 520 338
rect 520 292 522 338
rect 466 222 468 268
rect 468 222 520 268
rect 520 222 522 268
rect 466 212 522 222
<< metal3 >>
rect 117 348 527 357
rect 117 292 122 348
rect 178 292 294 348
rect 350 292 466 348
rect 522 292 527 348
rect 117 291 527 292
rect 117 268 183 291
rect 117 212 122 268
rect 178 212 183 268
rect 117 203 183 212
rect 289 268 355 291
rect 289 212 294 268
rect 350 212 355 268
rect 289 203 355 212
rect 461 268 527 291
rect 461 212 466 268
rect 522 212 527 268
rect 461 203 527 212
<< labels >>
flabel metal3 s 117 291 527 357 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 113 401 531 459 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 -89 603 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel pwell s 79 370 89 387 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 3302400
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3291330
string path 1.025 -1.475 15.075 -1.475 
<< end >>
