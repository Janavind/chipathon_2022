magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_0
timestamp 1666464484
transform 1 0 30 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_1
timestamp 1666464484
transform 1 0 116 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_2
timestamp 1666464484
transform 1 0 202 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808251  sky130_fd_pr__hvdfm1sd2__example_55959141808251_3
timestamp 1666464484
transform 1 0 288 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808250  sky130_fd_pr__hvdfm1sd__example_55959141808250_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808250  sky130_fd_pr__hvdfm1sd__example_55959141808250_1
timestamp 1666464484
transform 1 0 374 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 32722654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32719656
<< end >>
