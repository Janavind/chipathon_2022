magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 24 21 1256 203
rect 25 -17 59 21
<< locali >>
rect 136 333 179 493
rect 313 333 350 493
rect 17 292 350 333
rect 17 177 147 292
rect 556 271 630 339
rect 936 306 1271 340
rect 936 272 994 306
rect 556 211 715 271
rect 753 211 819 272
rect 853 211 994 272
rect 1028 211 1094 272
rect 1128 211 1271 306
rect 17 143 353 177
rect 136 131 353 143
rect 136 51 179 131
rect 313 51 353 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 367 102 527
rect 213 367 279 527
rect 384 292 450 527
rect 488 414 522 493
rect 556 448 622 527
rect 752 414 818 493
rect 488 374 818 414
rect 488 258 522 374
rect 852 340 902 493
rect 936 414 970 493
rect 1004 448 1070 527
rect 1104 414 1144 493
rect 936 374 1144 414
rect 1178 374 1271 493
rect 181 211 522 258
rect 664 306 902 340
rect 488 177 522 211
rect 17 17 102 109
rect 213 17 279 97
rect 387 17 450 177
rect 488 127 642 177
rect 676 127 1271 177
rect 676 93 714 127
rect 488 51 714 93
rect 752 17 818 89
rect 852 51 886 127
rect 920 17 986 89
rect 1020 51 1054 127
rect 1088 17 1154 89
rect 1188 51 1271 127
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< obsm1 >>
rect 845 456 903 465
rect 1213 456 1271 465
rect 845 428 1271 456
rect 845 419 903 428
rect 1213 419 1271 428
<< labels >>
rlabel locali s 1028 211 1094 272 6 A1
port 1 nsew signal input
rlabel locali s 1128 211 1271 306 6 A2
port 2 nsew signal input
rlabel locali s 853 211 994 272 6 A2
port 2 nsew signal input
rlabel locali s 936 272 994 306 6 A2
port 2 nsew signal input
rlabel locali s 936 306 1271 340 6 A2
port 2 nsew signal input
rlabel locali s 753 211 819 272 6 A3
port 3 nsew signal input
rlabel locali s 556 211 715 271 6 B1
port 4 nsew signal input
rlabel locali s 556 271 630 339 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 25 -17 59 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 24 21 1256 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 313 51 353 131 6 X
port 9 nsew signal output
rlabel locali s 136 51 179 131 6 X
port 9 nsew signal output
rlabel locali s 136 131 353 143 6 X
port 9 nsew signal output
rlabel locali s 17 143 353 177 6 X
port 9 nsew signal output
rlabel locali s 17 177 147 292 6 X
port 9 nsew signal output
rlabel locali s 17 292 350 333 6 X
port 9 nsew signal output
rlabel locali s 313 333 350 493 6 X
port 9 nsew signal output
rlabel locali s 136 333 179 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1288 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1423826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1412714
<< end >>
