magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -85 800 809 1568
<< pwell >>
rect 189 76 769 728
<< mvnmos >>
rect 268 102 388 702
rect 444 102 564 702
<< mvpmos >>
rect 126 866 246 1466
rect 302 866 422 1466
rect 478 866 598 1466
<< mvndiff >>
rect 215 624 268 702
rect 215 590 223 624
rect 257 590 268 624
rect 215 556 268 590
rect 215 522 223 556
rect 257 522 268 556
rect 215 488 268 522
rect 215 454 223 488
rect 257 454 268 488
rect 215 420 268 454
rect 215 386 223 420
rect 257 386 268 420
rect 215 352 268 386
rect 215 318 223 352
rect 257 318 268 352
rect 215 284 268 318
rect 215 250 223 284
rect 257 250 268 284
rect 215 216 268 250
rect 215 182 223 216
rect 257 182 268 216
rect 215 148 268 182
rect 215 114 223 148
rect 257 114 268 148
rect 215 102 268 114
rect 388 624 444 702
rect 388 590 399 624
rect 433 590 444 624
rect 388 556 444 590
rect 388 522 399 556
rect 433 522 444 556
rect 388 488 444 522
rect 388 454 399 488
rect 433 454 444 488
rect 388 420 444 454
rect 388 386 399 420
rect 433 386 444 420
rect 388 352 444 386
rect 388 318 399 352
rect 433 318 444 352
rect 388 284 444 318
rect 388 250 399 284
rect 433 250 444 284
rect 388 216 444 250
rect 388 182 399 216
rect 433 182 444 216
rect 388 148 444 182
rect 388 114 399 148
rect 433 114 444 148
rect 388 102 444 114
rect 564 624 617 702
rect 564 590 575 624
rect 609 590 617 624
rect 564 556 617 590
rect 564 522 575 556
rect 609 522 617 556
rect 564 488 617 522
rect 564 454 575 488
rect 609 454 617 488
rect 564 420 617 454
rect 564 386 575 420
rect 609 386 617 420
rect 564 352 617 386
rect 564 318 575 352
rect 609 318 617 352
rect 564 284 617 318
rect 564 250 575 284
rect 609 250 617 284
rect 564 216 617 250
rect 564 182 575 216
rect 609 182 617 216
rect 564 148 617 182
rect 564 114 575 148
rect 609 114 617 148
rect 564 102 617 114
<< mvpdiff >>
rect 73 1454 126 1466
rect 73 1420 81 1454
rect 115 1420 126 1454
rect 73 1386 126 1420
rect 73 1352 81 1386
rect 115 1352 126 1386
rect 73 1318 126 1352
rect 73 1284 81 1318
rect 115 1284 126 1318
rect 73 1250 126 1284
rect 73 1216 81 1250
rect 115 1216 126 1250
rect 73 1182 126 1216
rect 73 1148 81 1182
rect 115 1148 126 1182
rect 73 1114 126 1148
rect 73 1080 81 1114
rect 115 1080 126 1114
rect 73 1046 126 1080
rect 73 1012 81 1046
rect 115 1012 126 1046
rect 73 978 126 1012
rect 73 944 81 978
rect 115 944 126 978
rect 73 866 126 944
rect 246 1454 302 1466
rect 246 1420 257 1454
rect 291 1420 302 1454
rect 246 1386 302 1420
rect 246 1352 257 1386
rect 291 1352 302 1386
rect 246 1318 302 1352
rect 246 1284 257 1318
rect 291 1284 302 1318
rect 246 1250 302 1284
rect 246 1216 257 1250
rect 291 1216 302 1250
rect 246 1182 302 1216
rect 246 1148 257 1182
rect 291 1148 302 1182
rect 246 1114 302 1148
rect 246 1080 257 1114
rect 291 1080 302 1114
rect 246 1046 302 1080
rect 246 1012 257 1046
rect 291 1012 302 1046
rect 246 978 302 1012
rect 246 944 257 978
rect 291 944 302 978
rect 246 866 302 944
rect 422 1454 478 1466
rect 422 1420 433 1454
rect 467 1420 478 1454
rect 422 1386 478 1420
rect 422 1352 433 1386
rect 467 1352 478 1386
rect 422 1318 478 1352
rect 422 1284 433 1318
rect 467 1284 478 1318
rect 422 1250 478 1284
rect 422 1216 433 1250
rect 467 1216 478 1250
rect 422 1182 478 1216
rect 422 1148 433 1182
rect 467 1148 478 1182
rect 422 1114 478 1148
rect 422 1080 433 1114
rect 467 1080 478 1114
rect 422 1046 478 1080
rect 422 1012 433 1046
rect 467 1012 478 1046
rect 422 978 478 1012
rect 422 944 433 978
rect 467 944 478 978
rect 422 866 478 944
rect 598 1454 651 1466
rect 598 1420 609 1454
rect 643 1420 651 1454
rect 598 1386 651 1420
rect 598 1352 609 1386
rect 643 1352 651 1386
rect 598 1318 651 1352
rect 598 1284 609 1318
rect 643 1284 651 1318
rect 598 1250 651 1284
rect 598 1216 609 1250
rect 643 1216 651 1250
rect 598 1182 651 1216
rect 598 1148 609 1182
rect 643 1148 651 1182
rect 598 1114 651 1148
rect 598 1080 609 1114
rect 643 1080 651 1114
rect 598 1046 651 1080
rect 598 1012 609 1046
rect 643 1012 651 1046
rect 598 978 651 1012
rect 598 944 609 978
rect 643 944 651 978
rect 598 866 651 944
<< mvndiffc >>
rect 223 590 257 624
rect 223 522 257 556
rect 223 454 257 488
rect 223 386 257 420
rect 223 318 257 352
rect 223 250 257 284
rect 223 182 257 216
rect 223 114 257 148
rect 399 590 433 624
rect 399 522 433 556
rect 399 454 433 488
rect 399 386 433 420
rect 399 318 433 352
rect 399 250 433 284
rect 399 182 433 216
rect 399 114 433 148
rect 575 590 609 624
rect 575 522 609 556
rect 575 454 609 488
rect 575 386 609 420
rect 575 318 609 352
rect 575 250 609 284
rect 575 182 609 216
rect 575 114 609 148
<< mvpdiffc >>
rect 81 1420 115 1454
rect 81 1352 115 1386
rect 81 1284 115 1318
rect 81 1216 115 1250
rect 81 1148 115 1182
rect 81 1080 115 1114
rect 81 1012 115 1046
rect 81 944 115 978
rect 257 1420 291 1454
rect 257 1352 291 1386
rect 257 1284 291 1318
rect 257 1216 291 1250
rect 257 1148 291 1182
rect 257 1080 291 1114
rect 257 1012 291 1046
rect 257 944 291 978
rect 433 1420 467 1454
rect 433 1352 467 1386
rect 433 1284 467 1318
rect 433 1216 467 1250
rect 433 1148 467 1182
rect 433 1080 467 1114
rect 433 1012 467 1046
rect 433 944 467 978
rect 609 1420 643 1454
rect 609 1352 643 1386
rect 609 1284 643 1318
rect 609 1216 643 1250
rect 609 1148 643 1182
rect 609 1080 643 1114
rect 609 1012 643 1046
rect 609 944 643 978
<< mvpsubdiff >>
rect 705 665 743 702
rect 705 631 707 665
rect 741 631 743 665
rect 705 597 743 631
rect 705 563 707 597
rect 741 563 743 597
rect 705 529 743 563
rect 705 495 707 529
rect 741 495 743 529
rect 705 461 743 495
rect 705 427 707 461
rect 741 427 743 461
rect 705 393 743 427
rect 705 359 707 393
rect 741 359 743 393
rect 705 325 743 359
rect 705 291 707 325
rect 741 291 743 325
rect 705 257 743 291
rect 705 223 707 257
rect 741 223 743 257
rect 705 189 743 223
rect 705 155 707 189
rect 741 155 743 189
rect 705 102 743 155
<< mvnsubdiff >>
rect -19 1413 19 1462
rect -19 1379 -17 1413
rect 17 1379 19 1413
rect -19 1345 19 1379
rect -19 1311 -17 1345
rect 17 1311 19 1345
rect -19 1277 19 1311
rect -19 1243 -17 1277
rect 17 1243 19 1277
rect -19 1209 19 1243
rect -19 1175 -17 1209
rect 17 1175 19 1209
rect -19 1134 19 1175
rect -19 1100 -17 1134
rect 17 1100 19 1134
rect -19 1066 19 1100
rect -19 1032 -17 1066
rect 17 1032 19 1066
rect -19 998 19 1032
rect -19 964 -17 998
rect 17 964 19 998
rect -19 930 19 964
rect -19 896 -17 930
rect 17 896 19 930
rect -19 866 19 896
rect 705 1413 743 1462
rect 705 1379 707 1413
rect 741 1379 743 1413
rect 705 1345 743 1379
rect 705 1311 707 1345
rect 741 1311 743 1345
rect 705 1277 743 1311
rect 705 1243 707 1277
rect 741 1243 743 1277
rect 705 1209 743 1243
rect 705 1175 707 1209
rect 741 1175 743 1209
rect 705 1134 743 1175
rect 705 1100 707 1134
rect 741 1100 743 1134
rect 705 1066 743 1100
rect 705 1032 707 1066
rect 741 1032 743 1066
rect 705 998 743 1032
rect 705 964 707 998
rect 741 964 743 998
rect 705 930 743 964
rect 705 896 707 930
rect 741 896 743 930
rect 705 866 743 896
<< mvpsubdiffcont >>
rect 707 631 741 665
rect 707 563 741 597
rect 707 495 741 529
rect 707 427 741 461
rect 707 359 741 393
rect 707 291 741 325
rect 707 223 741 257
rect 707 155 741 189
<< mvnsubdiffcont >>
rect -17 1379 17 1413
rect -17 1311 17 1345
rect -17 1243 17 1277
rect -17 1175 17 1209
rect -17 1100 17 1134
rect -17 1032 17 1066
rect -17 964 17 998
rect -17 896 17 930
rect 707 1379 741 1413
rect 707 1311 741 1345
rect 707 1243 741 1277
rect 707 1175 741 1209
rect 707 1100 741 1134
rect 707 1032 741 1066
rect 707 964 741 998
rect 707 896 741 930
<< poly >>
rect 126 1548 422 1568
rect 126 1514 155 1548
rect 189 1514 223 1548
rect 257 1514 291 1548
rect 325 1514 359 1548
rect 393 1514 422 1548
rect 126 1492 422 1514
rect 126 1466 246 1492
rect 302 1466 422 1492
rect 478 1466 598 1492
rect 126 840 246 866
rect 302 840 422 866
rect 478 840 598 866
rect 126 793 388 840
rect 126 759 146 793
rect 180 759 214 793
rect 248 759 282 793
rect 316 759 388 793
rect 126 728 388 759
rect 478 783 634 840
rect 478 749 512 783
rect 546 749 580 783
rect 614 749 634 783
rect 478 728 634 749
rect 268 702 388 728
rect 444 702 564 728
rect 268 76 388 102
rect 246 58 388 76
rect 246 24 266 58
rect 300 24 334 58
rect 368 24 388 58
rect 246 8 388 24
rect 444 76 564 102
rect 444 58 588 76
rect 444 24 466 58
rect 500 24 534 58
rect 568 24 588 58
rect 444 8 588 24
<< polycont >>
rect 155 1514 189 1548
rect 223 1514 257 1548
rect 291 1514 325 1548
rect 359 1514 393 1548
rect 146 759 180 793
rect 214 759 248 793
rect 282 759 316 793
rect 512 749 546 783
rect 580 749 614 783
rect 266 24 300 58
rect 334 24 368 58
rect 466 24 500 58
rect 534 24 568 58
<< locali >>
rect 139 1514 155 1548
rect 189 1514 223 1548
rect 257 1514 291 1548
rect 325 1514 359 1548
rect 393 1514 409 1548
rect 81 1454 115 1470
rect -17 1413 17 1454
rect -17 1345 17 1379
rect -17 1277 17 1311
rect -17 1209 17 1243
rect -17 1134 17 1175
rect -17 1090 17 1100
rect -17 1018 17 1032
rect -17 946 17 964
rect 81 1386 115 1420
rect 81 1318 115 1352
rect 81 1250 115 1284
rect 81 1182 115 1216
rect 257 1454 291 1470
rect 257 1386 291 1420
rect 257 1318 291 1352
rect 257 1250 291 1284
rect 257 1182 291 1216
rect 81 1114 115 1148
rect 149 1144 187 1178
rect 433 1454 467 1470
rect 433 1386 467 1420
rect 609 1454 643 1470
rect 609 1386 643 1420
rect 433 1318 467 1352
rect 571 1340 609 1374
rect 433 1250 467 1284
rect 433 1182 467 1216
rect 81 1046 115 1080
rect 81 978 115 1012
rect 81 928 115 944
rect 257 1114 291 1148
rect 361 1144 399 1178
rect 257 1046 291 1056
rect 257 978 291 984
rect 433 1114 467 1148
rect 433 1046 467 1080
rect 433 978 467 1012
rect 433 928 467 944
rect 609 1318 643 1340
rect 609 1250 643 1284
rect 609 1182 643 1216
rect 609 1114 643 1148
rect 609 1046 643 1080
rect 609 978 643 1012
rect -17 874 17 896
rect 609 880 643 944
rect 399 846 643 880
rect 707 1413 741 1454
rect 707 1345 741 1379
rect 707 1277 741 1311
rect 707 1209 741 1243
rect 707 1134 741 1175
rect 707 1090 741 1100
rect 707 1018 741 1032
rect 707 946 741 964
rect 707 874 741 896
rect 130 759 146 793
rect 180 759 214 793
rect 248 759 282 793
rect 316 759 332 793
rect 223 624 257 640
rect 223 576 257 590
rect 223 504 257 522
rect 223 432 257 454
rect 223 352 257 386
rect 223 284 257 318
rect 223 216 257 250
rect 223 148 257 182
rect 223 98 257 114
rect 399 624 433 846
rect 496 749 512 783
rect 546 749 580 783
rect 614 749 630 783
rect 707 665 741 694
rect 399 556 433 590
rect 399 488 433 522
rect 399 420 433 454
rect 399 352 433 386
rect 399 284 433 318
rect 399 216 433 250
rect 399 148 433 182
rect 399 98 433 114
rect 575 624 609 640
rect 575 576 609 590
rect 575 504 609 522
rect 575 432 609 454
rect 575 352 609 386
rect 575 284 609 318
rect 575 216 609 250
rect 575 148 609 182
rect 575 98 609 114
rect 707 597 741 631
rect 707 529 741 536
rect 707 461 741 464
rect 707 426 741 427
rect 707 325 741 359
rect 707 257 741 291
rect 707 189 741 223
rect 707 110 741 155
rect 250 24 266 58
rect 300 24 334 58
rect 368 24 384 58
rect 450 24 466 58
rect 500 24 534 58
rect 568 24 584 58
<< viali >>
rect -17 1066 17 1090
rect -17 1056 17 1066
rect -17 998 17 1018
rect -17 984 17 998
rect -17 930 17 946
rect -17 912 17 930
rect 115 1144 149 1178
rect 187 1144 221 1178
rect 537 1340 571 1374
rect 609 1352 643 1374
rect 609 1340 643 1352
rect 327 1144 361 1178
rect 399 1144 433 1178
rect 257 1080 291 1090
rect 257 1056 291 1080
rect 257 1012 291 1018
rect 257 984 291 1012
rect 257 944 291 946
rect 257 912 291 944
rect 707 1066 741 1090
rect 707 1056 741 1066
rect 707 998 741 1018
rect 707 984 741 998
rect 707 930 741 946
rect 707 912 741 930
rect 223 556 257 576
rect 223 542 257 556
rect 223 488 257 504
rect 223 470 257 488
rect 223 420 257 432
rect 223 398 257 420
rect 575 556 609 576
rect 575 542 609 556
rect 575 488 609 504
rect 575 470 609 488
rect 575 420 609 432
rect 575 398 609 420
rect 707 563 741 570
rect 707 536 741 563
rect 707 495 741 498
rect 707 464 741 495
rect 707 393 741 426
rect 707 392 741 393
<< metal1 >>
rect 525 1374 655 1380
rect 525 1340 537 1374
rect 571 1340 609 1374
rect 643 1340 655 1374
rect 525 1334 655 1340
rect 103 1178 445 1184
rect 103 1144 115 1178
rect 149 1144 187 1178
rect 221 1144 327 1178
rect 361 1144 399 1178
rect 433 1144 445 1178
rect 103 1138 445 1144
rect -29 1090 753 1108
rect -29 1056 -17 1090
rect 17 1056 257 1090
rect 291 1056 707 1090
rect 741 1056 753 1090
rect -29 1018 753 1056
rect -29 984 -17 1018
rect 17 984 257 1018
rect 291 984 707 1018
rect 741 984 753 1018
rect -29 946 753 984
rect -29 912 -17 946
rect 17 912 257 946
rect 291 912 707 946
rect 741 912 753 946
rect -29 906 753 912
rect 0 576 753 582
rect 0 542 223 576
rect 257 542 575 576
rect 609 570 753 576
rect 609 542 707 570
rect 0 536 707 542
rect 741 536 753 570
rect 0 504 753 536
rect 0 470 223 504
rect 257 470 575 504
rect 609 498 753 504
rect 609 470 707 498
rect 0 464 707 470
rect 741 464 753 498
rect 0 432 753 464
rect 0 398 223 432
rect 257 398 575 432
rect 609 426 753 432
rect 609 398 707 426
rect 0 392 707 398
rect 741 392 753 426
rect 0 380 753 392
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_0
timestamp 1666464484
transform 1 0 268 0 1 102
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_1
timestamp 1666464484
transform -1 0 564 0 1 102
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808365  sky130_fd_pr__pfet_01v8__example_55959141808365_0
timestamp 1666464484
transform 1 0 478 0 -1 1466
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808366  sky130_fd_pr__pfet_01v8__example_55959141808366_0
timestamp 1666464484
transform 1 0 126 0 -1 1466
box -1 0 297 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1666464484
transform 1 0 537 0 1 1340
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1666464484
transform -1 0 433 0 1 1144
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1666464484
transform -1 0 221 0 1 1144
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1666464484
transform -1 0 741 0 1 392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1666464484
transform -1 0 741 0 1 912
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_2
timestamp 1666464484
transform 1 0 -17 0 1 912
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_3
timestamp 1666464484
transform 1 0 257 0 1 912
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_4
timestamp 1666464484
transform 1 0 575 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_5
timestamp 1666464484
transform 1 0 223 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1666464484
transform 0 1 496 1 0 733
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1666464484
transform 0 -1 384 1 0 8
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1666464484
transform 0 -1 584 1 0 8
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1666464484
transform 0 1 130 1 0 743
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1666464484
transform 0 1 139 1 0 1498
box 0 0 1 1
<< labels >>
flabel locali s 496 749 530 783 2 FreeSans 300 0 0 0 DRVLO_H_N
port 1 nsew
flabel locali s 294 759 331 793 6 FreeSans 300 0 0 0 PDEN_H_N
port 2 nsew
flabel metal1 s 0 380 42 582 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 711 380 753 582 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s -29 906 13 1108 6 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 711 906 753 1108 6 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 607 1350 607 1350 7 FreeSans 300 180 0 0 PD_H
port 5 nsew
flabel comment s 334 1166 334 1166 0 FreeSans 200 0 0 0 INT
<< properties >>
string GDS_END 32375178
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32369550
<< end >>
