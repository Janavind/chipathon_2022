magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 0 0 604 1214
<< pmoslvt >>
rect 204 102 274 1112
rect 330 102 400 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 274 1100 330 1112
rect 274 1066 285 1100
rect 319 1066 330 1100
rect 274 1032 330 1066
rect 274 998 285 1032
rect 319 998 330 1032
rect 274 964 330 998
rect 274 930 285 964
rect 319 930 330 964
rect 274 896 330 930
rect 274 862 285 896
rect 319 862 330 896
rect 274 828 330 862
rect 274 794 285 828
rect 319 794 330 828
rect 274 760 330 794
rect 274 726 285 760
rect 319 726 330 760
rect 274 692 330 726
rect 274 658 285 692
rect 319 658 330 692
rect 274 624 330 658
rect 274 590 285 624
rect 319 590 330 624
rect 274 556 330 590
rect 274 522 285 556
rect 319 522 330 556
rect 274 488 330 522
rect 274 454 285 488
rect 319 454 330 488
rect 274 420 330 454
rect 274 386 285 420
rect 319 386 330 420
rect 274 352 330 386
rect 274 318 285 352
rect 319 318 330 352
rect 274 284 330 318
rect 274 250 285 284
rect 319 250 330 284
rect 274 216 330 250
rect 274 182 285 216
rect 319 182 330 216
rect 274 148 330 182
rect 274 114 285 148
rect 319 114 330 148
rect 274 102 330 114
rect 400 1100 456 1112
rect 400 1066 411 1100
rect 445 1066 456 1100
rect 400 1032 456 1066
rect 400 998 411 1032
rect 445 998 456 1032
rect 400 964 456 998
rect 400 930 411 964
rect 445 930 456 964
rect 400 896 456 930
rect 400 862 411 896
rect 445 862 456 896
rect 400 828 456 862
rect 400 794 411 828
rect 445 794 456 828
rect 400 760 456 794
rect 400 726 411 760
rect 445 726 456 760
rect 400 692 456 726
rect 400 658 411 692
rect 445 658 456 692
rect 400 624 456 658
rect 400 590 411 624
rect 445 590 456 624
rect 400 556 456 590
rect 400 522 411 556
rect 445 522 456 556
rect 400 488 456 522
rect 400 454 411 488
rect 445 454 456 488
rect 400 420 456 454
rect 400 386 411 420
rect 445 386 456 420
rect 400 352 456 386
rect 400 318 411 352
rect 445 318 456 352
rect 400 284 456 318
rect 400 250 411 284
rect 445 250 456 284
rect 400 216 456 250
rect 400 182 411 216
rect 445 182 456 216
rect 400 148 456 182
rect 400 114 411 148
rect 445 114 456 148
rect 400 102 456 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 285 1066 319 1100
rect 285 998 319 1032
rect 285 930 319 964
rect 285 862 319 896
rect 285 794 319 828
rect 285 726 319 760
rect 285 658 319 692
rect 285 590 319 624
rect 285 522 319 556
rect 285 454 319 488
rect 285 386 319 420
rect 285 318 319 352
rect 285 250 319 284
rect 285 182 319 216
rect 285 114 319 148
rect 411 1066 445 1100
rect 411 998 445 1032
rect 411 930 445 964
rect 411 862 445 896
rect 411 794 445 828
rect 411 726 445 760
rect 411 658 445 692
rect 411 590 445 624
rect 411 522 445 556
rect 411 454 445 488
rect 411 386 445 420
rect 411 318 445 352
rect 411 250 445 284
rect 411 182 445 216
rect 411 114 445 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 510 1066 568 1112
rect 510 1032 522 1066
rect 556 1032 568 1066
rect 510 998 568 1032
rect 510 964 522 998
rect 556 964 568 998
rect 510 930 568 964
rect 510 896 522 930
rect 556 896 568 930
rect 510 862 568 896
rect 510 828 522 862
rect 556 828 568 862
rect 510 794 568 828
rect 510 760 522 794
rect 556 760 568 794
rect 510 726 568 760
rect 510 692 522 726
rect 556 692 568 726
rect 510 658 568 692
rect 510 624 522 658
rect 556 624 568 658
rect 510 590 568 624
rect 510 556 522 590
rect 556 556 568 590
rect 510 522 568 556
rect 510 488 522 522
rect 556 488 568 522
rect 510 454 568 488
rect 510 420 522 454
rect 556 420 568 454
rect 510 386 568 420
rect 510 352 522 386
rect 556 352 568 386
rect 510 318 568 352
rect 510 284 522 318
rect 556 284 568 318
rect 510 250 568 284
rect 510 216 522 250
rect 556 216 568 250
rect 510 182 568 216
rect 510 148 522 182
rect 556 148 568 182
rect 510 102 568 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 522 1032 556 1066
rect 522 964 556 998
rect 522 896 556 930
rect 522 828 556 862
rect 522 760 556 794
rect 522 692 556 726
rect 522 624 556 658
rect 522 556 556 590
rect 522 488 556 522
rect 522 420 556 454
rect 522 352 556 386
rect 522 284 556 318
rect 522 216 556 250
rect 522 148 556 182
<< poly >>
rect 165 1194 439 1214
rect 165 1160 183 1194
rect 217 1160 251 1194
rect 285 1160 319 1194
rect 353 1160 387 1194
rect 421 1160 439 1194
rect 165 1144 439 1160
rect 204 1112 274 1144
rect 330 1112 400 1144
rect 204 70 274 102
rect 330 70 400 102
rect 165 54 439 70
rect 165 20 183 54
rect 217 20 251 54
rect 285 20 319 54
rect 353 20 387 54
rect 421 20 439 54
rect 165 0 439 20
<< polycont >>
rect 183 1160 217 1194
rect 251 1160 285 1194
rect 319 1160 353 1194
rect 387 1160 421 1194
rect 183 20 217 54
rect 251 20 285 54
rect 319 20 353 54
rect 387 20 421 54
<< locali >>
rect 165 1160 177 1194
rect 217 1160 249 1194
rect 285 1160 319 1194
rect 355 1160 387 1194
rect 427 1160 439 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 285 1100 319 1116
rect 285 1032 319 1058
rect 285 964 319 986
rect 285 896 319 914
rect 285 828 319 842
rect 285 760 319 770
rect 285 692 319 698
rect 285 624 319 626
rect 285 588 319 590
rect 285 516 319 522
rect 285 444 319 454
rect 285 372 319 386
rect 285 300 319 318
rect 285 228 319 250
rect 285 156 319 182
rect 285 98 319 114
rect 411 1100 445 1116
rect 411 1032 445 1058
rect 411 964 445 986
rect 411 896 445 914
rect 411 828 445 842
rect 411 760 445 770
rect 411 692 445 698
rect 411 624 445 626
rect 411 588 445 590
rect 411 516 445 522
rect 411 444 445 454
rect 411 372 445 386
rect 411 300 445 318
rect 411 228 445 250
rect 411 156 445 182
rect 522 1020 556 1032
rect 522 948 556 964
rect 522 876 556 896
rect 522 804 556 828
rect 522 732 556 760
rect 522 660 556 692
rect 522 590 556 624
rect 522 522 556 554
rect 522 454 556 482
rect 522 386 556 410
rect 522 318 556 338
rect 522 250 556 266
rect 522 182 556 194
rect 411 98 445 114
rect 165 20 177 54
rect 217 20 249 54
rect 285 20 319 54
rect 355 20 387 54
rect 427 20 439 54
<< viali >>
rect 177 1160 183 1194
rect 183 1160 211 1194
rect 249 1160 251 1194
rect 251 1160 283 1194
rect 321 1160 353 1194
rect 353 1160 355 1194
rect 393 1160 421 1194
rect 421 1160 427 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 285 1066 319 1092
rect 285 1058 319 1066
rect 285 998 319 1020
rect 285 986 319 998
rect 285 930 319 948
rect 285 914 319 930
rect 285 862 319 876
rect 285 842 319 862
rect 285 794 319 804
rect 285 770 319 794
rect 285 726 319 732
rect 285 698 319 726
rect 285 658 319 660
rect 285 626 319 658
rect 285 556 319 588
rect 285 554 319 556
rect 285 488 319 516
rect 285 482 319 488
rect 285 420 319 444
rect 285 410 319 420
rect 285 352 319 372
rect 285 338 319 352
rect 285 284 319 300
rect 285 266 319 284
rect 285 216 319 228
rect 285 194 319 216
rect 285 148 319 156
rect 285 122 319 148
rect 411 1066 445 1092
rect 411 1058 445 1066
rect 411 998 445 1020
rect 411 986 445 998
rect 411 930 445 948
rect 411 914 445 930
rect 411 862 445 876
rect 411 842 445 862
rect 411 794 445 804
rect 411 770 445 794
rect 411 726 445 732
rect 411 698 445 726
rect 411 658 445 660
rect 411 626 445 658
rect 411 556 445 588
rect 411 554 445 556
rect 411 488 445 516
rect 411 482 445 488
rect 411 420 445 444
rect 411 410 445 420
rect 411 352 445 372
rect 411 338 445 352
rect 411 284 445 300
rect 411 266 445 284
rect 411 216 445 228
rect 411 194 445 216
rect 411 148 445 156
rect 411 122 445 148
rect 522 1066 556 1092
rect 522 1058 556 1066
rect 522 998 556 1020
rect 522 986 556 998
rect 522 930 556 948
rect 522 914 556 930
rect 522 862 556 876
rect 522 842 556 862
rect 522 794 556 804
rect 522 770 556 794
rect 522 726 556 732
rect 522 698 556 726
rect 522 658 556 660
rect 522 626 556 658
rect 522 556 556 588
rect 522 554 556 556
rect 522 488 556 516
rect 522 482 556 488
rect 522 420 556 444
rect 522 410 556 420
rect 522 352 556 372
rect 522 338 556 352
rect 522 284 556 300
rect 522 266 556 284
rect 522 216 556 228
rect 522 194 556 216
rect 522 148 556 156
rect 522 122 556 148
rect 177 20 183 54
rect 183 20 211 54
rect 249 20 251 54
rect 251 20 283 54
rect 321 20 353 54
rect 353 20 355 54
rect 393 20 421 54
rect 421 20 427 54
<< metal1 >>
rect 165 1194 439 1214
rect 165 1160 177 1194
rect 211 1160 249 1194
rect 283 1160 321 1194
rect 355 1160 393 1194
rect 427 1160 439 1194
rect 165 1148 439 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 276 1098 328 1104
rect 276 1034 328 1046
rect 276 970 328 982
rect 276 914 285 918
rect 319 914 328 918
rect 276 906 328 914
rect 276 842 285 854
rect 319 842 328 854
rect 276 778 285 790
rect 319 778 328 790
rect 276 714 285 726
rect 319 714 328 726
rect 276 660 328 662
rect 276 626 285 660
rect 319 626 328 660
rect 276 588 328 626
rect 276 554 285 588
rect 319 554 328 588
rect 276 516 328 554
rect 276 482 285 516
rect 319 482 328 516
rect 276 444 328 482
rect 276 410 285 444
rect 319 410 328 444
rect 276 372 328 410
rect 276 338 285 372
rect 319 338 328 372
rect 276 300 328 338
rect 276 266 285 300
rect 319 266 328 300
rect 276 228 328 266
rect 276 194 285 228
rect 319 194 328 228
rect 276 156 328 194
rect 276 122 285 156
rect 319 122 328 156
rect 276 110 328 122
rect 402 1092 454 1104
rect 402 1058 411 1092
rect 445 1058 454 1092
rect 402 1020 454 1058
rect 402 986 411 1020
rect 445 986 454 1020
rect 402 948 454 986
rect 402 914 411 948
rect 445 914 454 948
rect 402 876 454 914
rect 402 842 411 876
rect 445 842 454 876
rect 402 804 454 842
rect 402 770 411 804
rect 445 770 454 804
rect 402 732 454 770
rect 402 698 411 732
rect 445 698 454 732
rect 402 660 454 698
rect 402 626 411 660
rect 445 626 454 660
rect 402 588 454 626
rect 402 554 411 588
rect 445 554 454 588
rect 402 552 454 554
rect 402 488 411 500
rect 445 488 454 500
rect 402 424 411 436
rect 445 424 454 436
rect 402 360 411 372
rect 445 360 454 372
rect 402 300 454 308
rect 402 296 411 300
rect 445 296 454 300
rect 402 232 454 244
rect 402 168 454 180
rect 402 110 454 116
rect 510 1092 568 1104
rect 510 1058 522 1092
rect 556 1058 568 1092
rect 510 1020 568 1058
rect 510 986 522 1020
rect 556 986 568 1020
rect 510 948 568 986
rect 510 914 522 948
rect 556 914 568 948
rect 510 876 568 914
rect 510 842 522 876
rect 556 842 568 876
rect 510 804 568 842
rect 510 770 522 804
rect 556 770 568 804
rect 510 732 568 770
rect 510 698 522 732
rect 556 698 568 732
rect 510 660 568 698
rect 510 626 522 660
rect 556 626 568 660
rect 510 588 568 626
rect 510 554 522 588
rect 556 554 568 588
rect 510 516 568 554
rect 510 482 522 516
rect 556 482 568 516
rect 510 444 568 482
rect 510 410 522 444
rect 556 410 568 444
rect 510 372 568 410
rect 510 338 522 372
rect 556 338 568 372
rect 510 300 568 338
rect 510 266 522 300
rect 556 266 568 300
rect 510 228 568 266
rect 510 194 522 228
rect 556 194 568 228
rect 510 156 568 194
rect 510 122 522 156
rect 556 122 568 156
rect 510 110 568 122
rect 165 54 439 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 439 54
rect 165 0 439 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 276 1092 328 1098
rect 276 1058 285 1092
rect 285 1058 319 1092
rect 319 1058 328 1092
rect 276 1046 328 1058
rect 276 1020 328 1034
rect 276 986 285 1020
rect 285 986 319 1020
rect 319 986 328 1020
rect 276 982 328 986
rect 276 948 328 970
rect 276 918 285 948
rect 285 918 319 948
rect 319 918 328 948
rect 276 876 328 906
rect 276 854 285 876
rect 285 854 319 876
rect 319 854 328 876
rect 276 804 328 842
rect 276 790 285 804
rect 285 790 319 804
rect 319 790 328 804
rect 276 770 285 778
rect 285 770 319 778
rect 319 770 328 778
rect 276 732 328 770
rect 276 726 285 732
rect 285 726 319 732
rect 319 726 328 732
rect 276 698 285 714
rect 285 698 319 714
rect 319 698 328 714
rect 276 662 328 698
rect 402 516 454 552
rect 402 500 411 516
rect 411 500 445 516
rect 445 500 454 516
rect 402 482 411 488
rect 411 482 445 488
rect 445 482 454 488
rect 402 444 454 482
rect 402 436 411 444
rect 411 436 445 444
rect 445 436 454 444
rect 402 410 411 424
rect 411 410 445 424
rect 445 410 454 424
rect 402 372 454 410
rect 402 338 411 360
rect 411 338 445 360
rect 445 338 454 360
rect 402 308 454 338
rect 402 266 411 296
rect 411 266 445 296
rect 445 266 454 296
rect 402 244 454 266
rect 402 228 454 232
rect 402 194 411 228
rect 411 194 445 228
rect 445 194 454 228
rect 402 180 454 194
rect 402 156 454 168
rect 402 122 411 156
rect 411 122 445 156
rect 445 122 454 156
rect 402 116 454 122
<< metal2 >>
rect 10 1098 594 1104
rect 10 1046 276 1098
rect 328 1046 594 1098
rect 10 1034 594 1046
rect 10 982 276 1034
rect 328 982 594 1034
rect 10 970 594 982
rect 10 918 276 970
rect 328 918 594 970
rect 10 906 594 918
rect 10 854 276 906
rect 328 854 594 906
rect 10 842 594 854
rect 10 790 276 842
rect 328 790 594 842
rect 10 778 594 790
rect 10 726 276 778
rect 328 726 594 778
rect 10 714 594 726
rect 10 662 276 714
rect 328 662 594 714
rect 10 632 594 662
rect 10 552 594 582
rect 10 500 150 552
rect 202 500 402 552
rect 454 500 594 552
rect 10 488 594 500
rect 10 436 150 488
rect 202 436 402 488
rect 454 436 594 488
rect 10 424 594 436
rect 10 372 150 424
rect 202 372 402 424
rect 454 372 594 424
rect 10 360 594 372
rect 10 308 150 360
rect 202 308 402 360
rect 454 308 594 360
rect 10 296 594 308
rect 10 244 150 296
rect 202 244 402 296
rect 454 244 594 296
rect 10 232 594 244
rect 10 180 150 232
rect 202 180 402 232
rect 454 180 594 232
rect 10 168 594 180
rect 10 116 150 168
rect 202 116 402 168
rect 454 116 594 168
rect 10 110 594 116
<< labels >>
flabel metal2 s 12 781 31 851 0 FreeSans 400 90 0 0 DRAIN
port 1 nsew
flabel metal2 s 14 315 35 379 0 FreeSans 400 90 0 0 SOURCE
port 2 nsew
flabel metal1 s 165 0 439 66 0 FreeSans 300 0 0 0 GATE
port 3 nsew
flabel metal1 s 165 1148 439 1214 0 FreeSans 300 0 0 0 GATE
port 3 nsew
flabel metal1 s 60 732 60 732 7 FreeSans 400 90 0 0 BULK
port 4 nsew
flabel metal1 s 532 732 532 732 7 FreeSans 400 90 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9967686
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9952034
<< end >>
