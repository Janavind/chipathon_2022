magic
tech sky130A
magscale 1 2
timestamp 1669567954
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 348786 700340 348792 700392
rect 348844 700380 348850 700392
rect 364518 700380 364524 700392
rect 348844 700352 364524 700380
rect 348844 700340 348850 700352
rect 364518 700340 364524 700352
rect 364576 700340 364582 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 280798 700312 280804 700324
rect 24360 700284 280804 700312
rect 24360 700272 24366 700284
rect 280798 700272 280804 700284
rect 280856 700272 280862 700324
rect 283834 700272 283840 700324
rect 283892 700312 283898 700324
rect 304258 700312 304264 700324
rect 283892 700284 304264 700312
rect 283892 700272 283898 700284
rect 304258 700272 304264 700284
rect 304316 700272 304322 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 364426 700312 364432 700324
rect 332560 700284 364432 700312
rect 332560 700272 332566 700284
rect 364426 700272 364432 700284
rect 364484 700272 364490 700324
rect 218974 699660 218980 699712
rect 219032 699700 219038 699712
rect 220078 699700 220084 699712
rect 219032 699672 220084 699700
rect 219032 699660 219038 699672
rect 220078 699660 220084 699672
rect 220136 699660 220142 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 363598 698640 363604 698692
rect 363656 698680 363662 698692
rect 364978 698680 364984 698692
rect 363656 698652 364984 698680
rect 363656 698640 363662 698652
rect 364978 698640 364984 698652
rect 365036 698640 365042 698692
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 378778 696940 378784 696992
rect 378836 696980 378842 696992
rect 580166 696980 580172 696992
rect 378836 696952 580172 696980
rect 378836 696940 378842 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 369854 683176 369860 683188
rect 3476 683148 369860 683176
rect 3476 683136 3482 683148
rect 369854 683136 369860 683148
rect 369912 683136 369918 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 298738 670732 298744 670744
rect 3568 670704 298744 670732
rect 3568 670692 3574 670704
rect 298738 670692 298744 670704
rect 298796 670692 298802 670744
rect 360102 670692 360108 670744
rect 360160 670732 360166 670744
rect 580166 670732 580172 670744
rect 360160 670704 580172 670732
rect 360160 670692 360166 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 10318 656928 10324 656940
rect 3476 656900 10324 656928
rect 3476 656888 3482 656900
rect 10318 656888 10324 656900
rect 10376 656888 10382 656940
rect 359458 643084 359464 643136
rect 359516 643124 359522 643136
rect 580166 643124 580172 643136
rect 359516 643096 580172 643124
rect 359516 643084 359522 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 371234 632108 371240 632120
rect 3476 632080 371240 632108
rect 3476 632068 3482 632080
rect 371234 632068 371240 632080
rect 371292 632068 371298 632120
rect 359550 630640 359556 630692
rect 359608 630680 359614 630692
rect 579982 630680 579988 630692
rect 359608 630652 579988 630680
rect 359608 630640 359614 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 311158 618304 311164 618316
rect 3200 618276 311164 618304
rect 3200 618264 3206 618276
rect 311158 618264 311164 618276
rect 311216 618264 311222 618316
rect 382918 616836 382924 616888
rect 382976 616876 382982 616888
rect 580166 616876 580172 616888
rect 382976 616848 580172 616876
rect 382976 616836 382982 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 180058 605860 180064 605872
rect 3292 605832 180064 605860
rect 3292 605820 3298 605832
rect 180058 605820 180064 605832
rect 180116 605820 180122 605872
rect 367738 590656 367744 590708
rect 367796 590696 367802 590708
rect 580166 590696 580172 590708
rect 367796 590668 580172 590696
rect 367796 590656 367802 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 372614 579680 372620 579692
rect 3384 579652 372620 579680
rect 3384 579640 3390 579652
rect 372614 579640 372620 579652
rect 372672 579640 372678 579692
rect 358078 576852 358084 576904
rect 358136 576892 358142 576904
rect 580166 576892 580172 576904
rect 358136 576864 580172 576892
rect 358136 576852 358142 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 376018 563048 376024 563100
rect 376076 563088 376082 563100
rect 580166 563088 580172 563100
rect 376076 563060 580172 563088
rect 376076 563048 376082 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 377398 536800 377404 536852
rect 377456 536840 377462 536852
rect 579890 536840 579896 536852
rect 377456 536812 579896 536840
rect 377456 536800 377462 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 373994 527184 374000 527196
rect 3016 527156 374000 527184
rect 3016 527144 3022 527156
rect 373994 527144 374000 527156
rect 374052 527144 374058 527196
rect 392578 524424 392584 524476
rect 392636 524464 392642 524476
rect 580166 524464 580172 524476
rect 392636 524436 580172 524464
rect 392636 524424 392642 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 262858 514808 262864 514820
rect 3568 514780 262864 514808
rect 3568 514768 3574 514780
rect 262858 514768 262864 514780
rect 262916 514768 262922 514820
rect 361482 511232 361488 511284
rect 361540 511272 361546 511284
rect 580258 511272 580264 511284
rect 361540 511244 580264 511272
rect 361540 511232 361546 511244
rect 580258 511232 580264 511244
rect 580316 511232 580322 511284
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 51718 501004 51724 501016
rect 3108 500976 51724 501004
rect 3108 500964 3114 500976
rect 51718 500964 51724 500976
rect 51776 500964 51782 501016
rect 355318 484372 355324 484424
rect 355376 484412 355382 484424
rect 580166 484412 580172 484424
rect 355376 484384 580172 484412
rect 355376 484372 355382 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 374454 474756 374460 474768
rect 3108 474728 374460 474756
rect 3108 474716 3114 474728
rect 374454 474716 374460 474728
rect 374512 474716 374518 474768
rect 363966 473968 363972 474020
rect 364024 474008 364030 474020
rect 412634 474008 412640 474020
rect 364024 473980 412640 474008
rect 364024 473968 364030 473980
rect 412634 473968 412640 473980
rect 412692 473968 412698 474020
rect 356698 472608 356704 472660
rect 356756 472648 356762 472660
rect 392578 472648 392584 472660
rect 356756 472620 392584 472648
rect 356756 472608 356762 472620
rect 392578 472608 392584 472620
rect 392636 472608 392642 472660
rect 367830 470568 367836 470620
rect 367888 470608 367894 470620
rect 580074 470608 580080 470620
rect 367888 470580 580080 470608
rect 367888 470568 367894 470580
rect 580074 470568 580080 470580
rect 580132 470568 580138 470620
rect 360838 469820 360844 469872
rect 360896 469860 360902 469872
rect 527174 469860 527180 469872
rect 360896 469832 527180 469860
rect 360896 469820 360902 469832
rect 527174 469820 527180 469832
rect 527232 469820 527238 469872
rect 357710 468460 357716 468512
rect 357768 468500 357774 468512
rect 367738 468500 367744 468512
rect 357768 468472 367744 468500
rect 357768 468460 357774 468472
rect 367738 468460 367744 468472
rect 367796 468460 367802 468512
rect 40034 467100 40040 467152
rect 40092 467140 40098 467152
rect 368566 467140 368572 467152
rect 40092 467112 368572 467140
rect 40092 467100 40098 467112
rect 368566 467100 368572 467112
rect 368624 467100 368630 467152
rect 104894 465672 104900 465724
rect 104952 465712 104958 465724
rect 273254 465712 273260 465724
rect 104952 465684 273260 465712
rect 104952 465672 104958 465684
rect 273254 465672 273260 465684
rect 273312 465672 273318 465724
rect 362218 465672 362224 465724
rect 362276 465712 362282 465724
rect 477494 465712 477500 465724
rect 362276 465684 477500 465712
rect 362276 465672 362282 465684
rect 477494 465672 477500 465684
rect 477552 465672 477558 465724
rect 273254 465060 273260 465112
rect 273312 465100 273318 465112
rect 274542 465100 274548 465112
rect 273312 465072 274548 465100
rect 273312 465060 273318 465072
rect 274542 465060 274548 465072
rect 274600 465100 274606 465112
rect 368474 465100 368480 465112
rect 274600 465072 368480 465100
rect 274600 465060 274606 465072
rect 368474 465060 368480 465072
rect 368532 465060 368538 465112
rect 169754 464312 169760 464364
rect 169812 464352 169818 464364
rect 281442 464352 281448 464364
rect 169812 464324 281448 464352
rect 169812 464312 169818 464324
rect 281442 464312 281448 464324
rect 281500 464312 281506 464364
rect 362310 464312 362316 464364
rect 362368 464352 362374 464364
rect 542354 464352 542360 464364
rect 362368 464324 542360 464352
rect 362368 464312 362374 464324
rect 542354 464312 542360 464324
rect 542412 464312 542418 464364
rect 281442 463700 281448 463752
rect 281500 463740 281506 463752
rect 367278 463740 367284 463752
rect 281500 463712 367284 463740
rect 281500 463700 281506 463712
rect 367278 463700 367284 463712
rect 367336 463700 367342 463752
rect 356790 462952 356796 463004
rect 356848 462992 356854 463004
rect 377398 462992 377404 463004
rect 356848 462964 377404 462992
rect 356848 462952 356854 462964
rect 377398 462952 377404 462964
rect 377456 462952 377462 463004
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 315298 462380 315304 462392
rect 3568 462352 315304 462380
rect 3568 462340 3574 462352
rect 315298 462340 315304 462352
rect 315356 462340 315362 462392
rect 364150 461660 364156 461712
rect 364208 461700 364214 461712
rect 396718 461700 396724 461712
rect 364208 461672 396724 461700
rect 364208 461660 364214 461672
rect 396718 461660 396724 461672
rect 396776 461660 396782 461712
rect 234614 461592 234620 461644
rect 234672 461632 234678 461644
rect 365714 461632 365720 461644
rect 234672 461604 365720 461632
rect 234672 461592 234678 461604
rect 365714 461592 365720 461604
rect 365772 461592 365778 461644
rect 357342 460232 357348 460284
rect 357400 460272 357406 460284
rect 367830 460272 367836 460284
rect 357400 460244 367836 460272
rect 357400 460232 357406 460244
rect 367830 460232 367836 460244
rect 367888 460232 367894 460284
rect 363138 460164 363144 460216
rect 363196 460204 363202 460216
rect 429194 460204 429200 460216
rect 363196 460176 429200 460204
rect 363196 460164 363202 460176
rect 429194 460164 429200 460176
rect 429252 460164 429258 460216
rect 361114 458804 361120 458856
rect 361172 458844 361178 458856
rect 558914 458844 558920 458856
rect 361172 458816 558920 458844
rect 361172 458804 361178 458816
rect 558914 458804 558920 458816
rect 558972 458804 558978 458856
rect 334710 457240 334716 457292
rect 334768 457280 334774 457292
rect 373534 457280 373540 457292
rect 334768 457252 373540 457280
rect 334768 457240 334774 457252
rect 373534 457240 373540 457252
rect 373592 457240 373598 457292
rect 323762 457172 323768 457224
rect 323820 457212 323826 457224
rect 384206 457212 384212 457224
rect 323820 457184 384212 457212
rect 323820 457172 323826 457184
rect 384206 457172 384212 457184
rect 384264 457172 384270 457224
rect 320910 457104 320916 457156
rect 320968 457144 320974 457156
rect 381078 457144 381084 457156
rect 320968 457116 381084 457144
rect 320968 457104 320974 457116
rect 381078 457104 381084 457116
rect 381136 457104 381142 457156
rect 315298 457036 315304 457088
rect 315356 457076 315362 457088
rect 375742 457076 375748 457088
rect 315356 457048 375748 457076
rect 315356 457036 315362 457048
rect 375742 457036 375748 457048
rect 375800 457036 375806 457088
rect 320818 456968 320824 457020
rect 320876 457008 320882 457020
rect 381262 457008 381268 457020
rect 320876 456980 381268 457008
rect 320876 456968 320882 456980
rect 381262 456968 381268 456980
rect 381320 456968 381326 457020
rect 311158 456900 311164 456952
rect 311216 456940 311222 456952
rect 311802 456940 311808 456952
rect 311216 456912 311808 456940
rect 311216 456900 311222 456912
rect 311802 456900 311808 456912
rect 311860 456940 311866 456952
rect 372706 456940 372712 456952
rect 311860 456912 372712 456940
rect 311860 456900 311866 456912
rect 372706 456900 372712 456912
rect 372764 456900 372770 456952
rect 371418 456872 371424 456884
rect 306346 456844 371424 456872
rect 298738 456764 298744 456816
rect 298796 456804 298802 456816
rect 299382 456804 299388 456816
rect 298796 456776 299388 456804
rect 298796 456764 298802 456776
rect 299382 456764 299388 456776
rect 299440 456804 299446 456816
rect 306346 456804 306374 456844
rect 371418 456832 371424 456844
rect 371476 456832 371482 456884
rect 299440 456776 306374 456804
rect 299440 456764 299446 456776
rect 355962 456764 355968 456816
rect 356020 456804 356026 456816
rect 580166 456804 580172 456816
rect 356020 456776 580172 456804
rect 356020 456764 356026 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 357618 456084 357624 456136
rect 357676 456124 357682 456136
rect 382918 456124 382924 456136
rect 357676 456096 382924 456124
rect 357676 456084 357682 456096
rect 382918 456084 382924 456096
rect 382976 456084 382982 456136
rect 362862 456016 362868 456068
rect 362920 456056 362926 456068
rect 462314 456056 462320 456068
rect 362920 456028 462320 456056
rect 362920 456016 362926 456028
rect 462314 456016 462320 456028
rect 462372 456016 462378 456068
rect 361666 455948 361672 456000
rect 361724 455988 361730 456000
rect 362310 455988 362316 456000
rect 361724 455960 362316 455988
rect 361724 455948 361730 455960
rect 362310 455948 362316 455960
rect 362368 455948 362374 456000
rect 334618 455880 334624 455932
rect 334676 455920 334682 455932
rect 355502 455920 355508 455932
rect 334676 455892 355508 455920
rect 334676 455880 334682 455892
rect 355502 455880 355508 455892
rect 355560 455880 355566 455932
rect 332134 455812 332140 455864
rect 332192 455852 332198 455864
rect 356146 455852 356152 455864
rect 332192 455824 356152 455852
rect 332192 455812 332198 455824
rect 356146 455812 356152 455824
rect 356204 455852 356210 455864
rect 357342 455852 357348 455864
rect 356204 455824 357348 455852
rect 356204 455812 356210 455824
rect 357342 455812 357348 455824
rect 357400 455812 357406 455864
rect 332042 455744 332048 455796
rect 332100 455784 332106 455796
rect 359550 455784 359556 455796
rect 332100 455756 359556 455784
rect 332100 455744 332106 455756
rect 359550 455744 359556 455756
rect 359608 455744 359614 455796
rect 333330 455676 333336 455728
rect 333388 455716 333394 455728
rect 361666 455716 361672 455728
rect 333388 455688 361672 455716
rect 333388 455676 333394 455688
rect 361666 455676 361672 455688
rect 361724 455676 361730 455728
rect 332226 455608 332232 455660
rect 332284 455648 332290 455660
rect 364426 455648 364432 455660
rect 332284 455620 364432 455648
rect 332284 455608 332290 455620
rect 364426 455608 364432 455620
rect 364484 455608 364490 455660
rect 333422 455540 333428 455592
rect 333480 455580 333486 455592
rect 380158 455580 380164 455592
rect 333480 455552 380164 455580
rect 333480 455540 333486 455552
rect 380158 455540 380164 455552
rect 380216 455540 380222 455592
rect 302878 455472 302884 455524
rect 302936 455512 302942 455524
rect 362218 455512 362224 455524
rect 302936 455484 362224 455512
rect 302936 455472 302942 455484
rect 362218 455472 362224 455484
rect 362276 455472 362282 455524
rect 322290 455404 322296 455456
rect 322348 455444 322354 455456
rect 383102 455444 383108 455456
rect 322348 455416 383108 455444
rect 322348 455404 322354 455416
rect 383102 455404 383108 455416
rect 383160 455404 383166 455456
rect 281350 454928 281356 454980
rect 281408 454968 281414 454980
rect 351914 454968 351920 454980
rect 281408 454940 351920 454968
rect 281408 454928 281414 454940
rect 351914 454928 351920 454940
rect 351972 454928 351978 454980
rect 319530 454860 319536 454912
rect 319588 454900 319594 454912
rect 379790 454900 379796 454912
rect 319588 454872 379796 454900
rect 319588 454860 319594 454872
rect 379790 454860 379796 454872
rect 379848 454860 379854 454912
rect 294690 454792 294696 454844
rect 294748 454832 294754 454844
rect 354674 454832 354680 454844
rect 294748 454804 354680 454832
rect 294748 454792 294754 454804
rect 354674 454792 354680 454804
rect 354732 454792 354738 454844
rect 357434 454792 357440 454844
rect 357492 454832 357498 454844
rect 376018 454832 376024 454844
rect 357492 454804 376024 454832
rect 357492 454792 357498 454804
rect 376018 454792 376024 454804
rect 376076 454792 376082 454844
rect 337930 454724 337936 454776
rect 337988 454764 337994 454776
rect 357618 454764 357624 454776
rect 337988 454736 357624 454764
rect 337988 454724 337994 454736
rect 357618 454724 357624 454736
rect 357676 454764 357682 454776
rect 358446 454764 358452 454776
rect 357676 454736 358452 454764
rect 357676 454724 357682 454736
rect 358446 454724 358452 454736
rect 358504 454724 358510 454776
rect 337286 454656 337292 454708
rect 337344 454696 337350 454708
rect 362034 454696 362040 454708
rect 337344 454668 362040 454696
rect 337344 454656 337350 454668
rect 362034 454656 362040 454668
rect 362092 454696 362098 454708
rect 494054 454696 494060 454708
rect 362092 454668 494060 454696
rect 362092 454656 362098 454668
rect 494054 454656 494060 454668
rect 494112 454656 494118 454708
rect 337378 454588 337384 454640
rect 337436 454628 337442 454640
rect 363138 454628 363144 454640
rect 337436 454600 363144 454628
rect 337436 454588 337442 454600
rect 363138 454588 363144 454600
rect 363196 454588 363202 454640
rect 319622 454520 319628 454572
rect 319680 454560 319686 454572
rect 376754 454560 376760 454572
rect 319680 454532 376760 454560
rect 319680 454520 319686 454532
rect 376754 454520 376760 454532
rect 376812 454520 376818 454572
rect 319714 454452 319720 454504
rect 319772 454492 319778 454504
rect 378686 454492 378692 454504
rect 319772 454464 378692 454492
rect 319772 454452 319778 454464
rect 378686 454452 378692 454464
rect 378744 454452 378750 454504
rect 293862 454384 293868 454436
rect 293920 454424 293926 454436
rect 353294 454424 353300 454436
rect 293920 454396 353300 454424
rect 293920 454384 293926 454396
rect 353294 454384 353300 454396
rect 353352 454384 353358 454436
rect 318242 454316 318248 454368
rect 318300 454356 318306 454368
rect 378318 454356 378324 454368
rect 318300 454328 378324 454356
rect 318300 454316 318306 454328
rect 378318 454316 378324 454328
rect 378376 454316 378382 454368
rect 316862 454248 316868 454300
rect 316920 454288 316926 454300
rect 376938 454288 376944 454300
rect 316920 454260 376944 454288
rect 316920 454248 316926 454260
rect 376938 454248 376944 454260
rect 376996 454248 377002 454300
rect 340690 454180 340696 454232
rect 340748 454220 340754 454232
rect 357434 454220 357440 454232
rect 340748 454192 357440 454220
rect 340748 454180 340754 454192
rect 357434 454180 357440 454192
rect 357492 454180 357498 454232
rect 336458 454112 336464 454164
rect 336516 454152 336522 454164
rect 355042 454152 355048 454164
rect 336516 454124 355048 454152
rect 336516 454112 336522 454124
rect 355042 454112 355048 454124
rect 355100 454112 355106 454164
rect 337470 454044 337476 454096
rect 337528 454084 337534 454096
rect 374270 454084 374276 454096
rect 337528 454056 374276 454084
rect 337528 454044 337534 454056
rect 374270 454044 374276 454056
rect 374328 454044 374334 454096
rect 323578 453568 323584 453620
rect 323636 453608 323642 453620
rect 383838 453608 383844 453620
rect 323636 453580 383844 453608
rect 323636 453568 323642 453580
rect 383838 453568 383844 453580
rect 383896 453568 383902 453620
rect 318058 453500 318064 453552
rect 318116 453540 318122 453552
rect 378410 453540 378416 453552
rect 318116 453512 378416 453540
rect 318116 453500 318122 453512
rect 378410 453500 378416 453512
rect 378468 453500 378474 453552
rect 335262 453432 335268 453484
rect 335320 453472 335326 453484
rect 359090 453472 359096 453484
rect 335320 453444 359096 453472
rect 335320 453432 335326 453444
rect 359090 453432 359096 453444
rect 359148 453432 359154 453484
rect 361390 453432 361396 453484
rect 361448 453472 361454 453484
rect 378778 453472 378784 453484
rect 361448 453444 378784 453472
rect 361448 453432 361454 453444
rect 378778 453432 378784 453444
rect 378836 453432 378842 453484
rect 299474 453364 299480 453416
rect 299532 453404 299538 453416
rect 365070 453404 365076 453416
rect 299532 453376 365076 453404
rect 299532 453364 299538 453376
rect 365070 453364 365076 453376
rect 365128 453364 365134 453416
rect 356238 453296 356244 453348
rect 356296 453336 356302 453348
rect 580350 453336 580356 453348
rect 356296 453308 580356 453336
rect 356296 453296 356302 453308
rect 580350 453296 580356 453308
rect 580408 453296 580414 453348
rect 335170 453228 335176 453280
rect 335228 453268 335234 453280
rect 362402 453268 362408 453280
rect 335228 453240 362408 453268
rect 335228 453228 335234 453240
rect 362402 453228 362408 453240
rect 362460 453268 362466 453280
rect 362862 453268 362868 453280
rect 362460 453240 362868 453268
rect 362460 453228 362466 453240
rect 362862 453228 362868 453240
rect 362920 453228 362926 453280
rect 315390 453160 315396 453212
rect 315448 453200 315454 453212
rect 367094 453200 367100 453212
rect 315448 453172 367100 453200
rect 315448 453160 315454 453172
rect 367094 453160 367100 453172
rect 367152 453160 367158 453212
rect 316678 453092 316684 453144
rect 316736 453132 316742 453144
rect 371326 453132 371332 453144
rect 316736 453104 371332 453132
rect 316736 453092 316742 453104
rect 371326 453092 371332 453104
rect 371384 453092 371390 453144
rect 318150 453024 318156 453076
rect 318208 453064 318214 453076
rect 377214 453064 377220 453076
rect 318208 453036 377220 453064
rect 318208 453024 318214 453036
rect 377214 453024 377220 453036
rect 377272 453024 377278 453076
rect 316770 452956 316776 453008
rect 316828 452996 316834 453008
rect 376110 452996 376116 453008
rect 316828 452968 376116 452996
rect 316828 452956 316834 452968
rect 376110 452956 376116 452968
rect 376168 452956 376174 453008
rect 294782 452888 294788 452940
rect 294840 452928 294846 452940
rect 354122 452928 354128 452940
rect 294840 452900 354128 452928
rect 294840 452888 294846 452900
rect 354122 452888 354128 452900
rect 354180 452888 354186 452940
rect 322198 452820 322204 452872
rect 322256 452860 322262 452872
rect 381630 452860 381636 452872
rect 322256 452832 381636 452860
rect 322256 452820 322262 452832
rect 381630 452820 381636 452832
rect 381688 452820 381694 452872
rect 324958 452752 324964 452804
rect 325016 452792 325022 452804
rect 385034 452792 385040 452804
rect 325016 452764 385040 452792
rect 325016 452752 325022 452764
rect 385034 452752 385040 452764
rect 385092 452752 385098 452804
rect 341978 452684 341984 452736
rect 342036 452724 342042 452736
rect 353018 452724 353024 452736
rect 342036 452696 353024 452724
rect 342036 452684 342042 452696
rect 353018 452684 353024 452696
rect 353076 452684 353082 452736
rect 340046 452616 340052 452668
rect 340104 452656 340110 452668
rect 356238 452656 356244 452668
rect 340104 452628 356244 452656
rect 340104 452616 340110 452628
rect 356238 452616 356244 452628
rect 356296 452616 356302 452668
rect 355410 452548 355416 452600
rect 355468 452588 355474 452600
rect 355962 452588 355968 452600
rect 355468 452560 355968 452588
rect 355468 452548 355474 452560
rect 355962 452548 355968 452560
rect 356020 452548 356026 452600
rect 376754 452548 376760 452600
rect 376812 452588 376818 452600
rect 379054 452588 379060 452600
rect 376812 452560 379060 452588
rect 376812 452548 376818 452560
rect 379054 452548 379060 452560
rect 379112 452548 379118 452600
rect 278590 452140 278596 452192
rect 278648 452180 278654 452192
rect 348510 452180 348516 452192
rect 278648 452152 348516 452180
rect 278648 452140 278654 452152
rect 348510 452140 348516 452152
rect 348568 452140 348574 452192
rect 294598 452072 294604 452124
rect 294656 452112 294662 452124
rect 350626 452112 350632 452124
rect 294656 452084 350632 452112
rect 294656 452072 294662 452084
rect 350626 452072 350632 452084
rect 350684 452072 350690 452124
rect 340138 452004 340144 452056
rect 340196 452044 340202 452056
rect 385678 452044 385684 452056
rect 340196 452016 385684 452044
rect 340196 452004 340202 452016
rect 385678 452004 385684 452016
rect 385736 452004 385742 452056
rect 308490 451936 308496 451988
rect 308548 451976 308554 451988
rect 367186 451976 367192 451988
rect 308548 451948 367192 451976
rect 308548 451936 308554 451948
rect 367186 451936 367192 451948
rect 367244 451936 367250 451988
rect 371326 451936 371332 451988
rect 371384 451976 371390 451988
rect 376754 451976 376760 451988
rect 371384 451948 376760 451976
rect 371384 451936 371390 451948
rect 376754 451936 376760 451948
rect 376812 451936 376818 451988
rect 300118 451868 300124 451920
rect 300176 451908 300182 451920
rect 355410 451908 355416 451920
rect 300176 451880 355416 451908
rect 300176 451868 300182 451880
rect 355410 451868 355416 451880
rect 355468 451868 355474 451920
rect 363322 451868 363328 451920
rect 363380 451908 363386 451920
rect 365714 451908 365720 451920
rect 363380 451880 365720 451908
rect 363380 451868 363386 451880
rect 365714 451868 365720 451880
rect 365772 451908 365778 451920
rect 366174 451908 366180 451920
rect 365772 451880 366180 451908
rect 365772 451868 365778 451880
rect 366174 451868 366180 451880
rect 366232 451868 366238 451920
rect 342162 451800 342168 451852
rect 342220 451840 342226 451852
rect 353662 451840 353668 451852
rect 342220 451812 353668 451840
rect 342220 451800 342226 451812
rect 353662 451800 353668 451812
rect 353720 451800 353726 451852
rect 363598 451800 363604 451852
rect 363656 451840 363662 451852
rect 364058 451840 364064 451852
rect 363656 451812 364064 451840
rect 363656 451800 363662 451812
rect 364058 451800 364064 451812
rect 364116 451800 364122 451852
rect 342346 451732 342352 451784
rect 342404 451772 342410 451784
rect 365806 451772 365812 451784
rect 342404 451744 365812 451772
rect 342404 451732 342410 451744
rect 365806 451732 365812 451744
rect 365864 451732 365870 451784
rect 341518 451664 341524 451716
rect 341576 451704 341582 451716
rect 374638 451704 374644 451716
rect 341576 451676 374644 451704
rect 341576 451664 341582 451676
rect 374638 451664 374644 451676
rect 374696 451664 374702 451716
rect 340966 451596 340972 451648
rect 341024 451636 341030 451648
rect 341024 451608 373994 451636
rect 341024 451596 341030 451608
rect 309778 451528 309784 451580
rect 309836 451568 309842 451580
rect 352650 451568 352656 451580
rect 309836 451540 352656 451568
rect 309836 451528 309842 451540
rect 352650 451528 352656 451540
rect 352708 451528 352714 451580
rect 354582 451528 354588 451580
rect 354640 451568 354646 451580
rect 373966 451568 373994 451608
rect 384574 451568 384580 451580
rect 354640 451540 360194 451568
rect 373966 451540 384580 451568
rect 354640 451528 354646 451540
rect 337562 451460 337568 451512
rect 337620 451500 337626 451512
rect 349246 451500 349252 451512
rect 337620 451472 349252 451500
rect 337620 451460 337626 451472
rect 349246 451460 349252 451472
rect 349304 451460 349310 451512
rect 360166 451500 360194 451540
rect 384574 451528 384580 451540
rect 384632 451528 384638 451580
rect 366542 451500 366548 451512
rect 360166 451472 366548 451500
rect 366542 451460 366548 451472
rect 366600 451460 366606 451512
rect 341702 451392 341708 451444
rect 341760 451432 341766 451444
rect 382366 451432 382372 451444
rect 341760 451404 382372 451432
rect 341760 451392 341766 451404
rect 382366 451392 382372 451404
rect 382424 451392 382430 451444
rect 339402 451324 339408 451376
rect 339460 451364 339466 451376
rect 352558 451364 352564 451376
rect 339460 451336 352564 451364
rect 339460 451324 339466 451336
rect 352558 451324 352564 451336
rect 352616 451324 352622 451376
rect 352650 451324 352656 451376
rect 352708 451364 352714 451376
rect 364702 451364 364708 451376
rect 352708 451336 364708 451364
rect 352708 451324 352714 451336
rect 364702 451324 364708 451336
rect 364760 451324 364766 451376
rect 367094 451324 367100 451376
rect 367152 451364 367158 451376
rect 375374 451364 375380 451376
rect 367152 451336 375380 451364
rect 367152 451324 367158 451336
rect 375374 451324 375380 451336
rect 375432 451324 375438 451376
rect 338850 451256 338856 451308
rect 338908 451296 338914 451308
rect 351454 451296 351460 451308
rect 338908 451268 351460 451296
rect 338908 451256 338914 451268
rect 351454 451256 351460 451268
rect 351512 451256 351518 451308
rect 355042 451256 355048 451308
rect 355100 451296 355106 451308
rect 357434 451296 357440 451308
rect 355100 451268 357440 451296
rect 355100 451256 355106 451268
rect 357434 451256 357440 451268
rect 357492 451256 357498 451308
rect 365714 451256 365720 451308
rect 365772 451296 365778 451308
rect 369946 451296 369952 451308
rect 365772 451268 369952 451296
rect 365772 451256 365778 451268
rect 369946 451256 369952 451268
rect 370004 451256 370010 451308
rect 297450 450780 297456 450832
rect 297508 450820 297514 450832
rect 357710 450820 357716 450832
rect 297508 450792 357716 450820
rect 297508 450780 297514 450792
rect 357710 450780 357716 450792
rect 357768 450780 357774 450832
rect 300302 450712 300308 450764
rect 300360 450752 300366 450764
rect 360194 450752 360200 450764
rect 300360 450724 360200 450752
rect 300360 450712 300366 450724
rect 360194 450712 360200 450724
rect 360252 450752 360258 450764
rect 361390 450752 361396 450764
rect 360252 450724 361396 450752
rect 360252 450712 360258 450724
rect 361390 450712 361396 450724
rect 361448 450712 361454 450764
rect 266354 450644 266360 450696
rect 266412 450684 266418 450696
rect 304994 450684 305000 450696
rect 266412 450656 305000 450684
rect 266412 450644 266418 450656
rect 304994 450644 305000 450656
rect 305052 450644 305058 450696
rect 321002 450644 321008 450696
rect 321060 450684 321066 450696
rect 380526 450684 380532 450696
rect 321060 450656 380532 450684
rect 321060 450644 321066 450656
rect 380526 450644 380532 450656
rect 380584 450644 380590 450696
rect 201494 450576 201500 450628
rect 201552 450616 201558 450628
rect 201552 450588 296714 450616
rect 201552 450576 201558 450588
rect 136634 450508 136640 450560
rect 136692 450548 136698 450560
rect 296686 450548 296714 450588
rect 319438 450576 319444 450628
rect 319496 450616 319502 450628
rect 379422 450616 379428 450628
rect 319496 450588 379428 450616
rect 319496 450576 319502 450588
rect 379422 450576 379428 450588
rect 379480 450576 379486 450628
rect 306374 450548 306380 450560
rect 136692 450520 277394 450548
rect 296686 450520 306380 450548
rect 136692 450508 136698 450520
rect 277366 450208 277394 450520
rect 306374 450508 306380 450520
rect 306432 450548 306438 450560
rect 354582 450548 354588 450560
rect 306432 450520 354588 450548
rect 306432 450508 306438 450520
rect 354582 450508 354588 450520
rect 354640 450508 354646 450560
rect 357434 450508 357440 450560
rect 357492 450548 357498 450560
rect 580258 450548 580264 450560
rect 357492 450520 580264 450548
rect 357492 450508 357498 450520
rect 580258 450508 580264 450520
rect 580316 450508 580322 450560
rect 323670 450440 323676 450492
rect 323728 450480 323734 450492
rect 382734 450480 382740 450492
rect 323728 450452 382740 450480
rect 323728 450440 323734 450452
rect 382734 450440 382740 450452
rect 382792 450440 382798 450492
rect 314010 450372 314016 450424
rect 314068 450412 314074 450424
rect 373166 450412 373172 450424
rect 314068 450384 373172 450412
rect 314068 450372 314074 450384
rect 373166 450372 373172 450384
rect 373224 450372 373230 450424
rect 301498 450304 301504 450356
rect 301556 450344 301562 450356
rect 361022 450344 361028 450356
rect 301556 450316 361028 450344
rect 301556 450304 301562 450316
rect 361022 450304 361028 450316
rect 361080 450304 361086 450356
rect 297358 450236 297364 450288
rect 297416 450276 297422 450288
rect 356882 450276 356888 450288
rect 297416 450248 356888 450276
rect 297416 450236 297422 450248
rect 356882 450236 356888 450248
rect 356940 450236 356946 450288
rect 279878 450208 279884 450220
rect 277366 450180 279884 450208
rect 279878 450168 279884 450180
rect 279936 450208 279942 450220
rect 367876 450208 367882 450220
rect 279936 450180 367882 450208
rect 279936 450168 279942 450180
rect 367876 450168 367882 450180
rect 367934 450168 367940 450220
rect 371234 450168 371240 450220
rect 371292 450208 371298 450220
rect 371694 450208 371700 450220
rect 371292 450180 371700 450208
rect 371292 450168 371298 450180
rect 371694 450168 371700 450180
rect 371752 450168 371758 450220
rect 338758 450100 338764 450152
rect 338816 450140 338822 450152
rect 349108 450140 349114 450152
rect 338816 450112 349114 450140
rect 338816 450100 338822 450112
rect 349108 450100 349114 450112
rect 349166 450100 349172 450152
rect 354122 450100 354128 450152
rect 354180 450140 354186 450152
rect 388438 450140 388444 450152
rect 354180 450112 388444 450140
rect 354180 450100 354186 450112
rect 388438 450100 388444 450112
rect 388496 450100 388502 450152
rect 304994 450032 305000 450084
rect 305052 450072 305058 450084
rect 365438 450072 365444 450084
rect 305052 450044 365444 450072
rect 305052 450032 305058 450044
rect 365438 450032 365444 450044
rect 365496 450032 365502 450084
rect 340322 449964 340328 450016
rect 340380 450004 340386 450016
rect 372062 450004 372068 450016
rect 340380 449976 372068 450004
rect 340380 449964 340386 449976
rect 372062 449964 372068 449976
rect 372120 449964 372126 450016
rect 340782 449896 340788 449948
rect 340840 449936 340846 449948
rect 348142 449936 348148 449948
rect 340840 449908 348148 449936
rect 340840 449896 340846 449908
rect 348142 449896 348148 449908
rect 348200 449896 348206 449948
rect 354858 449896 354864 449948
rect 354916 449936 354922 449948
rect 389818 449936 389824 449948
rect 354916 449908 389824 449936
rect 354916 449896 354922 449908
rect 389818 449896 389824 449908
rect 389876 449896 389882 449948
rect 363322 449596 363328 449608
rect 350506 449568 363328 449596
rect 350506 449528 350534 449568
rect 363322 449556 363328 449568
rect 363380 449556 363386 449608
rect 331186 449500 350534 449528
rect 307018 449284 307024 449336
rect 307076 449324 307082 449336
rect 331186 449324 331214 449500
rect 342438 449420 342444 449472
rect 342496 449460 342502 449472
rect 349614 449460 349620 449472
rect 342496 449432 349620 449460
rect 342496 449420 342502 449432
rect 349614 449420 349620 449432
rect 349672 449420 349678 449472
rect 351086 449460 351092 449472
rect 349724 449432 351092 449460
rect 307076 449296 331214 449324
rect 307076 449284 307082 449296
rect 342070 449284 342076 449336
rect 342128 449324 342134 449336
rect 349724 449324 349752 449432
rect 351086 449420 351092 449432
rect 351144 449420 351150 449472
rect 369854 449420 369860 449472
rect 369912 449460 369918 449472
rect 370590 449460 370596 449472
rect 369912 449432 370596 449460
rect 369912 449420 369918 449432
rect 370590 449420 370596 449432
rect 370648 449420 370654 449472
rect 358078 449392 358084 449404
rect 350506 449364 358084 449392
rect 350506 449324 350534 449364
rect 358078 449352 358084 449364
rect 358136 449352 358142 449404
rect 363966 449392 363972 449404
rect 360166 449364 363972 449392
rect 342128 449296 349752 449324
rect 349816 449296 350534 449324
rect 342128 449284 342134 449296
rect 304350 449216 304356 449268
rect 304408 449256 304414 449268
rect 330202 449256 330208 449268
rect 304408 449228 330208 449256
rect 304408 449216 304414 449228
rect 330202 449216 330208 449228
rect 330260 449216 330266 449268
rect 333256 449228 338114 449256
rect 298738 449148 298744 449200
rect 298796 449188 298802 449200
rect 333256 449188 333284 449228
rect 298796 449160 333284 449188
rect 338086 449188 338114 449228
rect 349816 449188 349844 449296
rect 338086 449160 349844 449188
rect 298796 449148 298802 449160
rect 330202 449080 330208 449132
rect 330260 449120 330266 449132
rect 330260 449092 340874 449120
rect 330260 449080 330266 449092
rect 340846 449052 340874 449092
rect 360166 449052 360194 449364
rect 363966 449352 363972 449364
rect 364024 449352 364030 449404
rect 340846 449024 360194 449052
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 8938 448576 8944 448588
rect 3200 448548 8944 448576
rect 3200 448536 3206 448548
rect 8938 448536 8944 448548
rect 8996 448536 9002 448588
rect 277762 448536 277768 448588
rect 277820 448576 277826 448588
rect 342438 448576 342444 448588
rect 277820 448548 342444 448576
rect 277820 448536 277826 448548
rect 342438 448536 342444 448548
rect 342496 448536 342502 448588
rect 325050 445000 325056 445052
rect 325108 445040 325114 445052
rect 340966 445040 340972 445052
rect 325108 445012 340972 445040
rect 325108 445000 325114 445012
rect 340966 445000 340972 445012
rect 341024 445000 341030 445052
rect 322382 438132 322388 438184
rect 322440 438172 322446 438184
rect 340966 438172 340972 438184
rect 322440 438144 340972 438172
rect 322440 438132 322446 438144
rect 340966 438132 340972 438144
rect 341024 438132 341030 438184
rect 287698 435344 287704 435396
rect 287756 435384 287762 435396
rect 340874 435384 340880 435396
rect 287756 435356 340880 435384
rect 287756 435344 287762 435356
rect 340874 435344 340880 435356
rect 340932 435344 340938 435396
rect 389818 431876 389824 431928
rect 389876 431916 389882 431928
rect 580166 431916 580172 431928
rect 389876 431888 580172 431916
rect 389876 431876 389882 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 311158 422328 311164 422340
rect 3568 422300 311164 422328
rect 3568 422288 3574 422300
rect 311158 422288 311164 422300
rect 311216 422288 311222 422340
rect 289722 418752 289728 418804
rect 289780 418792 289786 418804
rect 337562 418792 337568 418804
rect 289780 418764 337568 418792
rect 289780 418752 289786 418764
rect 337562 418752 337568 418764
rect 337620 418752 337626 418804
rect 262858 417392 262864 417444
rect 262916 417432 262922 417444
rect 315482 417432 315488 417444
rect 262916 417404 315488 417432
rect 262916 417392 262922 417404
rect 315482 417392 315488 417404
rect 315540 417392 315546 417444
rect 8938 416712 8944 416764
rect 8996 416752 9002 416764
rect 314746 416752 314752 416764
rect 8996 416724 314752 416752
rect 8996 416712 9002 416724
rect 314746 416712 314752 416724
rect 314804 416752 314810 416764
rect 315390 416752 315396 416764
rect 314804 416724 315396 416752
rect 314804 416712 314810 416724
rect 315390 416712 315396 416724
rect 315448 416712 315454 416764
rect 311158 415420 311164 415472
rect 311216 415460 311222 415472
rect 316770 415460 316776 415472
rect 311216 415432 316776 415460
rect 311216 415420 311222 415432
rect 316770 415420 316776 415432
rect 316828 415420 316834 415472
rect 51718 414672 51724 414724
rect 51776 414712 51782 414724
rect 313918 414712 313924 414724
rect 51776 414684 313924 414712
rect 51776 414672 51782 414684
rect 313918 414672 313924 414684
rect 313976 414672 313982 414724
rect 313918 413924 313924 413976
rect 313976 413964 313982 413976
rect 337470 413964 337476 413976
rect 313976 413936 337476 413964
rect 313976 413924 313982 413936
rect 337470 413924 337476 413936
rect 337528 413924 337534 413976
rect 4798 413856 4804 413908
rect 4856 413896 4862 413908
rect 313274 413896 313280 413908
rect 4856 413868 313280 413896
rect 4856 413856 4862 413868
rect 313274 413856 313280 413868
rect 313332 413896 313338 413908
rect 314010 413896 314016 413908
rect 313332 413868 314016 413896
rect 313332 413856 313338 413868
rect 314010 413856 314016 413868
rect 314068 413856 314074 413908
rect 180058 411884 180064 411936
rect 180116 411924 180122 411936
rect 311894 411924 311900 411936
rect 180116 411896 311900 411924
rect 180116 411884 180122 411896
rect 311894 411884 311900 411896
rect 311952 411884 311958 411936
rect 311894 411204 311900 411256
rect 311952 411244 311958 411256
rect 312630 411244 312636 411256
rect 311952 411216 312636 411244
rect 311952 411204 311958 411216
rect 312630 411204 312636 411216
rect 312688 411244 312694 411256
rect 340322 411244 340328 411256
rect 312688 411216 340328 411244
rect 312688 411204 312694 411216
rect 340322 411204 340328 411216
rect 340380 411204 340386 411256
rect 10318 410524 10324 410576
rect 10376 410564 10382 410576
rect 311250 410564 311256 410576
rect 10376 410536 311256 410564
rect 10376 410524 10382 410536
rect 311250 410524 311256 410536
rect 311308 410524 311314 410576
rect 286410 409096 286416 409148
rect 286468 409136 286474 409148
rect 340230 409136 340236 409148
rect 286468 409108 340236 409136
rect 286468 409096 286474 409108
rect 340230 409096 340236 409108
rect 340288 409096 340294 409148
rect 326338 407736 326344 407788
rect 326396 407776 326402 407788
rect 340138 407776 340144 407788
rect 326396 407748 340144 407776
rect 326396 407736 326402 407748
rect 340138 407736 340144 407748
rect 340196 407736 340202 407788
rect 291930 406444 291936 406496
rect 291988 406484 291994 406496
rect 338850 406484 338856 406496
rect 291988 406456 338856 406484
rect 291988 406444 291994 406456
rect 338850 406444 338856 406456
rect 338908 406444 338914 406496
rect 88334 406376 88340 406428
rect 88392 406416 88398 406428
rect 309962 406416 309968 406428
rect 88392 406388 309968 406416
rect 88392 406376 88398 406388
rect 309962 406376 309968 406388
rect 310020 406376 310026 406428
rect 4154 405628 4160 405680
rect 4212 405668 4218 405680
rect 316034 405668 316040 405680
rect 4212 405640 316040 405668
rect 4212 405628 4218 405640
rect 316034 405628 316040 405640
rect 316092 405668 316098 405680
rect 316862 405668 316868 405680
rect 316092 405640 316868 405668
rect 316092 405628 316098 405640
rect 316862 405628 316868 405640
rect 316920 405628 316926 405680
rect 388990 405628 388996 405680
rect 389048 405668 389054 405680
rect 580166 405668 580172 405680
rect 389048 405640 580172 405668
rect 389048 405628 389054 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 309962 405560 309968 405612
rect 310020 405600 310026 405612
rect 334802 405600 334808 405612
rect 310020 405572 334808 405600
rect 310020 405560 310026 405572
rect 334802 405560 334808 405572
rect 334860 405560 334866 405612
rect 315482 404268 315488 404320
rect 315540 404308 315546 404320
rect 340966 404308 340972 404320
rect 315540 404280 340972 404308
rect 315540 404268 315546 404280
rect 340966 404268 340972 404280
rect 341024 404268 341030 404320
rect 299382 403588 299388 403640
rect 299440 403628 299446 403640
rect 310514 403628 310520 403640
rect 299440 403600 310520 403628
rect 299440 403588 299446 403600
rect 310514 403588 310520 403600
rect 310572 403588 310578 403640
rect 3418 402228 3424 402280
rect 3476 402268 3482 402280
rect 313274 402268 313280 402280
rect 3476 402240 313280 402268
rect 3476 402228 3482 402240
rect 313274 402228 313280 402240
rect 313332 402228 313338 402280
rect 316126 401616 316132 401668
rect 316184 401656 316190 401668
rect 316770 401656 316776 401668
rect 316184 401628 316776 401656
rect 316184 401616 316190 401628
rect 316770 401616 316776 401628
rect 316828 401616 316834 401668
rect 313274 401548 313280 401600
rect 313332 401588 313338 401600
rect 314010 401588 314016 401600
rect 313332 401560 314016 401588
rect 313332 401548 313338 401560
rect 314010 401548 314016 401560
rect 314068 401588 314074 401600
rect 334710 401588 334716 401600
rect 314068 401560 334716 401588
rect 314068 401548 314074 401560
rect 334710 401548 334716 401560
rect 334768 401548 334774 401600
rect 341794 400936 341800 400988
rect 341852 400976 341858 400988
rect 341852 400948 357434 400976
rect 341852 400936 341858 400948
rect 341426 400840 341432 400852
rect 338086 400812 341432 400840
rect 338086 400636 338114 400812
rect 341426 400800 341432 400812
rect 341484 400800 341490 400852
rect 341518 400800 341524 400852
rect 341576 400840 341582 400852
rect 342254 400840 342260 400852
rect 341576 400812 342260 400840
rect 341576 400800 341582 400812
rect 342254 400800 342260 400812
rect 342312 400800 342318 400852
rect 335326 400608 338114 400636
rect 357406 400636 357434 400948
rect 357406 400608 366496 400636
rect 281258 400528 281264 400580
rect 281316 400568 281322 400580
rect 335326 400568 335354 400608
rect 281316 400540 335354 400568
rect 281316 400528 281322 400540
rect 341886 400528 341892 400580
rect 341944 400568 341950 400580
rect 341944 400540 347866 400568
rect 341944 400528 341950 400540
rect 279970 400460 279976 400512
rect 280028 400500 280034 400512
rect 342254 400500 342260 400512
rect 280028 400472 342260 400500
rect 280028 400460 280034 400472
rect 342254 400460 342260 400472
rect 342312 400460 342318 400512
rect 347838 400500 347866 400540
rect 342364 400472 347774 400500
rect 347838 400472 357434 400500
rect 271690 400392 271696 400444
rect 271748 400432 271754 400444
rect 271748 400404 342208 400432
rect 271748 400392 271754 400404
rect 277118 400324 277124 400376
rect 277176 400364 277182 400376
rect 341426 400364 341432 400376
rect 277176 400336 341432 400364
rect 277176 400324 277182 400336
rect 341426 400324 341432 400336
rect 341484 400324 341490 400376
rect 281074 400256 281080 400308
rect 281132 400296 281138 400308
rect 341886 400296 341892 400308
rect 281132 400268 341892 400296
rect 281132 400256 281138 400268
rect 341886 400256 341892 400268
rect 341944 400256 341950 400308
rect 342180 400296 342208 400404
rect 342254 400324 342260 400376
rect 342312 400364 342318 400376
rect 342364 400364 342392 400472
rect 347746 400432 347774 400472
rect 342312 400336 342392 400364
rect 342456 400404 346716 400432
rect 347746 400404 349890 400432
rect 342312 400324 342318 400336
rect 342456 400296 342484 400404
rect 342180 400268 342484 400296
rect 345998 400336 346256 400364
rect 274266 400188 274272 400240
rect 274324 400228 274330 400240
rect 345998 400228 346026 400336
rect 274324 400200 346026 400228
rect 274324 400188 274330 400200
rect 341334 400120 341340 400172
rect 341392 400160 341398 400172
rect 341392 400132 346118 400160
rect 341392 400120 341398 400132
rect 335326 400064 338114 400092
rect 331858 399644 331864 399696
rect 331916 399684 331922 399696
rect 335326 399684 335354 400064
rect 338086 400024 338114 400064
rect 339862 400052 339868 400104
rect 339920 400092 339926 400104
rect 341610 400092 341616 400104
rect 339920 400064 341616 400092
rect 339920 400052 339926 400064
rect 341610 400052 341616 400064
rect 341668 400052 341674 400104
rect 338086 399996 345382 400024
rect 341518 399916 341524 399968
rect 341576 399956 341582 399968
rect 341576 399928 343726 399956
rect 341576 399916 341582 399928
rect 343698 399900 343726 399928
rect 343790 399928 344186 399956
rect 342346 399848 342352 399900
rect 342404 399888 342410 399900
rect 342576 399888 342582 399900
rect 342404 399860 342582 399888
rect 342404 399848 342410 399860
rect 342576 399848 342582 399860
rect 342634 399848 342640 399900
rect 342760 399848 342766 399900
rect 342818 399848 342824 399900
rect 343680 399848 343686 399900
rect 343738 399848 343744 399900
rect 340322 399712 340328 399764
rect 340380 399752 340386 399764
rect 342778 399752 342806 399848
rect 340380 399724 342806 399752
rect 340380 399712 340386 399724
rect 331916 399656 335354 399684
rect 331916 399644 331922 399656
rect 341242 399644 341248 399696
rect 341300 399684 341306 399696
rect 343790 399684 343818 399928
rect 344158 399900 344186 399928
rect 345354 399900 345382 399996
rect 344048 399848 344054 399900
rect 344106 399848 344112 399900
rect 344140 399848 344146 399900
rect 344198 399848 344204 399900
rect 344508 399848 344514 399900
rect 344566 399848 344572 399900
rect 344600 399848 344606 399900
rect 344658 399848 344664 399900
rect 344784 399848 344790 399900
rect 344842 399848 344848 399900
rect 345336 399848 345342 399900
rect 345394 399848 345400 399900
rect 346090 399888 346118 400132
rect 346228 399956 346256 400336
rect 346688 400228 346716 400404
rect 346688 400200 349798 400228
rect 347148 399996 348418 400024
rect 347148 399956 347176 399996
rect 346228 399928 347176 399956
rect 346164 399888 346170 399900
rect 346090 399860 346170 399888
rect 346164 399848 346170 399860
rect 346222 399848 346228 399900
rect 346348 399848 346354 399900
rect 346406 399848 346412 399900
rect 346716 399848 346722 399900
rect 346774 399848 346780 399900
rect 346992 399848 346998 399900
rect 347050 399848 347056 399900
rect 347176 399848 347182 399900
rect 347234 399848 347240 399900
rect 347360 399848 347366 399900
rect 347418 399848 347424 399900
rect 347820 399888 347826 399900
rect 347792 399848 347826 399888
rect 347878 399848 347884 399900
rect 347912 399848 347918 399900
rect 347970 399848 347976 399900
rect 348188 399848 348194 399900
rect 348246 399848 348252 399900
rect 348280 399848 348286 399900
rect 348338 399848 348344 399900
rect 341300 399656 343818 399684
rect 341300 399644 341306 399656
rect 310054 399576 310060 399628
rect 310112 399616 310118 399628
rect 341794 399616 341800 399628
rect 310112 399588 341800 399616
rect 310112 399576 310118 399588
rect 341794 399576 341800 399588
rect 341852 399576 341858 399628
rect 344066 399560 344094 399848
rect 344416 399780 344422 399832
rect 344474 399780 344480 399832
rect 344434 399696 344462 399780
rect 344370 399644 344376 399696
rect 344428 399656 344462 399696
rect 344428 399644 344434 399656
rect 344186 399576 344192 399628
rect 344244 399616 344250 399628
rect 344526 399616 344554 399848
rect 344618 399696 344646 399848
rect 344802 399764 344830 399848
rect 345980 399820 345986 399832
rect 344738 399712 344744 399764
rect 344796 399724 344830 399764
rect 345538 399792 345986 399820
rect 344796 399712 344802 399724
rect 344618 399656 344652 399696
rect 344646 399644 344652 399656
rect 344704 399644 344710 399696
rect 345538 399616 345566 399792
rect 345980 399780 345986 399792
rect 346038 399780 346044 399832
rect 346366 399684 346394 399848
rect 345998 399656 346394 399684
rect 345998 399628 346026 399656
rect 344244 399588 344554 399616
rect 345492 399588 345566 399616
rect 344244 399576 344250 399588
rect 311158 399508 311164 399560
rect 311216 399548 311222 399560
rect 342254 399548 342260 399560
rect 311216 399520 342260 399548
rect 311216 399508 311222 399520
rect 342254 399508 342260 399520
rect 342312 399508 342318 399560
rect 342806 399508 342812 399560
rect 342864 399548 342870 399560
rect 343818 399548 343824 399560
rect 342864 399520 343824 399548
rect 342864 399508 342870 399520
rect 343818 399508 343824 399520
rect 343876 399508 343882 399560
rect 344002 399508 344008 399560
rect 344060 399520 344094 399560
rect 344060 399508 344066 399520
rect 345290 399508 345296 399560
rect 345348 399548 345354 399560
rect 345492 399548 345520 399588
rect 345934 399576 345940 399628
rect 345992 399588 346026 399628
rect 346734 399616 346762 399848
rect 346090 399588 346762 399616
rect 345992 399576 345998 399588
rect 345348 399520 345520 399548
rect 345348 399508 345354 399520
rect 345566 399508 345572 399560
rect 345624 399548 345630 399560
rect 346090 399548 346118 399588
rect 347010 399548 347038 399848
rect 347194 399764 347222 399848
rect 347378 399764 347406 399848
rect 347544 399780 347550 399832
rect 347602 399780 347608 399832
rect 347636 399780 347642 399832
rect 347694 399780 347700 399832
rect 347194 399724 347228 399764
rect 347222 399712 347228 399724
rect 347280 399712 347286 399764
rect 347314 399712 347320 399764
rect 347372 399724 347406 399764
rect 347372 399712 347378 399724
rect 347562 399696 347590 399780
rect 347498 399644 347504 399696
rect 347556 399656 347590 399696
rect 347556 399644 347562 399656
rect 347654 399628 347682 399780
rect 347792 399764 347820 399848
rect 347774 399712 347780 399764
rect 347832 399712 347838 399764
rect 347930 399696 347958 399848
rect 348206 399820 348234 399848
rect 348160 399792 348234 399820
rect 348160 399696 348188 399792
rect 348298 399764 348326 399848
rect 348234 399712 348240 399764
rect 348292 399724 348326 399764
rect 348292 399712 348298 399724
rect 348390 399696 348418 399996
rect 349770 399956 349798 400200
rect 349862 400024 349890 400404
rect 357406 400092 357434 400472
rect 357406 400064 359642 400092
rect 349862 399996 357388 400024
rect 349770 399928 351914 399956
rect 351886 399900 351914 399928
rect 352438 399928 352696 399956
rect 352438 399900 352466 399928
rect 348832 399848 348838 399900
rect 348890 399848 348896 399900
rect 350580 399848 350586 399900
rect 350638 399848 350644 399900
rect 350672 399848 350678 399900
rect 350730 399888 350736 399900
rect 350730 399848 350764 399888
rect 350948 399848 350954 399900
rect 351006 399888 351012 399900
rect 351006 399848 351040 399888
rect 351408 399848 351414 399900
rect 351466 399888 351472 399900
rect 351466 399860 351592 399888
rect 351466 399848 351472 399860
rect 348740 399780 348746 399832
rect 348798 399780 348804 399832
rect 348758 399752 348786 399780
rect 347866 399644 347872 399696
rect 347924 399656 347958 399696
rect 347924 399644 347930 399656
rect 348142 399644 348148 399696
rect 348200 399644 348206 399696
rect 348326 399644 348332 399696
rect 348384 399656 348418 399696
rect 348712 399724 348786 399752
rect 348384 399644 348390 399656
rect 347590 399576 347596 399628
rect 347648 399588 347682 399628
rect 348712 399616 348740 399724
rect 348850 399696 348878 399848
rect 349016 399780 349022 399832
rect 349074 399820 349080 399832
rect 349476 399820 349482 399832
rect 349074 399780 349108 399820
rect 349080 399696 349108 399780
rect 349172 399792 349482 399820
rect 349172 399696 349200 399792
rect 349476 399780 349482 399792
rect 349534 399780 349540 399832
rect 349568 399780 349574 399832
rect 349626 399780 349632 399832
rect 349660 399780 349666 399832
rect 349718 399780 349724 399832
rect 349844 399780 349850 399832
rect 349902 399780 349908 399832
rect 349936 399780 349942 399832
rect 349994 399780 350000 399832
rect 350120 399780 350126 399832
rect 350178 399780 350184 399832
rect 350304 399780 350310 399832
rect 350362 399780 350368 399832
rect 350488 399820 350494 399832
rect 350460 399780 350494 399820
rect 350546 399780 350552 399832
rect 349586 399696 349614 399780
rect 348786 399644 348792 399696
rect 348844 399656 348878 399696
rect 348844 399644 348850 399656
rect 349062 399644 349068 399696
rect 349120 399644 349126 399696
rect 349154 399644 349160 399696
rect 349212 399644 349218 399696
rect 349522 399644 349528 399696
rect 349580 399656 349614 399696
rect 349580 399644 349586 399656
rect 348970 399616 348976 399628
rect 348712 399588 348976 399616
rect 347648 399576 347654 399588
rect 348970 399576 348976 399588
rect 349028 399576 349034 399628
rect 349430 399576 349436 399628
rect 349488 399616 349494 399628
rect 349678 399616 349706 399780
rect 349488 399588 349706 399616
rect 349488 399576 349494 399588
rect 349862 399560 349890 399780
rect 345624 399520 346118 399548
rect 346228 399520 347038 399548
rect 345624 399508 345630 399520
rect 312722 399440 312728 399492
rect 312780 399480 312786 399492
rect 312780 399452 344508 399480
rect 312780 399440 312786 399452
rect 277210 399372 277216 399424
rect 277268 399412 277274 399424
rect 344480 399412 344508 399452
rect 344554 399440 344560 399492
rect 344612 399480 344618 399492
rect 346228 399480 346256 399520
rect 347130 399508 347136 399560
rect 347188 399548 347194 399560
rect 348418 399548 348424 399560
rect 347188 399520 348424 399548
rect 347188 399508 347194 399520
rect 348418 399508 348424 399520
rect 348476 399508 348482 399560
rect 348510 399508 348516 399560
rect 348568 399508 348574 399560
rect 349798 399508 349804 399560
rect 349856 399520 349890 399560
rect 349856 399508 349862 399520
rect 344612 399452 346256 399480
rect 344612 399440 344618 399452
rect 346302 399440 346308 399492
rect 346360 399480 346366 399492
rect 348050 399480 348056 399492
rect 346360 399452 348056 399480
rect 346360 399440 346366 399452
rect 348050 399440 348056 399452
rect 348108 399440 348114 399492
rect 348528 399480 348556 399508
rect 349954 399492 349982 399780
rect 350138 399696 350166 399780
rect 350322 399752 350350 399780
rect 350322 399724 350396 399752
rect 350074 399644 350080 399696
rect 350132 399656 350166 399696
rect 350132 399644 350138 399656
rect 348160 399452 348556 399480
rect 346762 399412 346768 399424
rect 277268 399384 340874 399412
rect 344480 399384 346768 399412
rect 277268 399372 277274 399384
rect 275922 399304 275928 399356
rect 275980 399344 275986 399356
rect 340846 399344 340874 399384
rect 346762 399372 346768 399384
rect 346820 399372 346826 399424
rect 346946 399372 346952 399424
rect 347004 399412 347010 399424
rect 348160 399412 348188 399452
rect 349890 399440 349896 399492
rect 349948 399452 349982 399492
rect 349948 399440 349954 399452
rect 350258 399440 350264 399492
rect 350316 399480 350322 399492
rect 350368 399480 350396 399724
rect 350460 399628 350488 399780
rect 350598 399764 350626 399848
rect 350736 399764 350764 399848
rect 350598 399724 350632 399764
rect 350626 399712 350632 399724
rect 350684 399712 350690 399764
rect 350718 399712 350724 399764
rect 350776 399712 350782 399764
rect 351012 399628 351040 399848
rect 351224 399780 351230 399832
rect 351282 399780 351288 399832
rect 350442 399576 350448 399628
rect 350500 399576 350506 399628
rect 350994 399576 351000 399628
rect 351052 399576 351058 399628
rect 351242 399560 351270 399780
rect 351564 399684 351592 399860
rect 351684 399848 351690 399900
rect 351742 399848 351748 399900
rect 351868 399848 351874 399900
rect 351926 399848 351932 399900
rect 351960 399848 351966 399900
rect 352018 399848 352024 399900
rect 352236 399888 352242 399900
rect 352070 399860 352242 399888
rect 351702 399764 351730 399848
rect 351638 399712 351644 399764
rect 351696 399724 351730 399764
rect 351696 399712 351702 399724
rect 351730 399684 351736 399696
rect 351564 399656 351736 399684
rect 351730 399644 351736 399656
rect 351788 399644 351794 399696
rect 351978 399616 352006 399848
rect 352070 399696 352098 399860
rect 352236 399848 352242 399860
rect 352294 399848 352300 399900
rect 352420 399848 352426 399900
rect 352478 399848 352484 399900
rect 352512 399848 352518 399900
rect 352570 399888 352576 399900
rect 352570 399848 352604 399888
rect 352144 399780 352150 399832
rect 352202 399820 352208 399832
rect 352202 399792 352512 399820
rect 352202 399780 352208 399792
rect 352070 399656 352104 399696
rect 352098 399644 352104 399656
rect 352156 399644 352162 399696
rect 352190 399616 352196 399628
rect 351978 399588 352196 399616
rect 352190 399576 352196 399588
rect 352248 399576 352254 399628
rect 352374 399576 352380 399628
rect 352432 399616 352438 399628
rect 352484 399616 352512 399792
rect 352432 399588 352512 399616
rect 352432 399576 352438 399588
rect 351178 399508 351184 399560
rect 351236 399520 351270 399560
rect 351236 399508 351242 399520
rect 352006 399508 352012 399560
rect 352064 399548 352070 399560
rect 352576 399548 352604 399848
rect 352064 399520 352604 399548
rect 352064 399508 352070 399520
rect 350316 399452 350396 399480
rect 350316 399440 350322 399452
rect 352466 399440 352472 399492
rect 352524 399480 352530 399492
rect 352668 399480 352696 399928
rect 352760 399928 354674 399956
rect 352760 399560 352788 399928
rect 353248 399848 353254 399900
rect 353306 399888 353312 399900
rect 353616 399888 353622 399900
rect 353306 399848 353340 399888
rect 353312 399696 353340 399848
rect 353404 399860 353622 399888
rect 353294 399644 353300 399696
rect 353352 399644 353358 399696
rect 353404 399616 353432 399860
rect 353616 399848 353622 399860
rect 353674 399848 353680 399900
rect 353800 399848 353806 399900
rect 353858 399888 353864 399900
rect 354260 399888 354266 399900
rect 353858 399860 354030 399888
rect 353858 399848 353864 399860
rect 353892 399780 353898 399832
rect 353950 399780 353956 399832
rect 352944 399588 353432 399616
rect 352742 399508 352748 399560
rect 352800 399508 352806 399560
rect 352524 399452 352696 399480
rect 352524 399440 352530 399452
rect 349614 399412 349620 399424
rect 347004 399384 348188 399412
rect 348252 399384 349620 399412
rect 347004 399372 347010 399384
rect 348252 399344 348280 399384
rect 349614 399372 349620 399384
rect 349672 399372 349678 399424
rect 350902 399372 350908 399424
rect 350960 399412 350966 399424
rect 352944 399412 352972 399588
rect 353662 399576 353668 399628
rect 353720 399616 353726 399628
rect 353910 399616 353938 399780
rect 353720 399588 353938 399616
rect 353720 399576 353726 399588
rect 353846 399508 353852 399560
rect 353904 399548 353910 399560
rect 354002 399548 354030 399860
rect 354232 399848 354266 399888
rect 354318 399848 354324 399900
rect 354370 399860 354582 399888
rect 354076 399780 354082 399832
rect 354134 399820 354140 399832
rect 354134 399780 354168 399820
rect 354140 399560 354168 399780
rect 354232 399628 354260 399848
rect 354214 399576 354220 399628
rect 354272 399576 354278 399628
rect 353904 399520 354030 399548
rect 353904 399508 353910 399520
rect 354122 399508 354128 399560
rect 354180 399508 354186 399560
rect 353938 399440 353944 399492
rect 353996 399480 354002 399492
rect 354370 399480 354398 399860
rect 354444 399780 354450 399832
rect 354502 399780 354508 399832
rect 353996 399452 354398 399480
rect 353996 399440 354002 399452
rect 354462 399424 354490 399780
rect 354554 399616 354582 399860
rect 354646 399832 354674 399928
rect 355474 399928 355962 399956
rect 354720 399848 354726 399900
rect 354778 399848 354784 399900
rect 354904 399848 354910 399900
rect 354962 399848 354968 399900
rect 354628 399780 354634 399832
rect 354686 399780 354692 399832
rect 354738 399696 354766 399848
rect 354674 399644 354680 399696
rect 354732 399656 354766 399696
rect 354732 399644 354738 399656
rect 354922 399628 354950 399848
rect 355088 399780 355094 399832
rect 355146 399780 355152 399832
rect 354766 399616 354772 399628
rect 354554 399588 354772 399616
rect 354766 399576 354772 399588
rect 354824 399576 354830 399628
rect 354858 399576 354864 399628
rect 354916 399588 354950 399628
rect 354916 399576 354922 399588
rect 350960 399384 352972 399412
rect 350960 399372 350966 399384
rect 354398 399372 354404 399424
rect 354456 399384 354490 399424
rect 354456 399372 354462 399384
rect 354766 399372 354772 399424
rect 354824 399412 354830 399424
rect 355106 399412 355134 399780
rect 355474 399752 355502 399928
rect 355934 399900 355962 399928
rect 356164 399928 356606 399956
rect 355548 399848 355554 399900
rect 355606 399848 355612 399900
rect 355916 399848 355922 399900
rect 355974 399848 355980 399900
rect 355244 399724 355502 399752
rect 355244 399492 355272 399724
rect 355566 399696 355594 399848
rect 355502 399644 355508 399696
rect 355560 399656 355594 399696
rect 355560 399644 355566 399656
rect 355428 399588 356008 399616
rect 355428 399560 355456 399588
rect 355410 399508 355416 399560
rect 355468 399508 355474 399560
rect 355870 399548 355876 399560
rect 355520 399520 355876 399548
rect 355226 399440 355232 399492
rect 355284 399440 355290 399492
rect 354824 399384 355134 399412
rect 354824 399372 354830 399384
rect 354582 399344 354588 399356
rect 275980 399316 338114 399344
rect 340846 399316 348280 399344
rect 348344 399316 354588 399344
rect 275980 399304 275986 399316
rect 338086 399276 338114 399316
rect 348344 399276 348372 399316
rect 354582 399304 354588 399316
rect 354640 399304 354646 399356
rect 355134 399304 355140 399356
rect 355192 399344 355198 399356
rect 355520 399344 355548 399520
rect 355870 399508 355876 399520
rect 355928 399508 355934 399560
rect 355980 399480 356008 399588
rect 356164 399560 356192 399928
rect 356578 399900 356606 399928
rect 356284 399848 356290 399900
rect 356342 399888 356348 399900
rect 356342 399860 356514 399888
rect 356342 399848 356348 399860
rect 356486 399820 356514 399860
rect 356560 399848 356566 399900
rect 356618 399848 356624 399900
rect 356836 399848 356842 399900
rect 356894 399848 356900 399900
rect 357112 399848 357118 399900
rect 357170 399848 357176 399900
rect 356486 399792 356744 399820
rect 356606 399752 356612 399764
rect 356256 399724 356612 399752
rect 356146 399508 356152 399560
rect 356204 399508 356210 399560
rect 356256 399480 356284 399724
rect 356606 399712 356612 399724
rect 356664 399712 356670 399764
rect 356716 399616 356744 399792
rect 356440 399588 356744 399616
rect 356440 399548 356468 399588
rect 356348 399520 356468 399548
rect 356348 399492 356376 399520
rect 356514 399508 356520 399560
rect 356572 399548 356578 399560
rect 356854 399548 356882 399848
rect 356572 399520 356882 399548
rect 356572 399508 356578 399520
rect 355980 399452 356284 399480
rect 356330 399440 356336 399492
rect 356388 399440 356394 399492
rect 356422 399440 356428 399492
rect 356480 399480 356486 399492
rect 356790 399480 356796 399492
rect 356480 399452 356796 399480
rect 356480 399440 356486 399452
rect 356790 399440 356796 399452
rect 356848 399440 356854 399492
rect 355870 399372 355876 399424
rect 355928 399412 355934 399424
rect 357130 399412 357158 399848
rect 357360 399560 357388 399996
rect 357452 399928 358078 399956
rect 357342 399508 357348 399560
rect 357400 399508 357406 399560
rect 355928 399384 357158 399412
rect 355928 399372 355934 399384
rect 355192 399316 355548 399344
rect 355192 399304 355198 399316
rect 355686 399304 355692 399356
rect 355744 399344 355750 399356
rect 356238 399344 356244 399356
rect 355744 399316 356244 399344
rect 355744 399304 355750 399316
rect 356238 399304 356244 399316
rect 356296 399304 356302 399356
rect 356422 399304 356428 399356
rect 356480 399344 356486 399356
rect 357452 399344 357480 399928
rect 357572 399848 357578 399900
rect 357630 399848 357636 399900
rect 357756 399848 357762 399900
rect 357814 399848 357820 399900
rect 357848 399848 357854 399900
rect 357906 399848 357912 399900
rect 357940 399848 357946 399900
rect 357998 399848 358004 399900
rect 358050 399888 358078 399928
rect 359614 399900 359642 400064
rect 360948 399928 361574 399956
rect 358216 399888 358222 399900
rect 358050 399860 358222 399888
rect 358216 399848 358222 399860
rect 358274 399848 358280 399900
rect 358400 399848 358406 399900
rect 358458 399848 358464 399900
rect 358676 399848 358682 399900
rect 358734 399848 358740 399900
rect 358860 399848 358866 399900
rect 358918 399848 358924 399900
rect 359228 399848 359234 399900
rect 359286 399848 359292 399900
rect 359412 399848 359418 399900
rect 359470 399848 359476 399900
rect 359596 399848 359602 399900
rect 359654 399848 359660 399900
rect 360056 399848 360062 399900
rect 360114 399848 360120 399900
rect 360240 399848 360246 399900
rect 360298 399848 360304 399900
rect 360332 399848 360338 399900
rect 360390 399848 360396 399900
rect 360700 399848 360706 399900
rect 360758 399848 360764 399900
rect 360792 399848 360798 399900
rect 360850 399848 360856 399900
rect 357590 399560 357618 399848
rect 357590 399520 357624 399560
rect 357618 399508 357624 399520
rect 357676 399508 357682 399560
rect 356480 399316 357480 399344
rect 356480 399304 356486 399316
rect 338086 399248 348372 399276
rect 348418 399236 348424 399288
rect 348476 399276 348482 399288
rect 357158 399276 357164 399288
rect 348476 399248 357164 399276
rect 348476 399236 348482 399248
rect 357158 399236 357164 399248
rect 357216 399236 357222 399288
rect 357774 399276 357802 399848
rect 357866 399616 357894 399848
rect 357958 399696 357986 399848
rect 357958 399656 357992 399696
rect 357986 399644 357992 399656
rect 358044 399644 358050 399696
rect 358262 399644 358268 399696
rect 358320 399684 358326 399696
rect 358418 399684 358446 399848
rect 358492 399780 358498 399832
rect 358550 399780 358556 399832
rect 358320 399656 358446 399684
rect 358510 399696 358538 399780
rect 358510 399656 358544 399696
rect 358320 399644 358326 399656
rect 358538 399644 358544 399656
rect 358596 399644 358602 399696
rect 358446 399616 358452 399628
rect 357866 399588 358452 399616
rect 358446 399576 358452 399588
rect 358504 399576 358510 399628
rect 358170 399508 358176 399560
rect 358228 399548 358234 399560
rect 358694 399548 358722 399848
rect 358228 399520 358722 399548
rect 358228 399508 358234 399520
rect 358878 399480 358906 399848
rect 359136 399780 359142 399832
rect 359194 399780 359200 399832
rect 359154 399548 359182 399780
rect 359246 399628 359274 399848
rect 359246 399588 359280 399628
rect 359274 399576 359280 399588
rect 359332 399576 359338 399628
rect 359430 399616 359458 399848
rect 359688 399780 359694 399832
rect 359746 399780 359752 399832
rect 359780 399780 359786 399832
rect 359838 399780 359844 399832
rect 359872 399780 359878 399832
rect 359930 399780 359936 399832
rect 359706 399752 359734 399780
rect 359660 399724 359734 399752
rect 359660 399696 359688 399724
rect 359642 399644 359648 399696
rect 359700 399644 359706 399696
rect 359798 399684 359826 399780
rect 359752 399656 359826 399684
rect 359752 399628 359780 399656
rect 359890 399628 359918 399780
rect 359430 399588 359504 399616
rect 359476 399560 359504 399588
rect 359734 399576 359740 399628
rect 359792 399576 359798 399628
rect 359826 399576 359832 399628
rect 359884 399588 359918 399628
rect 359884 399576 359890 399588
rect 360074 399560 360102 399848
rect 360258 399684 360286 399848
rect 359366 399548 359372 399560
rect 359154 399520 359372 399548
rect 359366 399508 359372 399520
rect 359424 399508 359430 399560
rect 359458 399508 359464 399560
rect 359516 399508 359522 399560
rect 360010 399508 360016 399560
rect 360068 399520 360102 399560
rect 360212 399656 360286 399684
rect 360068 399508 360074 399520
rect 358878 399452 359136 399480
rect 359108 399424 359136 399452
rect 360102 399440 360108 399492
rect 360160 399480 360166 399492
rect 360212 399480 360240 399656
rect 360350 399628 360378 399848
rect 360286 399576 360292 399628
rect 360344 399588 360378 399628
rect 360344 399576 360350 399588
rect 360718 399492 360746 399848
rect 360160 399452 360240 399480
rect 360160 399440 360166 399452
rect 360654 399440 360660 399492
rect 360712 399452 360746 399492
rect 360810 399492 360838 399848
rect 360948 399560 360976 399928
rect 361546 399900 361574 399928
rect 361776 399928 362310 399956
rect 361068 399848 361074 399900
rect 361126 399848 361132 399900
rect 361160 399848 361166 399900
rect 361218 399848 361224 399900
rect 361252 399848 361258 399900
rect 361310 399848 361316 399900
rect 361528 399848 361534 399900
rect 361586 399848 361592 399900
rect 360930 399508 360936 399560
rect 360988 399508 360994 399560
rect 360810 399452 360844 399492
rect 360712 399440 360718 399452
rect 360838 399440 360844 399452
rect 360896 399440 360902 399492
rect 359090 399372 359096 399424
rect 359148 399372 359154 399424
rect 358722 399304 358728 399356
rect 358780 399344 358786 399356
rect 361086 399344 361114 399848
rect 358780 399316 361114 399344
rect 358780 399304 358786 399316
rect 358078 399276 358084 399288
rect 357774 399248 358084 399276
rect 358078 399236 358084 399248
rect 358136 399236 358142 399288
rect 360746 399236 360752 399288
rect 360804 399276 360810 399288
rect 361178 399276 361206 399848
rect 361270 399480 361298 399848
rect 361436 399780 361442 399832
rect 361494 399780 361500 399832
rect 361620 399780 361626 399832
rect 361678 399780 361684 399832
rect 361454 399560 361482 399780
rect 361638 399560 361666 399780
rect 361776 399560 361804 399928
rect 361896 399848 361902 399900
rect 361954 399848 361960 399900
rect 361390 399508 361396 399560
rect 361448 399520 361482 399560
rect 361448 399508 361454 399520
rect 361574 399508 361580 399560
rect 361632 399520 361666 399560
rect 361632 399508 361638 399520
rect 361758 399508 361764 399560
rect 361816 399508 361822 399560
rect 361914 399548 361942 399848
rect 362282 399832 362310 399928
rect 366146 399928 366404 399956
rect 366146 399900 366174 399928
rect 362724 399848 362730 399900
rect 362782 399848 362788 399900
rect 362908 399848 362914 399900
rect 362966 399888 362972 399900
rect 363092 399888 363098 399900
rect 362966 399848 363000 399888
rect 361988 399780 361994 399832
rect 362046 399780 362052 399832
rect 362264 399780 362270 399832
rect 362322 399780 362328 399832
rect 362356 399780 362362 399832
rect 362414 399780 362420 399832
rect 362448 399780 362454 399832
rect 362506 399780 362512 399832
rect 362006 399752 362034 399780
rect 362006 399724 362264 399752
rect 362126 399548 362132 399560
rect 361914 399520 362132 399548
rect 362126 399508 362132 399520
rect 362184 399508 362190 399560
rect 361482 399480 361488 399492
rect 361270 399452 361488 399480
rect 361482 399440 361488 399452
rect 361540 399440 361546 399492
rect 361666 399372 361672 399424
rect 361724 399412 361730 399424
rect 362236 399412 362264 399724
rect 362374 399696 362402 399780
rect 362310 399644 362316 399696
rect 362368 399656 362402 399696
rect 362368 399644 362374 399656
rect 362466 399628 362494 399780
rect 362586 399644 362592 399696
rect 362644 399684 362650 399696
rect 362742 399684 362770 399848
rect 362644 399656 362770 399684
rect 362644 399644 362650 399656
rect 362402 399576 362408 399628
rect 362460 399588 362494 399628
rect 362460 399576 362466 399588
rect 362494 399508 362500 399560
rect 362552 399548 362558 399560
rect 362972 399548 363000 399848
rect 363064 399848 363098 399888
rect 363150 399848 363156 399900
rect 363552 399848 363558 399900
rect 363610 399848 363616 399900
rect 363644 399848 363650 399900
rect 363702 399848 363708 399900
rect 364012 399848 364018 399900
rect 364070 399848 364076 399900
rect 364288 399848 364294 399900
rect 364346 399848 364352 399900
rect 364380 399848 364386 399900
rect 364438 399848 364444 399900
rect 364564 399848 364570 399900
rect 364622 399848 364628 399900
rect 365024 399848 365030 399900
rect 365082 399848 365088 399900
rect 365208 399888 365214 399900
rect 365180 399848 365214 399888
rect 365266 399848 365272 399900
rect 365300 399848 365306 399900
rect 365358 399848 365364 399900
rect 365484 399848 365490 399900
rect 365542 399848 365548 399900
rect 366036 399848 366042 399900
rect 366094 399848 366100 399900
rect 366128 399848 366134 399900
rect 366186 399848 366192 399900
rect 366220 399848 366226 399900
rect 366278 399848 366284 399900
rect 363064 399560 363092 399848
rect 362552 399520 363000 399548
rect 362552 399508 362558 399520
rect 363046 399508 363052 399560
rect 363104 399508 363110 399560
rect 363570 399480 363598 399848
rect 363248 399452 363598 399480
rect 363248 399424 363276 399452
rect 361724 399384 362264 399412
rect 361724 399372 361730 399384
rect 363230 399372 363236 399424
rect 363288 399372 363294 399424
rect 363322 399372 363328 399424
rect 363380 399412 363386 399424
rect 363662 399412 363690 399848
rect 364030 399820 364058 399848
rect 363984 399792 364058 399820
rect 363984 399696 364012 399792
rect 363966 399644 363972 399696
rect 364024 399644 364030 399696
rect 364306 399628 364334 399848
rect 364398 399696 364426 399848
rect 364398 399656 364432 399696
rect 364426 399644 364432 399656
rect 364484 399644 364490 399696
rect 364306 399588 364340 399628
rect 364334 399576 364340 399588
rect 364392 399576 364398 399628
rect 364058 399508 364064 399560
rect 364116 399548 364122 399560
rect 364582 399548 364610 399848
rect 364748 399780 364754 399832
rect 364806 399780 364812 399832
rect 364116 399520 364610 399548
rect 364116 399508 364122 399520
rect 363380 399384 363690 399412
rect 363380 399372 363386 399384
rect 361298 399304 361304 399356
rect 361356 399344 361362 399356
rect 364766 399344 364794 399780
rect 364886 399508 364892 399560
rect 364944 399548 364950 399560
rect 365042 399548 365070 399848
rect 365180 399696 365208 399848
rect 365318 399764 365346 399848
rect 365254 399712 365260 399764
rect 365312 399724 365346 399764
rect 365312 399712 365318 399724
rect 365502 399696 365530 399848
rect 365162 399644 365168 399696
rect 365220 399644 365226 399696
rect 365438 399644 365444 399696
rect 365496 399656 365530 399696
rect 365496 399644 365502 399656
rect 366054 399628 366082 399848
rect 365530 399576 365536 399628
rect 365588 399616 365594 399628
rect 365588 399588 365760 399616
rect 366054 399588 366088 399628
rect 365588 399576 365594 399588
rect 365732 399560 365760 399588
rect 366082 399576 366088 399588
rect 366140 399576 366146 399628
rect 364944 399520 365070 399548
rect 364944 399508 364950 399520
rect 365714 399508 365720 399560
rect 365772 399508 365778 399560
rect 365806 399508 365812 399560
rect 365864 399548 365870 399560
rect 366238 399548 366266 399848
rect 366376 399696 366404 399928
rect 366468 399820 366496 400608
rect 387794 400460 387800 400512
rect 387852 400500 387858 400512
rect 392118 400500 392124 400512
rect 387852 400472 392124 400500
rect 387852 400460 387858 400472
rect 392118 400460 392124 400472
rect 392176 400460 392182 400512
rect 390186 400324 390192 400376
rect 390244 400364 390250 400376
rect 394786 400364 394792 400376
rect 390244 400336 394792 400364
rect 390244 400324 390250 400336
rect 394786 400324 394792 400336
rect 394844 400324 394850 400376
rect 387886 400092 387892 400104
rect 384178 400064 387892 400092
rect 366606 399928 367048 399956
rect 366606 399900 366634 399928
rect 366588 399848 366594 399900
rect 366646 399848 366652 399900
rect 366864 399848 366870 399900
rect 366922 399888 366928 399900
rect 366922 399848 366956 399888
rect 366468 399792 366864 399820
rect 366836 399764 366864 399792
rect 366542 399712 366548 399764
rect 366600 399712 366606 399764
rect 366726 399752 366732 399764
rect 366652 399724 366732 399752
rect 366358 399644 366364 399696
rect 366416 399644 366422 399696
rect 365864 399520 366266 399548
rect 365864 399508 365870 399520
rect 366450 399508 366456 399560
rect 366508 399548 366514 399560
rect 366560 399548 366588 399712
rect 366652 399628 366680 399724
rect 366726 399712 366732 399724
rect 366784 399712 366790 399764
rect 366818 399712 366824 399764
rect 366876 399712 366882 399764
rect 366634 399576 366640 399628
rect 366692 399576 366698 399628
rect 366508 399520 366588 399548
rect 366508 399508 366514 399520
rect 366726 399508 366732 399560
rect 366784 399548 366790 399560
rect 366928 399548 366956 399848
rect 366784 399520 366956 399548
rect 366784 399508 366790 399520
rect 366542 399440 366548 399492
rect 366600 399480 366606 399492
rect 367020 399480 367048 399928
rect 371804 399928 372890 399956
rect 367600 399848 367606 399900
rect 367658 399848 367664 399900
rect 368704 399848 368710 399900
rect 368762 399848 368768 399900
rect 368796 399848 368802 399900
rect 368854 399848 368860 399900
rect 369164 399848 369170 399900
rect 369222 399848 369228 399900
rect 369900 399848 369906 399900
rect 369958 399848 369964 399900
rect 370084 399848 370090 399900
rect 370142 399848 370148 399900
rect 370360 399848 370366 399900
rect 370418 399848 370424 399900
rect 370728 399848 370734 399900
rect 370786 399848 370792 399900
rect 370912 399848 370918 399900
rect 370970 399848 370976 399900
rect 371280 399848 371286 399900
rect 371338 399888 371344 399900
rect 371338 399848 371372 399888
rect 371648 399848 371654 399900
rect 371706 399848 371712 399900
rect 367416 399780 367422 399832
rect 367474 399780 367480 399832
rect 367434 399696 367462 399780
rect 367434 399656 367468 399696
rect 367462 399644 367468 399656
rect 367520 399644 367526 399696
rect 367618 399616 367646 399848
rect 368244 399780 368250 399832
rect 368302 399780 368308 399832
rect 368336 399780 368342 399832
rect 368394 399780 368400 399832
rect 368262 399628 368290 399780
rect 367922 399616 367928 399628
rect 367618 399588 367928 399616
rect 367922 399576 367928 399588
rect 367980 399576 367986 399628
rect 368198 399576 368204 399628
rect 368256 399588 368290 399628
rect 368256 399576 368262 399588
rect 368354 399560 368382 399780
rect 368722 399696 368750 399848
rect 368658 399644 368664 399696
rect 368716 399656 368750 399696
rect 368716 399644 368722 399656
rect 368814 399616 368842 399848
rect 368814 399588 368980 399616
rect 368952 399560 368980 399588
rect 368290 399508 368296 399560
rect 368348 399520 368382 399560
rect 368348 399508 368354 399520
rect 368934 399508 368940 399560
rect 368992 399508 368998 399560
rect 369182 399548 369210 399848
rect 369044 399520 369210 399548
rect 366600 399452 367048 399480
rect 366600 399440 366606 399452
rect 367370 399372 367376 399424
rect 367428 399412 367434 399424
rect 367554 399412 367560 399424
rect 367428 399384 367560 399412
rect 367428 399372 367434 399384
rect 367554 399372 367560 399384
rect 367612 399372 367618 399424
rect 361356 399316 364794 399344
rect 361356 399304 361362 399316
rect 360804 399248 361206 399276
rect 360804 399236 360810 399248
rect 364058 399236 364064 399288
rect 364116 399276 364122 399288
rect 367554 399276 367560 399288
rect 364116 399248 367560 399276
rect 364116 399236 364122 399248
rect 367554 399236 367560 399248
rect 367612 399236 367618 399288
rect 367664 399248 367922 399276
rect 337746 399168 337752 399220
rect 337804 399208 337810 399220
rect 348694 399208 348700 399220
rect 337804 399180 348700 399208
rect 337804 399168 337810 399180
rect 348694 399168 348700 399180
rect 348752 399168 348758 399220
rect 349614 399168 349620 399220
rect 349672 399208 349678 399220
rect 353478 399208 353484 399220
rect 349672 399180 353484 399208
rect 349672 399168 349678 399180
rect 353478 399168 353484 399180
rect 353536 399168 353542 399220
rect 354030 399168 354036 399220
rect 354088 399208 354094 399220
rect 367664 399208 367692 399248
rect 354088 399180 367692 399208
rect 367894 399208 367922 399248
rect 368382 399236 368388 399288
rect 368440 399276 368446 399288
rect 369044 399276 369072 399520
rect 369670 399372 369676 399424
rect 369728 399412 369734 399424
rect 369918 399412 369946 399848
rect 369992 399780 369998 399832
rect 370050 399780 370056 399832
rect 370010 399560 370038 399780
rect 370102 399616 370130 399848
rect 370102 399588 370176 399616
rect 370010 399520 370044 399560
rect 370038 399508 370044 399520
rect 370096 399508 370102 399560
rect 369728 399384 369946 399412
rect 369728 399372 369734 399384
rect 369578 399304 369584 399356
rect 369636 399344 369642 399356
rect 370148 399344 370176 399588
rect 370222 399440 370228 399492
rect 370280 399480 370286 399492
rect 370378 399480 370406 399848
rect 370544 399780 370550 399832
rect 370602 399780 370608 399832
rect 370562 399628 370590 399780
rect 370746 399684 370774 399848
rect 370746 399656 370820 399684
rect 370498 399576 370504 399628
rect 370556 399588 370590 399628
rect 370556 399576 370562 399588
rect 370682 399576 370688 399628
rect 370740 399576 370746 399628
rect 370280 399452 370406 399480
rect 370280 399440 370286 399452
rect 370590 399440 370596 399492
rect 370648 399480 370654 399492
rect 370700 399480 370728 399576
rect 370648 399452 370728 399480
rect 370648 399440 370654 399452
rect 370682 399372 370688 399424
rect 370740 399412 370746 399424
rect 370792 399412 370820 399656
rect 370930 399560 370958 399848
rect 371344 399764 371372 399848
rect 371666 399764 371694 399848
rect 371326 399712 371332 399764
rect 371384 399712 371390 399764
rect 371666 399724 371700 399764
rect 371694 399712 371700 399724
rect 371752 399712 371758 399764
rect 370930 399520 370964 399560
rect 370958 399508 370964 399520
rect 371016 399508 371022 399560
rect 370740 399384 370820 399412
rect 370740 399372 370746 399384
rect 371050 399372 371056 399424
rect 371108 399412 371114 399424
rect 371804 399412 371832 399928
rect 372862 399900 372890 399928
rect 374426 399928 374960 399956
rect 374426 399900 374454 399928
rect 372016 399888 372022 399900
rect 371108 399384 371832 399412
rect 371896 399860 372022 399888
rect 371108 399372 371114 399384
rect 369636 399316 370176 399344
rect 369636 399304 369642 399316
rect 371510 399304 371516 399356
rect 371568 399344 371574 399356
rect 371896 399344 371924 399860
rect 372016 399848 372022 399860
rect 372074 399848 372080 399900
rect 372108 399848 372114 399900
rect 372166 399848 372172 399900
rect 372292 399848 372298 399900
rect 372350 399848 372356 399900
rect 372660 399848 372666 399900
rect 372718 399888 372724 399900
rect 372718 399848 372752 399888
rect 372844 399848 372850 399900
rect 372902 399848 372908 399900
rect 373028 399848 373034 399900
rect 373086 399848 373092 399900
rect 373212 399848 373218 399900
rect 373270 399888 373276 399900
rect 373270 399860 374040 399888
rect 373270 399848 373276 399860
rect 372126 399616 372154 399848
rect 372310 399696 372338 399848
rect 372476 399820 372482 399832
rect 372448 399780 372482 399820
rect 372534 399780 372540 399832
rect 372448 399696 372476 399780
rect 372310 399656 372344 399696
rect 372338 399644 372344 399656
rect 372396 399644 372402 399696
rect 372430 399644 372436 399696
rect 372488 399644 372494 399696
rect 372522 399616 372528 399628
rect 372126 399588 372528 399616
rect 372522 399576 372528 399588
rect 372580 399576 372586 399628
rect 371970 399508 371976 399560
rect 372028 399548 372034 399560
rect 372724 399548 372752 399848
rect 372798 399644 372804 399696
rect 372856 399684 372862 399696
rect 373046 399684 373074 399848
rect 373488 399820 373494 399832
rect 372856 399656 373074 399684
rect 373460 399780 373494 399820
rect 373546 399780 373552 399832
rect 373580 399780 373586 399832
rect 373638 399780 373644 399832
rect 373672 399780 373678 399832
rect 373730 399780 373736 399832
rect 373764 399780 373770 399832
rect 373822 399780 373828 399832
rect 373856 399780 373862 399832
rect 373914 399780 373920 399832
rect 372856 399644 372862 399656
rect 373460 399560 373488 399780
rect 373598 399752 373626 399780
rect 373552 399724 373626 399752
rect 373552 399628 373580 399724
rect 373690 399684 373718 399780
rect 373644 399656 373718 399684
rect 373534 399576 373540 399628
rect 373592 399576 373598 399628
rect 372028 399520 372752 399548
rect 372028 399508 372034 399520
rect 373442 399508 373448 399560
rect 373500 399508 373506 399560
rect 373644 399492 373672 399656
rect 373782 399628 373810 399780
rect 373874 399696 373902 399780
rect 373874 399656 373908 399696
rect 373902 399644 373908 399656
rect 373960 399644 373966 399696
rect 373718 399576 373724 399628
rect 373776 399588 373810 399628
rect 374012 399616 374040 399860
rect 374224 399848 374230 399900
rect 374282 399848 374288 399900
rect 374408 399848 374414 399900
rect 374466 399848 374472 399900
rect 374684 399848 374690 399900
rect 374742 399848 374748 399900
rect 373874 399588 374040 399616
rect 374242 399628 374270 399848
rect 374592 399780 374598 399832
rect 374650 399780 374656 399832
rect 374242 399588 374276 399628
rect 373776 399576 373782 399588
rect 373874 399560 373902 399588
rect 374270 399576 374276 399588
rect 374328 399576 374334 399628
rect 373810 399508 373816 399560
rect 373868 399520 373902 399560
rect 374454 399548 374460 399560
rect 374104 399520 374460 399548
rect 373868 399508 373874 399520
rect 374104 399492 374132 399520
rect 374454 399508 374460 399520
rect 374512 399508 374518 399560
rect 373626 399440 373632 399492
rect 373684 399440 373690 399492
rect 374086 399440 374092 399492
rect 374144 399440 374150 399492
rect 374610 399480 374638 399780
rect 374702 399548 374730 399848
rect 374776 399780 374782 399832
rect 374834 399780 374840 399832
rect 374794 399628 374822 399780
rect 374794 399588 374828 399628
rect 374822 399576 374828 399588
rect 374880 399576 374886 399628
rect 374702 399520 374868 399548
rect 374730 399480 374736 399492
rect 374610 399452 374736 399480
rect 374730 399440 374736 399452
rect 374788 399440 374794 399492
rect 374454 399372 374460 399424
rect 374512 399412 374518 399424
rect 374840 399412 374868 399520
rect 374932 399492 374960 399928
rect 378198 399928 379054 399956
rect 378198 399900 378226 399928
rect 375236 399848 375242 399900
rect 375294 399888 375300 399900
rect 375294 399848 375328 399888
rect 375880 399848 375886 399900
rect 375938 399848 375944 399900
rect 376064 399848 376070 399900
rect 376122 399848 376128 399900
rect 376340 399848 376346 399900
rect 376398 399848 376404 399900
rect 376432 399848 376438 399900
rect 376490 399848 376496 399900
rect 376800 399848 376806 399900
rect 376858 399848 376864 399900
rect 377720 399888 377726 399900
rect 377692 399848 377726 399888
rect 377778 399848 377784 399900
rect 377812 399848 377818 399900
rect 377870 399848 377876 399900
rect 378180 399848 378186 399900
rect 378238 399848 378244 399900
rect 378272 399848 378278 399900
rect 378330 399848 378336 399900
rect 378916 399848 378922 399900
rect 378974 399848 378980 399900
rect 375052 399780 375058 399832
rect 375110 399780 375116 399832
rect 375144 399780 375150 399832
rect 375202 399820 375208 399832
rect 375202 399780 375236 399820
rect 375070 399628 375098 399780
rect 375208 399696 375236 399780
rect 375190 399644 375196 399696
rect 375248 399644 375254 399696
rect 375070 399588 375104 399628
rect 375098 399576 375104 399588
rect 375156 399576 375162 399628
rect 375190 399508 375196 399560
rect 375248 399548 375254 399560
rect 375300 399548 375328 399848
rect 375604 399780 375610 399832
rect 375662 399780 375668 399832
rect 375248 399520 375328 399548
rect 375248 399508 375254 399520
rect 374914 399440 374920 399492
rect 374972 399440 374978 399492
rect 375374 399440 375380 399492
rect 375432 399480 375438 399492
rect 375622 399480 375650 399780
rect 375742 399508 375748 399560
rect 375800 399548 375806 399560
rect 375898 399548 375926 399848
rect 375800 399520 375926 399548
rect 375800 399508 375806 399520
rect 375432 399452 375650 399480
rect 375432 399440 375438 399452
rect 374512 399384 374868 399412
rect 374512 399372 374518 399384
rect 371568 399316 371924 399344
rect 371568 399304 371574 399316
rect 368440 399248 369072 399276
rect 376082 399276 376110 399848
rect 376202 399576 376208 399628
rect 376260 399616 376266 399628
rect 376358 399616 376386 399848
rect 376260 399588 376386 399616
rect 376260 399576 376266 399588
rect 376450 399560 376478 399848
rect 376818 399684 376846 399848
rect 377076 399780 377082 399832
rect 377134 399780 377140 399832
rect 377168 399780 377174 399832
rect 377226 399780 377232 399832
rect 377352 399780 377358 399832
rect 377410 399780 377416 399832
rect 377444 399780 377450 399832
rect 377502 399780 377508 399832
rect 377094 399696 377122 399780
rect 376938 399684 376944 399696
rect 376818 399656 376944 399684
rect 376938 399644 376944 399656
rect 376996 399644 377002 399696
rect 377030 399644 377036 399696
rect 377088 399656 377122 399696
rect 377088 399644 377094 399656
rect 376386 399508 376392 399560
rect 376444 399520 376478 399560
rect 376444 399508 376450 399520
rect 376294 399276 376300 399288
rect 376082 399248 376300 399276
rect 368440 399236 368446 399248
rect 376294 399236 376300 399248
rect 376352 399236 376358 399288
rect 377186 399276 377214 399780
rect 377370 399696 377398 399780
rect 377306 399644 377312 399696
rect 377364 399656 377398 399696
rect 377364 399644 377370 399656
rect 377462 399560 377490 399780
rect 377692 399764 377720 399848
rect 377830 399820 377858 399848
rect 377784 399792 377858 399820
rect 377784 399764 377812 399792
rect 377674 399712 377680 399764
rect 377732 399712 377738 399764
rect 377766 399712 377772 399764
rect 377824 399712 377830 399764
rect 378290 399752 378318 399848
rect 378290 399724 378640 399752
rect 378612 399560 378640 399724
rect 377398 399508 377404 399560
rect 377456 399520 377490 399560
rect 377456 399508 377462 399520
rect 378594 399508 378600 399560
rect 378652 399508 378658 399560
rect 378594 399372 378600 399424
rect 378652 399412 378658 399424
rect 378934 399412 378962 399848
rect 379026 399548 379054 399928
rect 384178 399900 384206 400064
rect 387886 400052 387892 400064
rect 387944 400052 387950 400104
rect 387978 400024 387984 400036
rect 385558 399996 387984 400024
rect 384270 399928 385494 399956
rect 384270 399900 384298 399928
rect 379100 399848 379106 399900
rect 379158 399848 379164 399900
rect 379376 399848 379382 399900
rect 379434 399848 379440 399900
rect 379744 399888 379750 399900
rect 379716 399848 379750 399888
rect 379802 399848 379808 399900
rect 380296 399848 380302 399900
rect 380354 399848 380360 399900
rect 380664 399848 380670 399900
rect 380722 399848 380728 399900
rect 381216 399848 381222 399900
rect 381274 399848 381280 399900
rect 381492 399848 381498 399900
rect 381550 399848 381556 399900
rect 381584 399848 381590 399900
rect 381642 399848 381648 399900
rect 381952 399848 381958 399900
rect 382010 399848 382016 399900
rect 382228 399848 382234 399900
rect 382286 399848 382292 399900
rect 382596 399848 382602 399900
rect 382654 399848 382660 399900
rect 382780 399848 382786 399900
rect 382838 399848 382844 399900
rect 383424 399848 383430 399900
rect 383482 399848 383488 399900
rect 383700 399888 383706 399900
rect 383672 399848 383706 399888
rect 383758 399848 383764 399900
rect 383792 399848 383798 399900
rect 383850 399848 383856 399900
rect 384160 399848 384166 399900
rect 384218 399848 384224 399900
rect 384252 399848 384258 399900
rect 384310 399848 384316 399900
rect 384436 399848 384442 399900
rect 384494 399848 384500 399900
rect 379118 399684 379146 399848
rect 379394 399764 379422 399848
rect 379716 399764 379744 399848
rect 379330 399712 379336 399764
rect 379388 399724 379422 399764
rect 379388 399712 379394 399724
rect 379698 399712 379704 399764
rect 379756 399712 379762 399764
rect 379974 399712 379980 399764
rect 380032 399712 380038 399764
rect 379422 399684 379428 399696
rect 379118 399656 379428 399684
rect 379422 399644 379428 399656
rect 379480 399644 379486 399696
rect 379606 399644 379612 399696
rect 379664 399684 379670 399696
rect 379992 399684 380020 399712
rect 379664 399656 380020 399684
rect 379664 399644 379670 399656
rect 379146 399548 379152 399560
rect 379026 399520 379152 399548
rect 379146 399508 379152 399520
rect 379204 399508 379210 399560
rect 379790 399548 379796 399560
rect 379532 399520 379796 399548
rect 378652 399384 378962 399412
rect 379532 399412 379560 399520
rect 379790 399508 379796 399520
rect 379848 399508 379854 399560
rect 380314 399492 380342 399848
rect 380480 399780 380486 399832
rect 380538 399780 380544 399832
rect 380498 399696 380526 399780
rect 380498 399656 380532 399696
rect 380526 399644 380532 399656
rect 380584 399644 380590 399696
rect 380434 399576 380440 399628
rect 380492 399616 380498 399628
rect 380682 399616 380710 399848
rect 380492 399588 380710 399616
rect 380492 399576 380498 399588
rect 380894 399508 380900 399560
rect 380952 399548 380958 399560
rect 381234 399548 381262 399848
rect 381354 399576 381360 399628
rect 381412 399616 381418 399628
rect 381510 399616 381538 399848
rect 381412 399588 381538 399616
rect 381412 399576 381418 399588
rect 381602 399560 381630 399848
rect 381970 399560 381998 399848
rect 380952 399520 381262 399548
rect 380952 399508 380958 399520
rect 381538 399508 381544 399560
rect 381596 399520 381630 399560
rect 381596 399508 381602 399520
rect 381906 399508 381912 399560
rect 381964 399520 381998 399560
rect 382246 399548 382274 399848
rect 382614 399764 382642 399848
rect 382614 399724 382648 399764
rect 382642 399712 382648 399724
rect 382700 399712 382706 399764
rect 382798 399616 382826 399848
rect 383442 399752 383470 399848
rect 383442 399724 383608 399752
rect 383580 399696 383608 399724
rect 383562 399644 383568 399696
rect 383620 399644 383626 399696
rect 383672 399616 383700 399848
rect 383810 399684 383838 399848
rect 383930 399684 383936 399696
rect 383810 399656 383936 399684
rect 383930 399644 383936 399656
rect 383988 399644 383994 399696
rect 384298 399644 384304 399696
rect 384356 399684 384362 399696
rect 384454 399684 384482 399848
rect 385080 399780 385086 399832
rect 385138 399780 385144 399832
rect 384712 399712 384718 399764
rect 384770 399712 384776 399764
rect 384356 399656 384482 399684
rect 384356 399644 384362 399656
rect 382798 399588 383332 399616
rect 383672 399588 384528 399616
rect 383304 399560 383332 399588
rect 382366 399548 382372 399560
rect 382246 399520 382372 399548
rect 381964 399508 381970 399520
rect 382366 399508 382372 399520
rect 382424 399508 382430 399560
rect 383286 399508 383292 399560
rect 383344 399508 383350 399560
rect 380250 399440 380256 399492
rect 380308 399452 380342 399492
rect 384500 399480 384528 399588
rect 384574 399508 384580 399560
rect 384632 399548 384638 399560
rect 384730 399548 384758 399712
rect 384632 399520 384758 399548
rect 384632 399508 384638 399520
rect 384758 399480 384764 399492
rect 384500 399452 384764 399480
rect 380308 399440 380314 399452
rect 384758 399440 384764 399452
rect 384816 399440 384822 399492
rect 385098 399480 385126 399780
rect 385466 399548 385494 399928
rect 385558 399900 385586 399996
rect 387978 399984 387984 399996
rect 388036 399984 388042 400036
rect 390186 399956 390192 399968
rect 387030 399928 390192 399956
rect 387030 399900 387058 399928
rect 390186 399916 390192 399928
rect 390244 399916 390250 399968
rect 385540 399848 385546 399900
rect 385598 399848 385604 399900
rect 385908 399848 385914 399900
rect 385966 399848 385972 399900
rect 386000 399848 386006 399900
rect 386058 399848 386064 399900
rect 386552 399848 386558 399900
rect 386610 399848 386616 399900
rect 387012 399848 387018 399900
rect 387070 399848 387076 399900
rect 387196 399848 387202 399900
rect 387254 399888 387260 399900
rect 387518 399888 387524 399900
rect 387254 399860 387524 399888
rect 387254 399848 387260 399860
rect 387518 399848 387524 399860
rect 387576 399848 387582 399900
rect 385632 399780 385638 399832
rect 385690 399780 385696 399832
rect 385650 399696 385678 399780
rect 385926 399696 385954 399848
rect 385650 399656 385684 399696
rect 385678 399644 385684 399656
rect 385736 399644 385742 399696
rect 385862 399644 385868 399696
rect 385920 399656 385954 399696
rect 385920 399644 385926 399656
rect 385770 399576 385776 399628
rect 385828 399616 385834 399628
rect 386018 399616 386046 399848
rect 386184 399780 386190 399832
rect 386242 399780 386248 399832
rect 385828 399588 386046 399616
rect 386202 399628 386230 399780
rect 386202 399588 386236 399628
rect 385828 399576 385834 399588
rect 386230 399576 386236 399588
rect 386288 399576 386294 399628
rect 386414 399576 386420 399628
rect 386472 399616 386478 399628
rect 386570 399616 386598 399848
rect 386736 399780 386742 399832
rect 386794 399780 386800 399832
rect 387104 399780 387110 399832
rect 387162 399780 387168 399832
rect 386754 399752 386782 399780
rect 386472 399588 386598 399616
rect 386708 399724 386782 399752
rect 386708 399616 386736 399724
rect 386782 399644 386788 399696
rect 386840 399684 386846 399696
rect 387122 399684 387150 399780
rect 386840 399656 387150 399684
rect 386840 399644 386846 399656
rect 386874 399616 386880 399628
rect 386708 399588 386880 399616
rect 386472 399576 386478 399588
rect 386874 399576 386880 399588
rect 386932 399576 386938 399628
rect 389174 399548 389180 399560
rect 385466 399520 389180 399548
rect 389174 399508 389180 399520
rect 389232 399508 389238 399560
rect 385586 399480 385592 399492
rect 385098 399452 385592 399480
rect 385586 399440 385592 399452
rect 385644 399440 385650 399492
rect 387794 399412 387800 399424
rect 379532 399384 387800 399412
rect 378652 399372 378658 399384
rect 387794 399372 387800 399384
rect 387852 399372 387858 399424
rect 378686 399304 378692 399356
rect 378744 399344 378750 399356
rect 379238 399344 379244 399356
rect 378744 399316 379244 399344
rect 378744 399304 378750 399316
rect 379238 399304 379244 399316
rect 379296 399304 379302 399356
rect 377674 399276 377680 399288
rect 377186 399248 377680 399276
rect 377674 399236 377680 399248
rect 377732 399236 377738 399288
rect 379606 399208 379612 399220
rect 367894 399180 379612 399208
rect 354088 399168 354094 399180
rect 379606 399168 379612 399180
rect 379664 399168 379670 399220
rect 338022 399100 338028 399152
rect 338080 399140 338086 399152
rect 366174 399140 366180 399152
rect 338080 399112 366180 399140
rect 338080 399100 338086 399112
rect 366174 399100 366180 399112
rect 366232 399100 366238 399152
rect 379238 399140 379244 399152
rect 371436 399112 379244 399140
rect 334986 399032 334992 399084
rect 335044 399072 335050 399084
rect 335044 399044 348694 399072
rect 335044 399032 335050 399044
rect 278682 398964 278688 399016
rect 278740 399004 278746 399016
rect 348510 399004 348516 399016
rect 278740 398976 348516 399004
rect 278740 398964 278746 398976
rect 348510 398964 348516 398976
rect 348568 398964 348574 399016
rect 348666 399004 348694 399044
rect 348758 399044 360194 399072
rect 348758 399004 348786 399044
rect 348666 398976 348786 399004
rect 349982 398964 349988 399016
rect 350040 399004 350046 399016
rect 360166 399004 360194 399044
rect 362862 399032 362868 399084
rect 362920 399072 362926 399084
rect 364518 399072 364524 399084
rect 362920 399044 364524 399072
rect 362920 399032 362926 399044
rect 364518 399032 364524 399044
rect 364576 399032 364582 399084
rect 371436 399072 371464 399112
rect 379238 399100 379244 399112
rect 379296 399100 379302 399152
rect 381630 399100 381636 399152
rect 381688 399140 381694 399152
rect 381906 399140 381912 399152
rect 381688 399112 381912 399140
rect 381688 399100 381694 399112
rect 381906 399100 381912 399112
rect 381964 399100 381970 399152
rect 365686 399044 371464 399072
rect 365686 399004 365714 399044
rect 350040 398976 358814 399004
rect 360166 398976 365714 399004
rect 350040 398964 350046 398976
rect 340506 398896 340512 398948
rect 340564 398936 340570 398948
rect 355962 398936 355968 398948
rect 340564 398908 355968 398936
rect 340564 398896 340570 398908
rect 355962 398896 355968 398908
rect 356020 398896 356026 398948
rect 356146 398896 356152 398948
rect 356204 398936 356210 398948
rect 356514 398936 356520 398948
rect 356204 398908 356520 398936
rect 356204 398896 356210 398908
rect 356514 398896 356520 398908
rect 356572 398896 356578 398948
rect 358786 398936 358814 398976
rect 366174 398964 366180 399016
rect 366232 399004 366238 399016
rect 366232 398976 376754 399004
rect 366232 398964 366238 398976
rect 365898 398936 365904 398948
rect 358786 398908 365904 398936
rect 365898 398896 365904 398908
rect 365956 398896 365962 398948
rect 375742 398936 375748 398948
rect 375484 398908 375748 398936
rect 375484 398880 375512 398908
rect 375742 398896 375748 398908
rect 375800 398896 375806 398948
rect 376726 398936 376754 398976
rect 381170 398936 381176 398948
rect 376726 398908 381176 398936
rect 381170 398896 381176 398908
rect 381228 398896 381234 398948
rect 382182 398896 382188 398948
rect 382240 398936 382246 398948
rect 382458 398936 382464 398948
rect 382240 398908 382464 398936
rect 382240 398896 382246 398908
rect 382458 398896 382464 398908
rect 382516 398896 382522 398948
rect 340414 398828 340420 398880
rect 340472 398868 340478 398880
rect 349982 398868 349988 398880
rect 340472 398840 349988 398868
rect 340472 398828 340478 398840
rect 349982 398828 349988 398840
rect 350040 398828 350046 398880
rect 354398 398828 354404 398880
rect 354456 398868 354462 398880
rect 355870 398868 355876 398880
rect 354456 398840 355876 398868
rect 354456 398828 354462 398840
rect 355870 398828 355876 398840
rect 355928 398828 355934 398880
rect 374270 398868 374276 398880
rect 363616 398840 374276 398868
rect 339126 398760 339132 398812
rect 339184 398800 339190 398812
rect 348142 398800 348148 398812
rect 339184 398772 348148 398800
rect 339184 398760 339190 398772
rect 348142 398760 348148 398772
rect 348200 398760 348206 398812
rect 348694 398760 348700 398812
rect 348752 398800 348758 398812
rect 352098 398800 352104 398812
rect 348752 398772 352104 398800
rect 348752 398760 348758 398772
rect 352098 398760 352104 398772
rect 352156 398760 352162 398812
rect 354030 398760 354036 398812
rect 354088 398800 354094 398812
rect 355410 398800 355416 398812
rect 354088 398772 355416 398800
rect 354088 398760 354094 398772
rect 355410 398760 355416 398772
rect 355468 398760 355474 398812
rect 356514 398760 356520 398812
rect 356572 398800 356578 398812
rect 363616 398800 363644 398840
rect 374270 398828 374276 398840
rect 374328 398828 374334 398880
rect 375466 398828 375472 398880
rect 375524 398828 375530 398880
rect 383010 398828 383016 398880
rect 383068 398868 383074 398880
rect 383562 398868 383568 398880
rect 383068 398840 383568 398868
rect 383068 398828 383074 398840
rect 383562 398828 383568 398840
rect 383620 398828 383626 398880
rect 385678 398828 385684 398880
rect 385736 398868 385742 398880
rect 394694 398868 394700 398880
rect 385736 398840 394700 398868
rect 385736 398828 385742 398840
rect 394694 398828 394700 398840
rect 394752 398828 394758 398880
rect 356572 398772 363644 398800
rect 356572 398760 356578 398772
rect 363690 398760 363696 398812
rect 363748 398800 363754 398812
rect 364058 398800 364064 398812
rect 363748 398772 364064 398800
rect 363748 398760 363754 398772
rect 364058 398760 364064 398772
rect 364116 398760 364122 398812
rect 365622 398760 365628 398812
rect 365680 398800 365686 398812
rect 365680 398772 374684 398800
rect 365680 398760 365686 398772
rect 343818 398692 343824 398744
rect 343876 398732 343882 398744
rect 344830 398732 344836 398744
rect 343876 398704 344836 398732
rect 343876 398692 343882 398704
rect 344830 398692 344836 398704
rect 344888 398692 344894 398744
rect 345124 398704 345428 398732
rect 330754 398624 330760 398676
rect 330812 398664 330818 398676
rect 345124 398664 345152 398704
rect 330812 398636 345152 398664
rect 345400 398664 345428 398704
rect 346026 398692 346032 398744
rect 346084 398732 346090 398744
rect 347774 398732 347780 398744
rect 346084 398704 347780 398732
rect 346084 398692 346090 398704
rect 347774 398692 347780 398704
rect 347832 398692 347838 398744
rect 348510 398692 348516 398744
rect 348568 398732 348574 398744
rect 356422 398732 356428 398744
rect 348568 398704 356428 398732
rect 348568 398692 348574 398704
rect 356422 398692 356428 398704
rect 356480 398692 356486 398744
rect 359182 398692 359188 398744
rect 359240 398732 359246 398744
rect 359550 398732 359556 398744
rect 359240 398704 359556 398732
rect 359240 398692 359246 398704
rect 359550 398692 359556 398704
rect 359608 398692 359614 398744
rect 374656 398732 374684 398772
rect 376938 398760 376944 398812
rect 376996 398800 377002 398812
rect 379054 398800 379060 398812
rect 376996 398772 379060 398800
rect 376996 398760 377002 398772
rect 379054 398760 379060 398772
rect 379112 398760 379118 398812
rect 381078 398732 381084 398744
rect 374656 398704 381084 398732
rect 381078 398692 381084 398704
rect 381136 398692 381142 398744
rect 365530 398664 365536 398676
rect 345400 398636 365536 398664
rect 330812 398624 330818 398636
rect 365530 398624 365536 398636
rect 365588 398624 365594 398676
rect 382550 398624 382556 398676
rect 382608 398664 382614 398676
rect 388070 398664 388076 398676
rect 382608 398636 388076 398664
rect 382608 398624 382614 398636
rect 388070 398624 388076 398636
rect 388128 398624 388134 398676
rect 305086 398556 305092 398608
rect 305144 398596 305150 398608
rect 340322 398596 340328 398608
rect 305144 398568 340328 398596
rect 305144 398556 305150 398568
rect 340322 398556 340328 398568
rect 340380 398556 340386 398608
rect 349246 398596 349252 398608
rect 344940 398568 349252 398596
rect 303614 398488 303620 398540
rect 303672 398528 303678 398540
rect 342898 398528 342904 398540
rect 303672 398500 342904 398528
rect 303672 398488 303678 398500
rect 342898 398488 342904 398500
rect 342956 398488 342962 398540
rect 295334 398420 295340 398472
rect 295392 398460 295398 398472
rect 343910 398460 343916 398472
rect 295392 398432 343916 398460
rect 295392 398420 295398 398432
rect 343910 398420 343916 398432
rect 343968 398420 343974 398472
rect 344940 398404 344968 398568
rect 349246 398556 349252 398568
rect 349304 398556 349310 398608
rect 351546 398556 351552 398608
rect 351604 398596 351610 398608
rect 371418 398596 371424 398608
rect 351604 398568 371424 398596
rect 351604 398556 351610 398568
rect 371418 398556 371424 398568
rect 371476 398556 371482 398608
rect 382366 398556 382372 398608
rect 382424 398596 382430 398608
rect 389266 398596 389272 398608
rect 382424 398568 389272 398596
rect 382424 398556 382430 398568
rect 389266 398556 389272 398568
rect 389324 398556 389330 398608
rect 345014 398488 345020 398540
rect 345072 398528 345078 398540
rect 345934 398528 345940 398540
rect 345072 398500 345940 398528
rect 345072 398488 345078 398500
rect 345934 398488 345940 398500
rect 345992 398488 345998 398540
rect 346118 398488 346124 398540
rect 346176 398528 346182 398540
rect 346176 398500 354674 398528
rect 346176 398488 346182 398500
rect 345658 398420 345664 398472
rect 345716 398460 345722 398472
rect 354398 398460 354404 398472
rect 345716 398432 354404 398460
rect 345716 398420 345722 398432
rect 354398 398420 354404 398432
rect 354456 398420 354462 398472
rect 354646 398460 354674 398500
rect 355502 398488 355508 398540
rect 355560 398528 355566 398540
rect 357342 398528 357348 398540
rect 355560 398500 357348 398528
rect 355560 398488 355566 398500
rect 357342 398488 357348 398500
rect 357400 398488 357406 398540
rect 359550 398488 359556 398540
rect 359608 398528 359614 398540
rect 363138 398528 363144 398540
rect 359608 398500 363144 398528
rect 359608 398488 359614 398500
rect 363138 398488 363144 398500
rect 363196 398488 363202 398540
rect 380986 398488 380992 398540
rect 381044 398528 381050 398540
rect 390646 398528 390652 398540
rect 381044 398500 390652 398528
rect 381044 398488 381050 398500
rect 390646 398488 390652 398500
rect 390704 398488 390710 398540
rect 360654 398460 360660 398472
rect 354646 398432 360660 398460
rect 360654 398420 360660 398432
rect 360712 398420 360718 398472
rect 382918 398420 382924 398472
rect 382976 398460 382982 398472
rect 389542 398460 389548 398472
rect 382976 398432 389548 398460
rect 382976 398420 382982 398432
rect 389542 398420 389548 398432
rect 389600 398420 389606 398472
rect 289078 398352 289084 398404
rect 289136 398392 289142 398404
rect 344094 398392 344100 398404
rect 289136 398364 344100 398392
rect 289136 398352 289142 398364
rect 344094 398352 344100 398364
rect 344152 398352 344158 398404
rect 344922 398352 344928 398404
rect 344980 398352 344986 398404
rect 348326 398352 348332 398404
rect 348384 398392 348390 398404
rect 362678 398392 362684 398404
rect 348384 398364 362684 398392
rect 348384 398352 348390 398364
rect 362678 398352 362684 398364
rect 362736 398352 362742 398404
rect 373810 398352 373816 398404
rect 373868 398392 373874 398404
rect 384482 398392 384488 398404
rect 373868 398364 384488 398392
rect 373868 398352 373874 398364
rect 384482 398352 384488 398364
rect 384540 398352 384546 398404
rect 386598 398352 386604 398404
rect 386656 398392 386662 398404
rect 392026 398392 392032 398404
rect 386656 398364 392032 398392
rect 386656 398352 386662 398364
rect 392026 398352 392032 398364
rect 392084 398352 392090 398404
rect 341886 398324 341892 398336
rect 331186 398296 341892 398324
rect 260742 398216 260748 398268
rect 260800 398256 260806 398268
rect 331186 398256 331214 398296
rect 341886 398284 341892 398296
rect 341944 398284 341950 398336
rect 345106 398324 345112 398336
rect 342824 398296 345112 398324
rect 260800 398228 331214 398256
rect 260800 398216 260806 398228
rect 304258 398148 304264 398200
rect 304316 398188 304322 398200
rect 305638 398188 305644 398200
rect 304316 398160 305644 398188
rect 304316 398148 304322 398160
rect 305638 398148 305644 398160
rect 305696 398148 305702 398200
rect 342824 398188 342852 398296
rect 345106 398284 345112 398296
rect 345164 398284 345170 398336
rect 346118 398324 346124 398336
rect 345400 398296 346124 398324
rect 342898 398216 342904 398268
rect 342956 398256 342962 398268
rect 345400 398256 345428 398296
rect 346118 398284 346124 398296
rect 346176 398284 346182 398336
rect 348142 398284 348148 398336
rect 348200 398324 348206 398336
rect 352098 398324 352104 398336
rect 348200 398296 352104 398324
rect 348200 398284 348206 398296
rect 352098 398284 352104 398296
rect 352156 398284 352162 398336
rect 354582 398284 354588 398336
rect 354640 398324 354646 398336
rect 360378 398324 360384 398336
rect 354640 398296 360384 398324
rect 354640 398284 354646 398296
rect 360378 398284 360384 398296
rect 360436 398284 360442 398336
rect 371418 398284 371424 398336
rect 371476 398324 371482 398336
rect 372430 398324 372436 398336
rect 371476 398296 372436 398324
rect 371476 398284 371482 398296
rect 372430 398284 372436 398296
rect 372488 398284 372494 398336
rect 342956 398228 345428 398256
rect 342956 398216 342962 398228
rect 363506 398216 363512 398268
rect 363564 398256 363570 398268
rect 365990 398256 365996 398268
rect 363564 398228 365996 398256
rect 363564 398216 363570 398228
rect 365990 398216 365996 398228
rect 366048 398216 366054 398268
rect 378778 398216 378784 398268
rect 378836 398256 378842 398268
rect 390554 398256 390560 398268
rect 378836 398228 390560 398256
rect 378836 398216 378842 398228
rect 390554 398216 390560 398228
rect 390612 398216 390618 398268
rect 354490 398188 354496 398200
rect 331186 398160 342852 398188
rect 342916 398160 354496 398188
rect 257982 398080 257988 398132
rect 258040 398120 258046 398132
rect 331186 398120 331214 398160
rect 258040 398092 331214 398120
rect 258040 398080 258046 398092
rect 341150 398080 341156 398132
rect 341208 398120 341214 398132
rect 342916 398120 342944 398160
rect 354490 398148 354496 398160
rect 354548 398148 354554 398200
rect 372430 398148 372436 398200
rect 372488 398188 372494 398200
rect 376846 398188 376852 398200
rect 372488 398160 376852 398188
rect 372488 398148 372494 398160
rect 376846 398148 376852 398160
rect 376904 398148 376910 398200
rect 386966 398148 386972 398200
rect 387024 398148 387030 398200
rect 341208 398092 342944 398120
rect 341208 398080 341214 398092
rect 353478 398080 353484 398132
rect 353536 398120 353542 398132
rect 358538 398120 358544 398132
rect 353536 398092 358544 398120
rect 353536 398080 353542 398092
rect 358538 398080 358544 398092
rect 358596 398080 358602 398132
rect 386984 398120 387012 398148
rect 386524 398092 387012 398120
rect 386524 398064 386552 398092
rect 341886 398012 341892 398064
rect 341944 398052 341950 398064
rect 357802 398052 357808 398064
rect 341944 398024 357808 398052
rect 341944 398012 341950 398024
rect 357802 398012 357808 398024
rect 357860 398012 357866 398064
rect 376846 398012 376852 398064
rect 376904 398052 376910 398064
rect 377306 398052 377312 398064
rect 376904 398024 377312 398052
rect 376904 398012 376910 398024
rect 377306 398012 377312 398024
rect 377364 398012 377370 398064
rect 377582 398012 377588 398064
rect 377640 398052 377646 398064
rect 378778 398052 378784 398064
rect 377640 398024 378784 398052
rect 377640 398012 377646 398024
rect 378778 398012 378784 398024
rect 378836 398012 378842 398064
rect 386506 398012 386512 398064
rect 386564 398012 386570 398064
rect 386966 398012 386972 398064
rect 387024 398052 387030 398064
rect 387702 398052 387708 398064
rect 387024 398024 387708 398052
rect 387024 398012 387030 398024
rect 387702 398012 387708 398024
rect 387760 398012 387766 398064
rect 342438 397944 342444 397996
rect 342496 397984 342502 397996
rect 343358 397984 343364 397996
rect 342496 397956 343364 397984
rect 342496 397944 342502 397956
rect 343358 397944 343364 397956
rect 343416 397944 343422 397996
rect 346026 397984 346032 397996
rect 343468 397956 346032 397984
rect 343468 397916 343496 397956
rect 346026 397944 346032 397956
rect 346084 397944 346090 397996
rect 352466 397944 352472 397996
rect 352524 397984 352530 397996
rect 352834 397984 352840 397996
rect 352524 397956 352840 397984
rect 352524 397944 352530 397956
rect 352834 397944 352840 397956
rect 352892 397944 352898 397996
rect 367830 397984 367836 397996
rect 355060 397956 367836 397984
rect 340846 397888 343496 397916
rect 333238 397740 333244 397792
rect 333296 397780 333302 397792
rect 340846 397780 340874 397888
rect 344830 397876 344836 397928
rect 344888 397916 344894 397928
rect 351086 397916 351092 397928
rect 344888 397888 351092 397916
rect 344888 397876 344894 397888
rect 351086 397876 351092 397888
rect 351144 397876 351150 397928
rect 352098 397876 352104 397928
rect 352156 397916 352162 397928
rect 354582 397916 354588 397928
rect 352156 397888 354588 397916
rect 352156 397876 352162 397888
rect 354582 397876 354588 397888
rect 354640 397876 354646 397928
rect 341518 397808 341524 397860
rect 341576 397848 341582 397860
rect 343082 397848 343088 397860
rect 341576 397820 343088 397848
rect 341576 397808 341582 397820
rect 343082 397808 343088 397820
rect 343140 397808 343146 397860
rect 349614 397808 349620 397860
rect 349672 397848 349678 397860
rect 350074 397848 350080 397860
rect 349672 397820 350080 397848
rect 349672 397808 349678 397820
rect 350074 397808 350080 397820
rect 350132 397808 350138 397860
rect 333296 397752 340874 397780
rect 333296 397740 333302 397752
rect 348418 397740 348424 397792
rect 348476 397780 348482 397792
rect 352374 397780 352380 397792
rect 348476 397752 352380 397780
rect 348476 397740 348482 397752
rect 352374 397740 352380 397752
rect 352432 397740 352438 397792
rect 274450 397672 274456 397724
rect 274508 397712 274514 397724
rect 345658 397712 345664 397724
rect 274508 397684 333376 397712
rect 274508 397672 274514 397684
rect 277026 397604 277032 397656
rect 277084 397644 277090 397656
rect 333238 397644 333244 397656
rect 277084 397616 333244 397644
rect 277084 397604 277090 397616
rect 333238 397604 333244 397616
rect 333296 397604 333302 397656
rect 333348 397644 333376 397684
rect 338086 397684 345664 397712
rect 338086 397644 338114 397684
rect 345658 397672 345664 397684
rect 345716 397672 345722 397724
rect 345842 397672 345848 397724
rect 345900 397712 345906 397724
rect 349430 397712 349436 397724
rect 345900 397684 349436 397712
rect 345900 397672 345906 397684
rect 349430 397672 349436 397684
rect 349488 397672 349494 397724
rect 350074 397672 350080 397724
rect 350132 397712 350138 397724
rect 355060 397712 355088 397956
rect 367830 397944 367836 397956
rect 367888 397944 367894 397996
rect 374178 397944 374184 397996
rect 374236 397984 374242 397996
rect 382918 397984 382924 397996
rect 374236 397956 382924 397984
rect 374236 397944 374242 397956
rect 382918 397944 382924 397956
rect 382976 397944 382982 397996
rect 381538 397876 381544 397928
rect 381596 397916 381602 397928
rect 381906 397916 381912 397928
rect 381596 397888 381912 397916
rect 381596 397876 381602 397888
rect 381906 397876 381912 397888
rect 381964 397876 381970 397928
rect 372246 397740 372252 397792
rect 372304 397780 372310 397792
rect 374362 397780 374368 397792
rect 372304 397752 374368 397780
rect 372304 397740 372310 397752
rect 374362 397740 374368 397752
rect 374420 397740 374426 397792
rect 381262 397740 381268 397792
rect 381320 397780 381326 397792
rect 381538 397780 381544 397792
rect 381320 397752 381544 397780
rect 381320 397740 381326 397752
rect 381538 397740 381544 397752
rect 381596 397740 381602 397792
rect 350132 397684 355088 397712
rect 350132 397672 350138 397684
rect 356422 397672 356428 397724
rect 356480 397712 356486 397724
rect 356882 397712 356888 397724
rect 356480 397684 356888 397712
rect 356480 397672 356486 397684
rect 356882 397672 356888 397684
rect 356940 397672 356946 397724
rect 361114 397672 361120 397724
rect 361172 397712 361178 397724
rect 361482 397712 361488 397724
rect 361172 397684 361488 397712
rect 361172 397672 361178 397684
rect 361482 397672 361488 397684
rect 361540 397672 361546 397724
rect 376754 397712 376760 397724
rect 371988 397684 376760 397712
rect 333348 397616 338114 397644
rect 338942 397604 338948 397656
rect 339000 397644 339006 397656
rect 355042 397644 355048 397656
rect 339000 397616 355048 397644
rect 339000 397604 339006 397616
rect 355042 397604 355048 397616
rect 355100 397604 355106 397656
rect 330846 397536 330852 397588
rect 330904 397576 330910 397588
rect 353478 397576 353484 397588
rect 330904 397548 353484 397576
rect 330904 397536 330910 397548
rect 353478 397536 353484 397548
rect 353536 397536 353542 397588
rect 355594 397536 355600 397588
rect 355652 397576 355658 397588
rect 357802 397576 357808 397588
rect 355652 397548 357808 397576
rect 355652 397536 355658 397548
rect 357802 397536 357808 397548
rect 357860 397536 357866 397588
rect 360930 397536 360936 397588
rect 360988 397576 360994 397588
rect 363598 397576 363604 397588
rect 360988 397548 363604 397576
rect 360988 397536 360994 397548
rect 363598 397536 363604 397548
rect 363656 397536 363662 397588
rect 340966 397468 340972 397520
rect 341024 397508 341030 397520
rect 346946 397508 346952 397520
rect 341024 397480 346952 397508
rect 341024 397468 341030 397480
rect 346946 397468 346952 397480
rect 347004 397468 347010 397520
rect 349430 397468 349436 397520
rect 349488 397508 349494 397520
rect 349706 397508 349712 397520
rect 349488 397480 349712 397508
rect 349488 397468 349494 397480
rect 349706 397468 349712 397480
rect 349764 397468 349770 397520
rect 351086 397468 351092 397520
rect 351144 397508 351150 397520
rect 351362 397508 351368 397520
rect 351144 397480 351368 397508
rect 351144 397468 351150 397480
rect 351362 397468 351368 397480
rect 351420 397468 351426 397520
rect 356790 397468 356796 397520
rect 356848 397508 356854 397520
rect 357986 397508 357992 397520
rect 356848 397480 357992 397508
rect 356848 397468 356854 397480
rect 357986 397468 357992 397480
rect 358044 397468 358050 397520
rect 358354 397468 358360 397520
rect 358412 397508 358418 397520
rect 362310 397508 362316 397520
rect 358412 397480 362316 397508
rect 358412 397468 358418 397480
rect 362310 397468 362316 397480
rect 362368 397468 362374 397520
rect 371988 397508 372016 397684
rect 376754 397672 376760 397684
rect 376812 397672 376818 397724
rect 386414 397672 386420 397724
rect 386472 397712 386478 397724
rect 387334 397712 387340 397724
rect 386472 397684 387340 397712
rect 386472 397672 386478 397684
rect 387334 397672 387340 397684
rect 387392 397672 387398 397724
rect 371988 397480 372108 397508
rect 372080 397452 372108 397480
rect 385310 397468 385316 397520
rect 385368 397508 385374 397520
rect 389450 397508 389456 397520
rect 385368 397480 389456 397508
rect 385368 397468 385374 397480
rect 389450 397468 389456 397480
rect 389508 397468 389514 397520
rect 334710 397400 334716 397452
rect 334768 397440 334774 397452
rect 359090 397440 359096 397452
rect 334768 397412 359096 397440
rect 334768 397400 334774 397412
rect 359090 397400 359096 397412
rect 359148 397400 359154 397452
rect 372062 397400 372068 397452
rect 372120 397400 372126 397452
rect 386414 397400 386420 397452
rect 386472 397440 386478 397452
rect 387518 397440 387524 397452
rect 386472 397412 387524 397440
rect 386472 397400 386478 397412
rect 387518 397400 387524 397412
rect 387576 397400 387582 397452
rect 345658 397332 345664 397384
rect 345716 397372 345722 397384
rect 362494 397372 362500 397384
rect 345716 397344 362500 397372
rect 345716 397332 345722 397344
rect 362494 397332 362500 397344
rect 362552 397332 362558 397384
rect 364518 397332 364524 397384
rect 364576 397372 364582 397384
rect 364702 397372 364708 397384
rect 364576 397344 364708 397372
rect 364576 397332 364582 397344
rect 364702 397332 364708 397344
rect 364760 397332 364766 397384
rect 365990 397332 365996 397384
rect 366048 397372 366054 397384
rect 366174 397372 366180 397384
rect 366048 397344 366180 397372
rect 366048 397332 366054 397344
rect 366174 397332 366180 397344
rect 366232 397332 366238 397384
rect 382366 397332 382372 397384
rect 382424 397372 382430 397384
rect 382734 397372 382740 397384
rect 382424 397344 382740 397372
rect 382424 397332 382430 397344
rect 382734 397332 382740 397344
rect 382792 397332 382798 397384
rect 385678 397332 385684 397384
rect 385736 397372 385742 397384
rect 385954 397372 385960 397384
rect 385736 397344 385960 397372
rect 385736 397332 385742 397344
rect 385954 397332 385960 397344
rect 386012 397332 386018 397384
rect 332318 397264 332324 397316
rect 332376 397304 332382 397316
rect 359642 397304 359648 397316
rect 332376 397276 359648 397304
rect 332376 397264 332382 397276
rect 359642 397264 359648 397276
rect 359700 397264 359706 397316
rect 330662 397196 330668 397248
rect 330720 397236 330726 397248
rect 358630 397236 358636 397248
rect 330720 397208 358636 397236
rect 330720 397196 330726 397208
rect 358630 397196 358636 397208
rect 358688 397196 358694 397248
rect 383746 397196 383752 397248
rect 383804 397236 383810 397248
rect 389358 397236 389364 397248
rect 383804 397208 389364 397236
rect 383804 397196 383810 397208
rect 389358 397196 389364 397208
rect 389416 397196 389422 397248
rect 337838 397128 337844 397180
rect 337896 397168 337902 397180
rect 380618 397168 380624 397180
rect 337896 397140 380624 397168
rect 337896 397128 337902 397140
rect 380618 397128 380624 397140
rect 380676 397128 380682 397180
rect 380986 397128 380992 397180
rect 381044 397168 381050 397180
rect 382642 397168 382648 397180
rect 381044 397140 382648 397168
rect 381044 397128 381050 397140
rect 382642 397128 382648 397140
rect 382700 397128 382706 397180
rect 384298 397128 384304 397180
rect 384356 397168 384362 397180
rect 384574 397168 384580 397180
rect 384356 397140 384580 397168
rect 384356 397128 384362 397140
rect 384574 397128 384580 397140
rect 384632 397128 384638 397180
rect 336182 397060 336188 397112
rect 336240 397100 336246 397112
rect 383286 397100 383292 397112
rect 336240 397072 383292 397100
rect 336240 397060 336246 397072
rect 383286 397060 383292 397072
rect 383344 397060 383350 397112
rect 306282 396992 306288 397044
rect 306340 397032 306346 397044
rect 366358 397032 366364 397044
rect 306340 397004 366364 397032
rect 306340 396992 306346 397004
rect 366358 396992 366364 397004
rect 366416 396992 366422 397044
rect 386690 396992 386696 397044
rect 386748 397032 386754 397044
rect 387242 397032 387248 397044
rect 386748 397004 387248 397032
rect 386748 396992 386754 397004
rect 387242 396992 387248 397004
rect 387300 396992 387306 397044
rect 276934 396924 276940 396976
rect 276992 396964 276998 396976
rect 339862 396964 339868 396976
rect 276992 396936 339868 396964
rect 276992 396924 276998 396936
rect 339862 396924 339868 396936
rect 339920 396924 339926 396976
rect 349154 396924 349160 396976
rect 349212 396964 349218 396976
rect 349522 396964 349528 396976
rect 349212 396936 349528 396964
rect 349212 396924 349218 396936
rect 349522 396924 349528 396936
rect 349580 396924 349586 396976
rect 377858 396924 377864 396976
rect 377916 396964 377922 396976
rect 381078 396964 381084 396976
rect 377916 396936 381084 396964
rect 377916 396924 377922 396936
rect 381078 396924 381084 396936
rect 381136 396924 381142 396976
rect 280982 396856 280988 396908
rect 281040 396896 281046 396908
rect 350442 396896 350448 396908
rect 281040 396868 350448 396896
rect 281040 396856 281046 396868
rect 350442 396856 350448 396868
rect 350500 396856 350506 396908
rect 355686 396856 355692 396908
rect 355744 396896 355750 396908
rect 360838 396896 360844 396908
rect 355744 396868 360844 396896
rect 355744 396856 355750 396868
rect 360838 396856 360844 396868
rect 360896 396856 360902 396908
rect 362310 396856 362316 396908
rect 362368 396896 362374 396908
rect 371970 396896 371976 396908
rect 362368 396868 371976 396896
rect 362368 396856 362374 396868
rect 371970 396856 371976 396868
rect 372028 396856 372034 396908
rect 378502 396856 378508 396908
rect 378560 396896 378566 396908
rect 381262 396896 381268 396908
rect 378560 396868 381268 396896
rect 378560 396856 378566 396868
rect 381262 396856 381268 396868
rect 381320 396856 381326 396908
rect 390002 396856 390008 396908
rect 390060 396896 390066 396908
rect 394878 396896 394884 396908
rect 390060 396868 394884 396896
rect 390060 396856 390066 396868
rect 394878 396856 394884 396868
rect 394936 396856 394942 396908
rect 271506 396788 271512 396840
rect 271564 396828 271570 396840
rect 353110 396828 353116 396840
rect 271564 396800 353116 396828
rect 271564 396788 271570 396800
rect 353110 396788 353116 396800
rect 353168 396788 353174 396840
rect 354490 396788 354496 396840
rect 354548 396828 354554 396840
rect 354950 396828 354956 396840
rect 354548 396800 354956 396828
rect 354548 396788 354554 396800
rect 354950 396788 354956 396800
rect 355008 396788 355014 396840
rect 377858 396788 377864 396840
rect 377916 396828 377922 396840
rect 379698 396828 379704 396840
rect 377916 396800 379704 396828
rect 377916 396788 377922 396800
rect 379698 396788 379704 396800
rect 379756 396788 379762 396840
rect 340598 396720 340604 396772
rect 340656 396760 340662 396772
rect 345658 396760 345664 396772
rect 340656 396732 345664 396760
rect 340656 396720 340662 396732
rect 345658 396720 345664 396732
rect 345716 396720 345722 396772
rect 355134 396720 355140 396772
rect 355192 396760 355198 396772
rect 360746 396760 360752 396772
rect 355192 396732 360752 396760
rect 355192 396720 355198 396732
rect 360746 396720 360752 396732
rect 360804 396720 360810 396772
rect 367922 396720 367928 396772
rect 367980 396760 367986 396772
rect 368658 396760 368664 396772
rect 367980 396732 368664 396760
rect 367980 396720 367986 396732
rect 368658 396720 368664 396732
rect 368716 396720 368722 396772
rect 377306 396720 377312 396772
rect 377364 396760 377370 396772
rect 381446 396760 381452 396772
rect 377364 396732 381452 396760
rect 377364 396720 377370 396732
rect 381446 396720 381452 396732
rect 381504 396720 381510 396772
rect 346026 396652 346032 396704
rect 346084 396692 346090 396704
rect 351178 396692 351184 396704
rect 346084 396664 351184 396692
rect 346084 396652 346090 396664
rect 351178 396652 351184 396664
rect 351236 396652 351242 396704
rect 358262 396652 358268 396704
rect 358320 396692 358326 396704
rect 358814 396692 358820 396704
rect 358320 396664 358820 396692
rect 358320 396652 358326 396664
rect 358814 396652 358820 396664
rect 358872 396652 358878 396704
rect 363506 396652 363512 396704
rect 363564 396692 363570 396704
rect 363966 396692 363972 396704
rect 363564 396664 363972 396692
rect 363564 396652 363570 396664
rect 363966 396652 363972 396664
rect 364024 396652 364030 396704
rect 377398 396652 377404 396704
rect 377456 396692 377462 396704
rect 377674 396692 377680 396704
rect 377456 396664 377680 396692
rect 377456 396652 377462 396664
rect 377674 396652 377680 396664
rect 377732 396652 377738 396704
rect 383930 396652 383936 396704
rect 383988 396692 383994 396704
rect 384114 396692 384120 396704
rect 383988 396664 384120 396692
rect 383988 396652 383994 396664
rect 384114 396652 384120 396664
rect 384172 396652 384178 396704
rect 385218 396652 385224 396704
rect 385276 396692 385282 396704
rect 385862 396692 385868 396704
rect 385276 396664 385868 396692
rect 385276 396652 385282 396664
rect 385862 396652 385868 396664
rect 385920 396652 385926 396704
rect 257798 396584 257804 396636
rect 257856 396624 257862 396636
rect 343634 396624 343640 396636
rect 257856 396596 343640 396624
rect 257856 396584 257862 396596
rect 343634 396584 343640 396596
rect 343692 396584 343698 396636
rect 363414 396584 363420 396636
rect 363472 396624 363478 396636
rect 363874 396624 363880 396636
rect 363472 396596 363880 396624
rect 363472 396584 363478 396596
rect 363874 396584 363880 396596
rect 363932 396584 363938 396636
rect 335998 396516 336004 396568
rect 336056 396556 336062 396568
rect 352006 396556 352012 396568
rect 336056 396528 352012 396556
rect 336056 396516 336062 396528
rect 352006 396516 352012 396528
rect 352064 396516 352070 396568
rect 382642 396516 382648 396568
rect 382700 396556 382706 396568
rect 383378 396556 383384 396568
rect 382700 396528 383384 396556
rect 382700 396516 382706 396528
rect 383378 396516 383384 396528
rect 383436 396516 383442 396568
rect 355870 396448 355876 396500
rect 355928 396488 355934 396500
rect 361574 396488 361580 396500
rect 355928 396460 361580 396488
rect 355928 396448 355934 396460
rect 361574 396448 361580 396460
rect 361632 396448 361638 396500
rect 383930 396448 383936 396500
rect 383988 396488 383994 396500
rect 384666 396488 384672 396500
rect 383988 396460 384672 396488
rect 383988 396448 383994 396460
rect 384666 396448 384672 396460
rect 384724 396448 384730 396500
rect 360838 396312 360844 396364
rect 360896 396352 360902 396364
rect 362954 396352 362960 396364
rect 360896 396324 362960 396352
rect 360896 396312 360902 396324
rect 362954 396312 362960 396324
rect 363012 396312 363018 396364
rect 351178 396176 351184 396228
rect 351236 396216 351242 396228
rect 355318 396216 355324 396228
rect 351236 396188 355324 396216
rect 351236 396176 351242 396188
rect 355318 396176 355324 396188
rect 355376 396176 355382 396228
rect 372706 396176 372712 396228
rect 372764 396216 372770 396228
rect 373258 396216 373264 396228
rect 372764 396188 373264 396216
rect 372764 396176 372770 396188
rect 373258 396176 373264 396188
rect 373316 396176 373322 396228
rect 341794 396108 341800 396160
rect 341852 396148 341858 396160
rect 354766 396148 354772 396160
rect 341852 396120 354772 396148
rect 341852 396108 341858 396120
rect 354766 396108 354772 396120
rect 354824 396108 354830 396160
rect 385494 396108 385500 396160
rect 385552 396148 385558 396160
rect 386230 396148 386236 396160
rect 385552 396120 386236 396148
rect 385552 396108 385558 396120
rect 386230 396108 386236 396120
rect 386288 396108 386294 396160
rect 346486 396040 346492 396092
rect 346544 396080 346550 396092
rect 346854 396080 346860 396092
rect 346544 396052 346860 396080
rect 346544 396040 346550 396052
rect 346854 396040 346860 396052
rect 346912 396040 346918 396092
rect 361850 396080 361856 396092
rect 354646 396052 361856 396080
rect 335078 395972 335084 396024
rect 335136 396012 335142 396024
rect 354646 396012 354674 396052
rect 361850 396040 361856 396052
rect 361908 396040 361914 396092
rect 335136 395984 354674 396012
rect 335136 395972 335142 395984
rect 360102 395972 360108 396024
rect 360160 396012 360166 396024
rect 363690 396012 363696 396024
rect 360160 395984 363696 396012
rect 360160 395972 360166 395984
rect 363690 395972 363696 395984
rect 363748 395972 363754 396024
rect 379514 395972 379520 396024
rect 379572 396012 379578 396024
rect 379790 396012 379796 396024
rect 379572 395984 379796 396012
rect 379572 395972 379578 395984
rect 379790 395972 379796 395984
rect 379848 395972 379854 396024
rect 341702 395904 341708 395956
rect 341760 395944 341766 395956
rect 368934 395944 368940 395956
rect 341760 395916 368940 395944
rect 341760 395904 341766 395916
rect 368934 395904 368940 395916
rect 368992 395904 368998 395956
rect 381446 395904 381452 395956
rect 381504 395944 381510 395956
rect 381998 395944 382004 395956
rect 381504 395916 382004 395944
rect 381504 395904 381510 395916
rect 381998 395904 382004 395916
rect 382056 395904 382062 395956
rect 340138 395836 340144 395888
rect 340196 395876 340202 395888
rect 368014 395876 368020 395888
rect 340196 395848 368020 395876
rect 340196 395836 340202 395848
rect 368014 395836 368020 395848
rect 368072 395836 368078 395888
rect 336366 395768 336372 395820
rect 336424 395808 336430 395820
rect 369670 395808 369676 395820
rect 336424 395780 369676 395808
rect 336424 395768 336430 395780
rect 369670 395768 369676 395780
rect 369728 395768 369734 395820
rect 330570 395700 330576 395752
rect 330628 395740 330634 395752
rect 365438 395740 365444 395752
rect 330628 395712 365444 395740
rect 330628 395700 330634 395712
rect 365438 395700 365444 395712
rect 365496 395700 365502 395752
rect 281626 395632 281632 395684
rect 281684 395672 281690 395684
rect 303614 395672 303620 395684
rect 281684 395644 303620 395672
rect 281684 395632 281690 395644
rect 303614 395632 303620 395644
rect 303672 395632 303678 395684
rect 329282 395632 329288 395684
rect 329340 395672 329346 395684
rect 368198 395672 368204 395684
rect 329340 395644 368204 395672
rect 329340 395632 329346 395644
rect 368198 395632 368204 395644
rect 368256 395632 368262 395684
rect 369026 395632 369032 395684
rect 369084 395672 369090 395684
rect 369762 395672 369768 395684
rect 369084 395644 369768 395672
rect 369084 395632 369090 395644
rect 369762 395632 369768 395644
rect 369820 395632 369826 395684
rect 372522 395632 372528 395684
rect 372580 395672 372586 395684
rect 374546 395672 374552 395684
rect 372580 395644 374552 395672
rect 372580 395632 372586 395644
rect 374546 395632 374552 395644
rect 374604 395632 374610 395684
rect 383654 395632 383660 395684
rect 383712 395672 383718 395684
rect 384390 395672 384396 395684
rect 383712 395644 384396 395672
rect 383712 395632 383718 395644
rect 384390 395632 384396 395644
rect 384448 395632 384454 395684
rect 281534 395564 281540 395616
rect 281592 395604 281598 395616
rect 305086 395604 305092 395616
rect 281592 395576 305092 395604
rect 281592 395564 281598 395576
rect 305086 395564 305092 395576
rect 305144 395564 305150 395616
rect 339310 395564 339316 395616
rect 339368 395604 339374 395616
rect 381630 395604 381636 395616
rect 339368 395576 381636 395604
rect 339368 395564 339374 395576
rect 381630 395564 381636 395576
rect 381688 395564 381694 395616
rect 385402 395564 385408 395616
rect 385460 395604 385466 395616
rect 386322 395604 386328 395616
rect 385460 395576 386328 395604
rect 385460 395564 385466 395576
rect 386322 395564 386328 395576
rect 386380 395564 386386 395616
rect 278406 395496 278412 395548
rect 278464 395536 278470 395548
rect 347958 395536 347964 395548
rect 278464 395508 347964 395536
rect 278464 395496 278470 395508
rect 347958 395496 347964 395508
rect 348016 395496 348022 395548
rect 350902 395496 350908 395548
rect 350960 395536 350966 395548
rect 351730 395536 351736 395548
rect 350960 395508 351736 395536
rect 350960 395496 350966 395508
rect 351730 395496 351736 395508
rect 351788 395496 351794 395548
rect 356974 395496 356980 395548
rect 357032 395536 357038 395548
rect 361022 395536 361028 395548
rect 357032 395508 361028 395536
rect 357032 395496 357038 395508
rect 361022 395496 361028 395508
rect 361080 395496 361086 395548
rect 366358 395496 366364 395548
rect 366416 395536 366422 395548
rect 370590 395536 370596 395548
rect 366416 395508 370596 395536
rect 366416 395496 366422 395508
rect 370590 395496 370596 395508
rect 370648 395496 370654 395548
rect 275554 395428 275560 395480
rect 275612 395468 275618 395480
rect 353662 395468 353668 395480
rect 275612 395440 353668 395468
rect 275612 395428 275618 395440
rect 353662 395428 353668 395440
rect 353720 395428 353726 395480
rect 378134 395428 378140 395480
rect 378192 395468 378198 395480
rect 379974 395468 379980 395480
rect 378192 395440 379980 395468
rect 378192 395428 378198 395440
rect 379974 395428 379980 395440
rect 380032 395428 380038 395480
rect 346854 395360 346860 395412
rect 346912 395400 346918 395412
rect 347406 395400 347412 395412
rect 346912 395372 347412 395400
rect 346912 395360 346918 395372
rect 347406 395360 347412 395372
rect 347464 395360 347470 395412
rect 354858 395360 354864 395412
rect 354916 395400 354922 395412
rect 356054 395400 356060 395412
rect 354916 395372 356060 395400
rect 354916 395360 354922 395372
rect 356054 395360 356060 395372
rect 356112 395360 356118 395412
rect 361022 395360 361028 395412
rect 361080 395400 361086 395412
rect 374638 395400 374644 395412
rect 361080 395372 374644 395400
rect 361080 395360 361086 395372
rect 374638 395360 374644 395372
rect 374696 395360 374702 395412
rect 275738 395292 275744 395344
rect 275796 395332 275802 395344
rect 341794 395332 341800 395344
rect 275796 395304 341800 395332
rect 275796 395292 275802 395304
rect 341794 395292 341800 395304
rect 341852 395292 341858 395344
rect 352742 395332 352748 395344
rect 343560 395304 352748 395332
rect 337654 395224 337660 395276
rect 337712 395264 337718 395276
rect 343560 395264 343588 395304
rect 352742 395292 352748 395304
rect 352800 395292 352806 395344
rect 355962 395292 355968 395344
rect 356020 395332 356026 395344
rect 356020 395304 368704 395332
rect 356020 395292 356026 395304
rect 337712 395236 343588 395264
rect 337712 395224 337718 395236
rect 343634 395224 343640 395276
rect 343692 395264 343698 395276
rect 350810 395264 350816 395276
rect 343692 395236 350816 395264
rect 343692 395224 343698 395236
rect 350810 395224 350816 395236
rect 350868 395224 350874 395276
rect 353478 395224 353484 395276
rect 353536 395264 353542 395276
rect 354306 395264 354312 395276
rect 353536 395236 354312 395264
rect 353536 395224 353542 395236
rect 354306 395224 354312 395236
rect 354364 395224 354370 395276
rect 367738 395224 367744 395276
rect 367796 395264 367802 395276
rect 368566 395264 368572 395276
rect 367796 395236 368572 395264
rect 367796 395224 367802 395236
rect 368566 395224 368572 395236
rect 368624 395224 368630 395276
rect 368676 395264 368704 395304
rect 369762 395292 369768 395344
rect 369820 395332 369826 395344
rect 371602 395332 371608 395344
rect 369820 395304 371608 395332
rect 369820 395292 369826 395304
rect 371602 395292 371608 395304
rect 371660 395292 371666 395344
rect 371786 395292 371792 395344
rect 371844 395332 371850 395344
rect 372154 395332 372160 395344
rect 371844 395304 372160 395332
rect 371844 395292 371850 395304
rect 372154 395292 372160 395304
rect 372212 395292 372218 395344
rect 374270 395292 374276 395344
rect 374328 395332 374334 395344
rect 375282 395332 375288 395344
rect 374328 395304 375288 395332
rect 374328 395292 374334 395304
rect 375282 395292 375288 395304
rect 375340 395292 375346 395344
rect 369946 395264 369952 395276
rect 368676 395236 369952 395264
rect 369946 395224 369952 395236
rect 370004 395224 370010 395276
rect 374638 395224 374644 395276
rect 374696 395264 374702 395276
rect 375558 395264 375564 395276
rect 374696 395236 375564 395264
rect 374696 395224 374702 395236
rect 375558 395224 375564 395236
rect 375616 395224 375622 395276
rect 375834 395224 375840 395276
rect 375892 395264 375898 395276
rect 376386 395264 376392 395276
rect 375892 395236 376392 395264
rect 375892 395224 375898 395236
rect 376386 395224 376392 395236
rect 376444 395224 376450 395276
rect 327994 395156 328000 395208
rect 328052 395196 328058 395208
rect 343542 395196 343548 395208
rect 328052 395168 343548 395196
rect 328052 395156 328058 395168
rect 343542 395156 343548 395168
rect 343600 395156 343606 395208
rect 374178 395156 374184 395208
rect 374236 395196 374242 395208
rect 375098 395196 375104 395208
rect 374236 395168 375104 395196
rect 374236 395156 374242 395168
rect 375098 395156 375104 395168
rect 375156 395156 375162 395208
rect 267642 395088 267648 395140
rect 267700 395128 267706 395140
rect 345014 395128 345020 395140
rect 267700 395100 345020 395128
rect 267700 395088 267706 395100
rect 345014 395088 345020 395100
rect 345072 395088 345078 395140
rect 364886 395088 364892 395140
rect 364944 395128 364950 395140
rect 365070 395128 365076 395140
rect 364944 395100 365076 395128
rect 364944 395088 364950 395100
rect 365070 395088 365076 395100
rect 365128 395088 365134 395140
rect 370038 395088 370044 395140
rect 370096 395128 370102 395140
rect 371602 395128 371608 395140
rect 370096 395100 371608 395128
rect 370096 395088 370102 395100
rect 371602 395088 371608 395100
rect 371660 395088 371666 395140
rect 378226 395088 378232 395140
rect 378284 395128 378290 395140
rect 390738 395128 390744 395140
rect 378284 395100 390744 395128
rect 378284 395088 378290 395100
rect 390738 395088 390744 395100
rect 390796 395088 390802 395140
rect 361758 395020 361764 395072
rect 361816 395060 361822 395072
rect 362218 395060 362224 395072
rect 361816 395032 362224 395060
rect 361816 395020 361822 395032
rect 362218 395020 362224 395032
rect 362276 395020 362282 395072
rect 345014 394952 345020 395004
rect 345072 394992 345078 395004
rect 350626 394992 350632 395004
rect 345072 394964 350632 394992
rect 345072 394952 345078 394964
rect 350626 394952 350632 394964
rect 350684 394952 350690 395004
rect 353018 394952 353024 395004
rect 353076 394992 353082 395004
rect 354214 394992 354220 395004
rect 353076 394964 354220 394992
rect 353076 394952 353082 394964
rect 354214 394952 354220 394964
rect 354272 394952 354278 395004
rect 361850 394680 361856 394732
rect 361908 394720 361914 394732
rect 362586 394720 362592 394732
rect 361908 394692 362592 394720
rect 361908 394680 361914 394692
rect 362586 394680 362592 394692
rect 362644 394680 362650 394732
rect 341610 394612 341616 394664
rect 341668 394652 341674 394664
rect 360010 394652 360016 394664
rect 341668 394624 360016 394652
rect 341668 394612 341674 394624
rect 360010 394612 360016 394624
rect 360068 394612 360074 394664
rect 334894 394544 334900 394596
rect 334952 394584 334958 394596
rect 359182 394584 359188 394596
rect 334952 394556 359188 394584
rect 334952 394544 334958 394556
rect 359182 394544 359188 394556
rect 359240 394544 359246 394596
rect 336550 394476 336556 394528
rect 336608 394516 336614 394528
rect 368934 394516 368940 394528
rect 336608 394488 368940 394516
rect 336608 394476 336614 394488
rect 368934 394476 368940 394488
rect 368992 394476 368998 394528
rect 339218 394408 339224 394460
rect 339276 394448 339282 394460
rect 378962 394448 378968 394460
rect 339276 394420 378968 394448
rect 339276 394408 339282 394420
rect 378962 394408 378968 394420
rect 379020 394408 379026 394460
rect 322842 394340 322848 394392
rect 322900 394380 322906 394392
rect 382274 394380 382280 394392
rect 322900 394352 382280 394380
rect 322900 394340 322906 394352
rect 382274 394340 382280 394352
rect 382332 394340 382338 394392
rect 272978 394272 272984 394324
rect 273036 394312 273042 394324
rect 345750 394312 345756 394324
rect 273036 394284 345756 394312
rect 273036 394272 273042 394284
rect 345750 394272 345756 394284
rect 345808 394272 345814 394324
rect 358906 394312 358912 394324
rect 352024 394284 358912 394312
rect 276750 394204 276756 394256
rect 276808 394244 276814 394256
rect 339862 394244 339868 394256
rect 276808 394216 339868 394244
rect 276808 394204 276814 394216
rect 339862 394204 339868 394216
rect 339920 394204 339926 394256
rect 279694 394136 279700 394188
rect 279752 394176 279758 394188
rect 352024 394176 352052 394284
rect 358906 394272 358912 394284
rect 358964 394272 358970 394324
rect 358998 394272 359004 394324
rect 359056 394312 359062 394324
rect 359734 394312 359740 394324
rect 359056 394284 359740 394312
rect 359056 394272 359062 394284
rect 359734 394272 359740 394284
rect 359792 394272 359798 394324
rect 352742 394204 352748 394256
rect 352800 394244 352806 394256
rect 374822 394244 374828 394256
rect 352800 394216 374828 394244
rect 352800 394204 352806 394216
rect 374822 394204 374828 394216
rect 374880 394204 374886 394256
rect 375558 394204 375564 394256
rect 375616 394244 375622 394256
rect 376478 394244 376484 394256
rect 375616 394216 376484 394244
rect 375616 394204 375622 394216
rect 376478 394204 376484 394216
rect 376536 394204 376542 394256
rect 380066 394204 380072 394256
rect 380124 394244 380130 394256
rect 380342 394244 380348 394256
rect 380124 394216 380348 394244
rect 380124 394204 380130 394216
rect 380342 394204 380348 394216
rect 380400 394204 380406 394256
rect 279752 394148 352052 394176
rect 279752 394136 279758 394148
rect 354122 394136 354128 394188
rect 354180 394176 354186 394188
rect 354180 394148 360194 394176
rect 354180 394136 354186 394148
rect 264790 394068 264796 394120
rect 264848 394108 264854 394120
rect 342438 394108 342444 394120
rect 264848 394080 342444 394108
rect 264848 394068 264854 394080
rect 342438 394068 342444 394080
rect 342496 394068 342502 394120
rect 360166 394108 360194 394148
rect 385126 394136 385132 394188
rect 385184 394176 385190 394188
rect 385770 394176 385776 394188
rect 385184 394148 385776 394176
rect 385184 394136 385190 394148
rect 385770 394136 385776 394148
rect 385828 394136 385834 394188
rect 376846 394108 376852 394120
rect 342916 394080 352788 394108
rect 360166 394080 376852 394108
rect 272610 394000 272616 394052
rect 272668 394040 272674 394052
rect 342916 394040 342944 394080
rect 272668 394012 342944 394040
rect 272668 394000 272674 394012
rect 342990 394000 342996 394052
rect 343048 394040 343054 394052
rect 347038 394040 347044 394052
rect 343048 394012 347044 394040
rect 343048 394000 343054 394012
rect 347038 394000 347044 394012
rect 347096 394000 347102 394052
rect 352374 394000 352380 394052
rect 352432 394040 352438 394052
rect 352650 394040 352656 394052
rect 352432 394012 352656 394040
rect 352432 394000 352438 394012
rect 352650 394000 352656 394012
rect 352708 394000 352714 394052
rect 352760 394040 352788 394080
rect 376846 394068 376852 394080
rect 376904 394068 376910 394120
rect 386046 394068 386052 394120
rect 386104 394108 386110 394120
rect 389634 394108 389640 394120
rect 386104 394080 389640 394108
rect 386104 394068 386110 394080
rect 389634 394068 389640 394080
rect 389692 394068 389698 394120
rect 355226 394040 355232 394052
rect 352760 394012 355232 394040
rect 355226 394000 355232 394012
rect 355284 394000 355290 394052
rect 356238 394000 356244 394052
rect 356296 394040 356302 394052
rect 357250 394040 357256 394052
rect 356296 394012 357256 394040
rect 356296 394000 356302 394012
rect 357250 394000 357256 394012
rect 357308 394000 357314 394052
rect 273990 393932 273996 393984
rect 274048 393972 274054 393984
rect 274048 393944 350534 393972
rect 274048 393932 274054 393944
rect 342530 393864 342536 393916
rect 342588 393904 342594 393916
rect 343266 393904 343272 393916
rect 342588 393876 343272 393904
rect 342588 393864 342594 393876
rect 343266 393864 343272 393876
rect 343324 393864 343330 393916
rect 342438 393796 342444 393848
rect 342496 393836 342502 393848
rect 344370 393836 344376 393848
rect 342496 393808 344376 393836
rect 342496 393796 342502 393808
rect 344370 393796 344376 393808
rect 344428 393796 344434 393848
rect 350506 393768 350534 393944
rect 357158 393932 357164 393984
rect 357216 393972 357222 393984
rect 359458 393972 359464 393984
rect 357216 393944 359464 393972
rect 357216 393932 357222 393944
rect 359458 393932 359464 393944
rect 359516 393932 359522 393984
rect 376018 393932 376024 393984
rect 376076 393972 376082 393984
rect 376294 393972 376300 393984
rect 376076 393944 376300 393972
rect 376076 393932 376082 393944
rect 376294 393932 376300 393944
rect 376352 393932 376358 393984
rect 350626 393796 350632 393848
rect 350684 393836 350690 393848
rect 351362 393836 351368 393848
rect 350684 393808 351368 393836
rect 350684 393796 350690 393808
rect 351362 393796 351368 393808
rect 351420 393796 351426 393848
rect 352098 393796 352104 393848
rect 352156 393836 352162 393848
rect 352558 393836 352564 393848
rect 352156 393808 352564 393836
rect 352156 393796 352162 393808
rect 352558 393796 352564 393808
rect 352616 393796 352622 393848
rect 376018 393796 376024 393848
rect 376076 393836 376082 393848
rect 376570 393836 376576 393848
rect 376076 393808 376576 393836
rect 376076 393796 376082 393808
rect 376570 393796 376576 393808
rect 376628 393796 376634 393848
rect 377214 393796 377220 393848
rect 377272 393836 377278 393848
rect 377766 393836 377772 393848
rect 377272 393808 377772 393836
rect 377272 393796 377278 393808
rect 377766 393796 377772 393808
rect 377824 393796 377830 393848
rect 364886 393768 364892 393780
rect 350506 393740 364892 393768
rect 364886 393728 364892 393740
rect 364944 393728 364950 393780
rect 374822 393728 374828 393780
rect 374880 393768 374886 393780
rect 377490 393768 377496 393780
rect 374880 393740 377496 393768
rect 374880 393728 374886 393740
rect 377490 393728 377496 393740
rect 377548 393728 377554 393780
rect 378870 393592 378876 393644
rect 378928 393632 378934 393644
rect 379238 393632 379244 393644
rect 378928 393604 379244 393632
rect 378928 393592 378934 393604
rect 379238 393592 379244 393604
rect 379296 393592 379302 393644
rect 345658 393524 345664 393576
rect 345716 393564 345722 393576
rect 347498 393564 347504 393576
rect 345716 393536 347504 393564
rect 345716 393524 345722 393536
rect 347498 393524 347504 393536
rect 347556 393524 347562 393576
rect 348694 393524 348700 393576
rect 348752 393564 348758 393576
rect 349246 393564 349252 393576
rect 348752 393536 349252 393564
rect 348752 393524 348758 393536
rect 349246 393524 349252 393536
rect 349304 393524 349310 393576
rect 363414 393524 363420 393576
rect 363472 393564 363478 393576
rect 364242 393564 364248 393576
rect 363472 393536 364248 393564
rect 363472 393524 363478 393536
rect 364242 393524 364248 393536
rect 364300 393524 364306 393576
rect 345290 393456 345296 393508
rect 345348 393496 345354 393508
rect 346670 393496 346676 393508
rect 345348 393468 346676 393496
rect 345348 393456 345354 393468
rect 346670 393456 346676 393468
rect 346728 393456 346734 393508
rect 351362 393456 351368 393508
rect 351420 393496 351426 393508
rect 353846 393496 353852 393508
rect 351420 393468 353852 393496
rect 351420 393456 351426 393468
rect 353846 393456 353852 393468
rect 353904 393456 353910 393508
rect 363138 393456 363144 393508
rect 363196 393496 363202 393508
rect 364150 393496 364156 393508
rect 363196 393468 364156 393496
rect 363196 393456 363202 393468
rect 364150 393456 364156 393468
rect 364208 393456 364214 393508
rect 364518 393456 364524 393508
rect 364576 393496 364582 393508
rect 364886 393496 364892 393508
rect 364576 393468 364892 393496
rect 364576 393456 364582 393468
rect 364886 393456 364892 393468
rect 364944 393456 364950 393508
rect 367462 393456 367468 393508
rect 367520 393496 367526 393508
rect 368842 393496 368848 393508
rect 367520 393468 368848 393496
rect 367520 393456 367526 393468
rect 368842 393456 368848 393468
rect 368900 393456 368906 393508
rect 339034 393388 339040 393440
rect 339092 393428 339098 393440
rect 346578 393428 346584 393440
rect 339092 393400 346584 393428
rect 339092 393388 339098 393400
rect 346578 393388 346584 393400
rect 346636 393388 346642 393440
rect 347958 393388 347964 393440
rect 348016 393428 348022 393440
rect 349062 393428 349068 393440
rect 348016 393400 349068 393428
rect 348016 393388 348022 393400
rect 349062 393388 349068 393400
rect 349120 393388 349126 393440
rect 349522 393388 349528 393440
rect 349580 393428 349586 393440
rect 349798 393428 349804 393440
rect 349580 393400 349804 393428
rect 349580 393388 349586 393400
rect 349798 393388 349804 393400
rect 349856 393388 349862 393440
rect 360470 393388 360476 393440
rect 360528 393428 360534 393440
rect 361482 393428 361488 393440
rect 360528 393400 361488 393428
rect 360528 393388 360534 393400
rect 361482 393388 361488 393400
rect 361540 393388 361546 393440
rect 362218 393388 362224 393440
rect 362276 393428 362282 393440
rect 370222 393428 370228 393440
rect 362276 393400 370228 393428
rect 362276 393388 362282 393400
rect 370222 393388 370228 393400
rect 370280 393388 370286 393440
rect 321370 393320 321376 393372
rect 321428 393360 321434 393372
rect 378134 393360 378140 393372
rect 321428 393332 378140 393360
rect 321428 393320 321434 393332
rect 378134 393320 378140 393332
rect 378192 393320 378198 393372
rect 282914 393252 282920 393304
rect 282972 393292 282978 393304
rect 344370 393292 344376 393304
rect 282972 393264 344376 393292
rect 282972 393252 282978 393264
rect 344370 393252 344376 393264
rect 344428 393252 344434 393304
rect 346762 393252 346768 393304
rect 346820 393292 346826 393304
rect 347314 393292 347320 393304
rect 346820 393264 347320 393292
rect 346820 393252 346826 393264
rect 347314 393252 347320 393264
rect 347372 393252 347378 393304
rect 348786 393252 348792 393304
rect 348844 393292 348850 393304
rect 349062 393292 349068 393304
rect 348844 393264 349068 393292
rect 348844 393252 348850 393264
rect 349062 393252 349068 393264
rect 349120 393252 349126 393304
rect 349246 393252 349252 393304
rect 349304 393292 349310 393304
rect 350534 393292 350540 393304
rect 349304 393264 350540 393292
rect 349304 393252 349310 393264
rect 350534 393252 350540 393264
rect 350592 393252 350598 393304
rect 350718 393252 350724 393304
rect 350776 393292 350782 393304
rect 350994 393292 351000 393304
rect 350776 393264 351000 393292
rect 350776 393252 350782 393264
rect 350994 393252 351000 393264
rect 351052 393252 351058 393304
rect 353386 393252 353392 393304
rect 353444 393292 353450 393304
rect 354306 393292 354312 393304
rect 353444 393264 354312 393292
rect 353444 393252 353450 393264
rect 354306 393252 354312 393264
rect 354364 393252 354370 393304
rect 359734 393252 359740 393304
rect 359792 393292 359798 393304
rect 360194 393292 360200 393304
rect 359792 393264 360200 393292
rect 359792 393252 359798 393264
rect 360194 393252 360200 393264
rect 360252 393252 360258 393304
rect 364518 393252 364524 393304
rect 364576 393292 364582 393304
rect 364794 393292 364800 393304
rect 364576 393264 364800 393292
rect 364576 393252 364582 393264
rect 364794 393252 364800 393264
rect 364852 393252 364858 393304
rect 365990 393252 365996 393304
rect 366048 393292 366054 393304
rect 366910 393292 366916 393304
rect 366048 393264 366916 393292
rect 366048 393252 366054 393264
rect 366910 393252 366916 393264
rect 366968 393252 366974 393304
rect 367830 393252 367836 393304
rect 367888 393292 367894 393304
rect 370222 393292 370228 393304
rect 367888 393264 370228 393292
rect 367888 393252 367894 393264
rect 370222 393252 370228 393264
rect 370280 393252 370286 393304
rect 341794 393184 341800 393236
rect 341852 393224 341858 393236
rect 386506 393224 386512 393236
rect 341852 393196 386512 393224
rect 341852 393184 341858 393196
rect 386506 393184 386512 393196
rect 386564 393184 386570 393236
rect 341426 393116 341432 393168
rect 341484 393156 341490 393168
rect 366450 393156 366456 393168
rect 341484 393128 366456 393156
rect 341484 393116 341490 393128
rect 366450 393116 366456 393128
rect 366508 393116 366514 393168
rect 373166 393116 373172 393168
rect 373224 393156 373230 393168
rect 373718 393156 373724 393168
rect 373224 393128 373724 393156
rect 373224 393116 373230 393128
rect 373718 393116 373724 393128
rect 373776 393116 373782 393168
rect 336642 393048 336648 393100
rect 336700 393088 336706 393100
rect 364242 393088 364248 393100
rect 336700 393060 364248 393088
rect 336700 393048 336706 393060
rect 364242 393048 364248 393060
rect 364300 393048 364306 393100
rect 364426 393048 364432 393100
rect 364484 393088 364490 393100
rect 364702 393088 364708 393100
rect 364484 393060 364708 393088
rect 364484 393048 364490 393060
rect 364702 393048 364708 393060
rect 364760 393048 364766 393100
rect 364794 393048 364800 393100
rect 364852 393088 364858 393100
rect 365714 393088 365720 393100
rect 364852 393060 365720 393088
rect 364852 393048 364858 393060
rect 365714 393048 365720 393060
rect 365772 393048 365778 393100
rect 315850 392980 315856 393032
rect 315908 393020 315914 393032
rect 375098 393020 375104 393032
rect 315908 392992 375104 393020
rect 315908 392980 315914 392992
rect 375098 392980 375104 392992
rect 375156 392980 375162 393032
rect 282362 392912 282368 392964
rect 282420 392952 282426 392964
rect 342714 392952 342720 392964
rect 282420 392924 342720 392952
rect 282420 392912 282426 392924
rect 342714 392912 342720 392924
rect 342772 392912 342778 392964
rect 343450 392912 343456 392964
rect 343508 392952 343514 392964
rect 345474 392952 345480 392964
rect 343508 392924 345480 392952
rect 343508 392912 343514 392924
rect 345474 392912 345480 392924
rect 345532 392912 345538 392964
rect 346118 392912 346124 392964
rect 346176 392952 346182 392964
rect 350258 392952 350264 392964
rect 346176 392924 350264 392952
rect 346176 392912 346182 392924
rect 350258 392912 350264 392924
rect 350316 392912 350322 392964
rect 358262 392912 358268 392964
rect 358320 392952 358326 392964
rect 358722 392952 358728 392964
rect 358320 392924 358728 392952
rect 358320 392912 358326 392924
rect 358722 392912 358728 392924
rect 358780 392912 358786 392964
rect 359458 392912 359464 392964
rect 359516 392952 359522 392964
rect 364978 392952 364984 392964
rect 359516 392924 364984 392952
rect 359516 392912 359522 392924
rect 364978 392912 364984 392924
rect 365036 392912 365042 392964
rect 279786 392844 279792 392896
rect 279844 392884 279850 392896
rect 345198 392884 345204 392896
rect 279844 392856 345204 392884
rect 279844 392844 279850 392856
rect 345198 392844 345204 392856
rect 345256 392844 345262 392896
rect 349154 392844 349160 392896
rect 349212 392884 349218 392896
rect 349338 392884 349344 392896
rect 349212 392856 349344 392884
rect 349212 392844 349218 392856
rect 349338 392844 349344 392856
rect 349396 392844 349402 392896
rect 363598 392844 363604 392896
rect 363656 392884 363662 392896
rect 366726 392884 366732 392896
rect 363656 392856 366732 392884
rect 363656 392844 363662 392856
rect 366726 392844 366732 392856
rect 366784 392844 366790 392896
rect 276290 392776 276296 392828
rect 276348 392816 276354 392828
rect 350074 392816 350080 392828
rect 276348 392788 350080 392816
rect 276348 392776 276354 392788
rect 350074 392776 350080 392788
rect 350132 392776 350138 392828
rect 370590 392776 370596 392828
rect 370648 392816 370654 392828
rect 370958 392816 370964 392828
rect 370648 392788 370964 392816
rect 370648 392776 370654 392788
rect 370958 392776 370964 392788
rect 371016 392776 371022 392828
rect 347038 392708 347044 392760
rect 347096 392748 347102 392760
rect 348878 392748 348884 392760
rect 347096 392720 348884 392748
rect 347096 392708 347102 392720
rect 348878 392708 348884 392720
rect 348936 392708 348942 392760
rect 352742 392708 352748 392760
rect 352800 392748 352806 392760
rect 381722 392748 381728 392760
rect 352800 392720 381728 392748
rect 352800 392708 352806 392720
rect 381722 392708 381728 392720
rect 381780 392708 381786 392760
rect 274082 392640 274088 392692
rect 274140 392680 274146 392692
rect 353202 392680 353208 392692
rect 274140 392652 353208 392680
rect 274140 392640 274146 392652
rect 353202 392640 353208 392652
rect 353260 392640 353266 392692
rect 271414 392572 271420 392624
rect 271472 392612 271478 392624
rect 363322 392612 363328 392624
rect 271472 392584 363328 392612
rect 271472 392572 271478 392584
rect 363322 392572 363328 392584
rect 363380 392572 363386 392624
rect 371878 392572 371884 392624
rect 371936 392612 371942 392624
rect 382366 392612 382372 392624
rect 371936 392584 382372 392612
rect 371936 392572 371942 392584
rect 382366 392572 382372 392584
rect 382424 392572 382430 392624
rect 330478 392504 330484 392556
rect 330536 392544 330542 392556
rect 343542 392544 343548 392556
rect 330536 392516 343548 392544
rect 330536 392504 330542 392516
rect 343542 392504 343548 392516
rect 343600 392504 343606 392556
rect 359550 392504 359556 392556
rect 359608 392544 359614 392556
rect 360102 392544 360108 392556
rect 359608 392516 360108 392544
rect 359608 392504 359614 392516
rect 360102 392504 360108 392516
rect 360160 392504 360166 392556
rect 271598 392436 271604 392488
rect 271656 392476 271662 392488
rect 361666 392476 361672 392488
rect 271656 392448 361672 392476
rect 271656 392436 271662 392448
rect 361666 392436 361672 392448
rect 361724 392436 361730 392488
rect 344278 392368 344284 392420
rect 344336 392408 344342 392420
rect 353570 392408 353576 392420
rect 344336 392380 353576 392408
rect 344336 392368 344342 392380
rect 353570 392368 353576 392380
rect 353628 392368 353634 392420
rect 375742 392368 375748 392420
rect 375800 392408 375806 392420
rect 376110 392408 376116 392420
rect 375800 392380 376116 392408
rect 375800 392368 375806 392380
rect 376110 392368 376116 392380
rect 376168 392368 376174 392420
rect 365070 392300 365076 392352
rect 365128 392340 365134 392352
rect 369854 392340 369860 392352
rect 365128 392312 369860 392340
rect 365128 392300 365134 392312
rect 369854 392300 369860 392312
rect 369912 392300 369918 392352
rect 367830 392232 367836 392284
rect 367888 392272 367894 392284
rect 368474 392272 368480 392284
rect 367888 392244 368480 392272
rect 367888 392232 367894 392244
rect 368474 392232 368480 392244
rect 368532 392232 368538 392284
rect 355502 392028 355508 392080
rect 355560 392068 355566 392080
rect 364334 392068 364340 392080
rect 355560 392040 364340 392068
rect 355560 392028 355566 392040
rect 364334 392028 364340 392040
rect 364392 392028 364398 392080
rect 364978 391960 364984 392012
rect 365036 392000 365042 392012
rect 370406 392000 370412 392012
rect 365036 391972 370412 392000
rect 365036 391960 365042 391972
rect 370406 391960 370412 391972
rect 370464 391960 370470 392012
rect 360746 391824 360752 391876
rect 360804 391864 360810 391876
rect 361114 391864 361120 391876
rect 360804 391836 361120 391864
rect 360804 391824 360810 391836
rect 361114 391824 361120 391836
rect 361172 391824 361178 391876
rect 367186 391756 367192 391808
rect 367244 391796 367250 391808
rect 369854 391796 369860 391808
rect 367244 391768 369860 391796
rect 367244 391756 367250 391768
rect 369854 391756 369860 391768
rect 369912 391756 369918 391808
rect 311802 391416 311808 391468
rect 311860 391456 311866 391468
rect 371694 391456 371700 391468
rect 311860 391428 371700 391456
rect 311860 391416 311866 391428
rect 371694 391416 371700 391428
rect 371752 391416 371758 391468
rect 281718 391348 281724 391400
rect 281776 391388 281782 391400
rect 342254 391388 342260 391400
rect 281776 391360 342260 391388
rect 281776 391348 281782 391360
rect 342254 391348 342260 391360
rect 342312 391348 342318 391400
rect 344646 391388 344652 391400
rect 343284 391360 344652 391388
rect 270310 391280 270316 391332
rect 270368 391320 270374 391332
rect 343284 391320 343312 391360
rect 344646 391348 344652 391360
rect 344704 391348 344710 391400
rect 381078 391388 381084 391400
rect 350506 391360 381084 391388
rect 270368 391292 343312 391320
rect 270368 391280 270374 391292
rect 343358 391280 343364 391332
rect 343416 391320 343422 391332
rect 350506 391320 350534 391360
rect 381078 391348 381084 391360
rect 381136 391348 381142 391400
rect 343416 391292 350534 391320
rect 343416 391280 343422 391292
rect 368658 391280 368664 391332
rect 368716 391320 368722 391332
rect 369302 391320 369308 391332
rect 368716 391292 369308 391320
rect 368716 391280 368722 391292
rect 369302 391280 369308 391292
rect 369360 391280 369366 391332
rect 369394 391280 369400 391332
rect 369452 391320 369458 391332
rect 371694 391320 371700 391332
rect 369452 391292 371700 391320
rect 369452 391280 369458 391292
rect 371694 391280 371700 391292
rect 371752 391280 371758 391332
rect 267550 391212 267556 391264
rect 267608 391252 267614 391264
rect 348234 391252 348240 391264
rect 267608 391224 348240 391252
rect 267608 391212 267614 391224
rect 348234 391212 348240 391224
rect 348292 391212 348298 391264
rect 359182 391212 359188 391264
rect 359240 391252 359246 391264
rect 359826 391252 359832 391264
rect 359240 391224 359832 391252
rect 359240 391212 359246 391224
rect 359826 391212 359832 391224
rect 359884 391212 359890 391264
rect 363690 391212 363696 391264
rect 363748 391252 363754 391264
rect 383102 391252 383108 391264
rect 363748 391224 383108 391252
rect 363748 391212 363754 391224
rect 383102 391212 383108 391224
rect 383160 391212 383166 391264
rect 374454 391076 374460 391128
rect 374512 391116 374518 391128
rect 374914 391116 374920 391128
rect 374512 391088 374920 391116
rect 374512 391076 374518 391088
rect 374914 391076 374920 391088
rect 374972 391076 374978 391128
rect 341794 391008 341800 391060
rect 341852 391048 341858 391060
rect 354950 391048 354956 391060
rect 341852 391020 354956 391048
rect 341852 391008 341858 391020
rect 354950 391008 354956 391020
rect 355008 391008 355014 391060
rect 313182 390600 313188 390652
rect 313240 390640 313246 390652
rect 372614 390640 372620 390652
rect 313240 390612 372620 390640
rect 313240 390600 313246 390612
rect 372614 390600 372620 390612
rect 372672 390600 372678 390652
rect 314378 390532 314384 390584
rect 314436 390572 314442 390584
rect 373994 390572 374000 390584
rect 314436 390544 374000 390572
rect 314436 390532 314442 390544
rect 373994 390532 374000 390544
rect 374052 390532 374058 390584
rect 345934 390464 345940 390516
rect 345992 390504 345998 390516
rect 375466 390504 375472 390516
rect 345992 390476 375472 390504
rect 345992 390464 345998 390476
rect 375466 390464 375472 390476
rect 375524 390464 375530 390516
rect 356698 390328 356704 390380
rect 356756 390368 356762 390380
rect 360562 390368 360568 390380
rect 356756 390340 360568 390368
rect 356756 390328 356762 390340
rect 360562 390328 360568 390340
rect 360620 390328 360626 390380
rect 337562 390192 337568 390244
rect 337620 390232 337626 390244
rect 345566 390232 345572 390244
rect 337620 390204 345572 390232
rect 337620 390192 337626 390204
rect 345566 390192 345572 390204
rect 345624 390192 345630 390244
rect 319162 390124 319168 390176
rect 319220 390164 319226 390176
rect 379330 390164 379336 390176
rect 319220 390136 379336 390164
rect 319220 390124 319226 390136
rect 379330 390124 379336 390136
rect 379388 390124 379394 390176
rect 319806 390056 319812 390108
rect 319864 390096 319870 390108
rect 378134 390096 378140 390108
rect 319864 390068 378140 390096
rect 319864 390056 319870 390068
rect 378134 390056 378140 390068
rect 378192 390056 378198 390108
rect 319898 389988 319904 390040
rect 319956 390028 319962 390040
rect 380158 390028 380164 390040
rect 319956 390000 380164 390028
rect 319956 389988 319962 390000
rect 380158 389988 380164 390000
rect 380216 389988 380222 390040
rect 281810 389920 281816 389972
rect 281868 389960 281874 389972
rect 342622 389960 342628 389972
rect 281868 389932 342628 389960
rect 281868 389920 281874 389932
rect 342622 389920 342628 389932
rect 342680 389920 342686 389972
rect 343082 389920 343088 389972
rect 343140 389960 343146 389972
rect 367002 389960 367008 389972
rect 343140 389932 367008 389960
rect 343140 389920 343146 389932
rect 367002 389920 367008 389932
rect 367060 389920 367066 389972
rect 269850 389852 269856 389904
rect 269908 389892 269914 389904
rect 342438 389892 342444 389904
rect 269908 389864 342444 389892
rect 269908 389852 269914 389864
rect 342438 389852 342444 389864
rect 342496 389852 342502 389904
rect 259270 389784 259276 389836
rect 259328 389824 259334 389836
rect 347130 389824 347136 389836
rect 259328 389796 347136 389824
rect 259328 389784 259334 389796
rect 347130 389784 347136 389796
rect 347188 389784 347194 389836
rect 351270 389716 351276 389768
rect 351328 389756 351334 389768
rect 361758 389756 361764 389768
rect 351328 389728 361764 389756
rect 351328 389716 351334 389728
rect 361758 389716 361764 389728
rect 361816 389716 361822 389768
rect 347130 389512 347136 389564
rect 347188 389552 347194 389564
rect 354490 389552 354496 389564
rect 347188 389524 354496 389552
rect 347188 389512 347194 389524
rect 354490 389512 354496 389524
rect 354548 389512 354554 389564
rect 349798 389308 349804 389360
rect 349856 389348 349862 389360
rect 355134 389348 355140 389360
rect 349856 389320 355140 389348
rect 349856 389308 349862 389320
rect 355134 389308 355140 389320
rect 355192 389308 355198 389360
rect 318702 389172 318708 389224
rect 318760 389212 318766 389224
rect 378134 389212 378140 389224
rect 318760 389184 378140 389212
rect 318760 389172 318766 389184
rect 378134 389172 378140 389184
rect 378192 389172 378198 389224
rect 350994 388968 351000 389020
rect 351052 389008 351058 389020
rect 351454 389008 351460 389020
rect 351052 388980 351460 389008
rect 351052 388968 351058 388980
rect 351454 388968 351460 388980
rect 351512 388968 351518 389020
rect 333514 388696 333520 388748
rect 333572 388736 333578 388748
rect 365162 388736 365168 388748
rect 333572 388708 365168 388736
rect 333572 388696 333578 388708
rect 365162 388696 365168 388708
rect 365220 388696 365226 388748
rect 343542 388628 343548 388680
rect 343600 388668 343606 388680
rect 383654 388668 383660 388680
rect 343600 388640 383660 388668
rect 343600 388628 343606 388640
rect 383654 388628 383660 388640
rect 383712 388628 383718 388680
rect 276658 388560 276664 388612
rect 276716 388600 276722 388612
rect 343174 388600 343180 388612
rect 276716 388572 343180 388600
rect 276716 388560 276722 388572
rect 343174 388560 343180 388572
rect 343232 388560 343238 388612
rect 262122 388492 262128 388544
rect 262180 388532 262186 388544
rect 348050 388532 348056 388544
rect 262180 388504 348056 388532
rect 262180 388492 262186 388504
rect 348050 388492 348056 388504
rect 348108 388492 348114 388544
rect 349890 388492 349896 388544
rect 349948 388532 349954 388544
rect 381446 388532 381452 388544
rect 349948 388504 381452 388532
rect 349948 388492 349954 388504
rect 381446 388492 381452 388504
rect 381504 388492 381510 388544
rect 257890 388424 257896 388476
rect 257948 388464 257954 388476
rect 347590 388464 347596 388476
rect 257948 388436 347596 388464
rect 257948 388424 257954 388436
rect 347590 388424 347596 388436
rect 347648 388424 347654 388476
rect 354214 388424 354220 388476
rect 354272 388464 354278 388476
rect 386414 388464 386420 388476
rect 354272 388436 386420 388464
rect 354272 388424 354278 388436
rect 386414 388424 386420 388436
rect 386472 388424 386478 388476
rect 356698 388016 356704 388068
rect 356756 388056 356762 388068
rect 356974 388056 356980 388068
rect 356756 388028 356980 388056
rect 356756 388016 356762 388028
rect 356974 388016 356980 388028
rect 357032 388016 357038 388068
rect 352558 387880 352564 387932
rect 352616 387920 352622 387932
rect 354858 387920 354864 387932
rect 352616 387892 354864 387920
rect 352616 387880 352622 387892
rect 354858 387880 354864 387892
rect 354916 387880 354922 387932
rect 321738 387744 321744 387796
rect 321796 387784 321802 387796
rect 322474 387784 322480 387796
rect 321796 387756 322480 387784
rect 321796 387744 321802 387756
rect 322474 387744 322480 387756
rect 322532 387744 322538 387796
rect 348510 387744 348516 387796
rect 348568 387784 348574 387796
rect 355686 387784 355692 387796
rect 348568 387756 355692 387784
rect 348568 387744 348574 387756
rect 355686 387744 355692 387756
rect 355744 387744 355750 387796
rect 348602 387608 348608 387660
rect 348660 387648 348666 387660
rect 357158 387648 357164 387660
rect 348660 387620 357164 387648
rect 348660 387608 348666 387620
rect 357158 387608 357164 387620
rect 357216 387608 357222 387660
rect 331030 387540 331036 387592
rect 331088 387580 331094 387592
rect 355226 387580 355232 387592
rect 331088 387552 355232 387580
rect 331088 387540 331094 387552
rect 355226 387540 355232 387552
rect 355284 387540 355290 387592
rect 305086 387472 305092 387524
rect 305144 387512 305150 387524
rect 305638 387512 305644 387524
rect 305144 387484 305644 387512
rect 305144 387472 305150 387484
rect 305638 387472 305644 387484
rect 305696 387472 305702 387524
rect 329374 387472 329380 387524
rect 329432 387512 329438 387524
rect 365346 387512 365352 387524
rect 329432 387484 365352 387512
rect 329432 387472 329438 387484
rect 365346 387472 365352 387484
rect 365404 387472 365410 387524
rect 333606 387404 333612 387456
rect 333664 387444 333670 387456
rect 373442 387444 373448 387456
rect 333664 387416 373448 387444
rect 333664 387404 333670 387416
rect 373442 387404 373448 387416
rect 373500 387404 373506 387456
rect 332410 387336 332416 387388
rect 332468 387376 332474 387388
rect 374822 387376 374828 387388
rect 332468 387348 374828 387376
rect 332468 387336 332474 387348
rect 374822 387336 374828 387348
rect 374880 387336 374886 387388
rect 329466 387268 329472 387320
rect 329524 387308 329530 387320
rect 371970 387308 371976 387320
rect 329524 387280 371976 387308
rect 329524 387268 329530 387280
rect 371970 387268 371976 387280
rect 372028 387268 372034 387320
rect 275462 387200 275468 387252
rect 275520 387240 275526 387252
rect 341242 387240 341248 387252
rect 275520 387212 341248 387240
rect 275520 387200 275526 387212
rect 341242 387200 341248 387212
rect 341300 387200 341306 387252
rect 347314 387200 347320 387252
rect 347372 387240 347378 387252
rect 359366 387240 359372 387252
rect 347372 387212 359372 387240
rect 347372 387200 347378 387212
rect 359366 387200 359372 387212
rect 359424 387200 359430 387252
rect 263410 387132 263416 387184
rect 263468 387172 263474 387184
rect 342806 387172 342812 387184
rect 263468 387144 342812 387172
rect 263468 387132 263474 387144
rect 342806 387132 342812 387144
rect 342864 387132 342870 387184
rect 344554 387132 344560 387184
rect 344612 387172 344618 387184
rect 357710 387172 357716 387184
rect 344612 387144 357716 387172
rect 344612 387132 344618 387144
rect 357710 387132 357716 387144
rect 357768 387132 357774 387184
rect 275370 387064 275376 387116
rect 275428 387104 275434 387116
rect 363506 387104 363512 387116
rect 275428 387076 363512 387104
rect 275428 387064 275434 387076
rect 363506 387064 363512 387076
rect 363564 387064 363570 387116
rect 262858 386452 262864 386504
rect 262916 386492 262922 386504
rect 321738 386492 321744 386504
rect 262916 386464 321744 386492
rect 262916 386452 262922 386464
rect 321738 386452 321744 386464
rect 321796 386452 321802 386504
rect 279142 386384 279148 386436
rect 279200 386424 279206 386436
rect 292574 386424 292580 386436
rect 279200 386396 292580 386424
rect 279200 386384 279206 386396
rect 292574 386384 292580 386396
rect 292632 386424 292638 386436
rect 293862 386424 293868 386436
rect 292632 386396 293868 386424
rect 292632 386384 292638 386396
rect 293862 386384 293868 386396
rect 293920 386424 293926 386436
rect 580258 386424 580264 386436
rect 293920 386396 580264 386424
rect 293920 386384 293926 386396
rect 580258 386384 580264 386396
rect 580316 386384 580322 386436
rect 320450 386316 320456 386368
rect 320508 386356 320514 386368
rect 320910 386356 320916 386368
rect 320508 386328 320916 386356
rect 320508 386316 320514 386328
rect 320910 386316 320916 386328
rect 320968 386316 320974 386368
rect 277854 385976 277860 386028
rect 277912 386016 277918 386028
rect 349982 386016 349988 386028
rect 277912 385988 349988 386016
rect 277912 385976 277918 385988
rect 349982 385976 349988 385988
rect 350040 385976 350046 386028
rect 280706 385908 280712 385960
rect 280764 385948 280770 385960
rect 358354 385948 358360 385960
rect 280764 385920 358360 385948
rect 280764 385908 280770 385920
rect 358354 385908 358360 385920
rect 358412 385908 358418 385960
rect 279510 385840 279516 385892
rect 279568 385880 279574 385892
rect 360746 385880 360752 385892
rect 279568 385852 360752 385880
rect 279568 385840 279574 385852
rect 360746 385840 360752 385852
rect 360804 385840 360810 385892
rect 268930 385772 268936 385824
rect 268988 385812 268994 385824
rect 353018 385812 353024 385824
rect 268988 385784 353024 385812
rect 268988 385772 268994 385784
rect 353018 385772 353024 385784
rect 353076 385772 353082 385824
rect 279602 385704 279608 385756
rect 279660 385744 279666 385756
rect 368106 385744 368112 385756
rect 279660 385716 368112 385744
rect 279660 385704 279666 385716
rect 368106 385704 368112 385716
rect 368164 385704 368170 385756
rect 3418 385636 3424 385688
rect 3476 385676 3482 385688
rect 255314 385676 255320 385688
rect 3476 385648 255320 385676
rect 3476 385636 3482 385648
rect 255314 385636 255320 385648
rect 255372 385636 255378 385688
rect 278222 385636 278228 385688
rect 278280 385676 278286 385688
rect 366358 385676 366364 385688
rect 278280 385648 366364 385676
rect 278280 385636 278286 385648
rect 366358 385636 366364 385648
rect 366416 385636 366422 385688
rect 269942 385160 269948 385212
rect 270000 385200 270006 385212
rect 320450 385200 320456 385212
rect 270000 385172 320456 385200
rect 270000 385160 270006 385172
rect 320450 385160 320456 385172
rect 320508 385160 320514 385212
rect 264514 385092 264520 385144
rect 264572 385132 264578 385144
rect 323762 385132 323768 385144
rect 264572 385104 323768 385132
rect 264572 385092 264578 385104
rect 323762 385092 323768 385104
rect 323820 385092 323826 385144
rect 255314 385024 255320 385076
rect 255372 385064 255378 385076
rect 316218 385064 316224 385076
rect 255372 385036 316224 385064
rect 255372 385024 255378 385036
rect 316218 385024 316224 385036
rect 316276 385064 316282 385076
rect 316678 385064 316684 385076
rect 316276 385036 316684 385064
rect 316276 385024 316282 385036
rect 316678 385024 316684 385036
rect 316736 385024 316742 385076
rect 319070 384956 319076 385008
rect 319128 384996 319134 385008
rect 319714 384996 319720 385008
rect 319128 384968 319720 384996
rect 319128 384956 319134 384968
rect 319714 384956 319720 384968
rect 319772 384956 319778 385008
rect 325694 384956 325700 385008
rect 325752 384996 325758 385008
rect 326338 384996 326344 385008
rect 325752 384968 326344 384996
rect 325752 384956 325758 384968
rect 326338 384956 326344 384968
rect 326396 384956 326402 385008
rect 344462 384956 344468 385008
rect 344520 384996 344526 385008
rect 358262 384996 358268 385008
rect 344520 384968 358268 384996
rect 344520 384956 344526 384968
rect 358262 384956 358268 384968
rect 358320 384956 358326 385008
rect 345934 384888 345940 384940
rect 345992 384928 345998 384940
rect 361206 384928 361212 384940
rect 345992 384900 361212 384928
rect 345992 384888 345998 384900
rect 361206 384888 361212 384900
rect 361264 384888 361270 384940
rect 348694 384820 348700 384872
rect 348752 384860 348758 384872
rect 363230 384860 363236 384872
rect 348752 384832 363236 384860
rect 348752 384820 348758 384832
rect 363230 384820 363236 384832
rect 363288 384820 363294 384872
rect 346210 384752 346216 384804
rect 346268 384792 346274 384804
rect 361850 384792 361856 384804
rect 346268 384764 361856 384792
rect 346268 384752 346274 384764
rect 361850 384752 361856 384764
rect 361908 384752 361914 384804
rect 344830 384684 344836 384736
rect 344888 384724 344894 384736
rect 362402 384724 362408 384736
rect 344888 384696 362408 384724
rect 344888 384684 344894 384696
rect 362402 384684 362408 384696
rect 362460 384684 362466 384736
rect 343174 384616 343180 384668
rect 343232 384656 343238 384668
rect 363138 384656 363144 384668
rect 343232 384628 363144 384656
rect 343232 384616 343238 384628
rect 363138 384616 363144 384628
rect 363196 384616 363202 384668
rect 345842 384548 345848 384600
rect 345900 384588 345906 384600
rect 366082 384588 366088 384600
rect 345900 384560 366088 384588
rect 345900 384548 345906 384560
rect 366082 384548 366088 384560
rect 366140 384548 366146 384600
rect 347406 384480 347412 384532
rect 347464 384520 347470 384532
rect 370682 384520 370688 384532
rect 347464 384492 370688 384520
rect 347464 384480 347470 384492
rect 370682 384480 370688 384492
rect 370740 384480 370746 384532
rect 338666 384412 338672 384464
rect 338724 384452 338730 384464
rect 364702 384452 364708 384464
rect 338724 384424 364708 384452
rect 338724 384412 338730 384424
rect 364702 384412 364708 384424
rect 364760 384412 364766 384464
rect 329190 384344 329196 384396
rect 329248 384384 329254 384396
rect 379974 384384 379980 384396
rect 329248 384356 379980 384384
rect 329248 384344 329254 384356
rect 379974 384344 379980 384356
rect 380032 384344 380038 384396
rect 283558 384276 283564 384328
rect 283616 384316 283622 384328
rect 352834 384316 352840 384328
rect 283616 384288 352840 384316
rect 283616 384276 283622 384288
rect 352834 384276 352840 384288
rect 352892 384276 352898 384328
rect 262950 383800 262956 383852
rect 263008 383840 263014 383852
rect 322290 383840 322296 383852
rect 263008 383812 322296 383840
rect 263008 383800 263014 383812
rect 322290 383800 322296 383812
rect 322348 383800 322354 383852
rect 265894 383732 265900 383784
rect 265952 383772 265958 383784
rect 325694 383772 325700 383784
rect 265952 383744 325700 383772
rect 265952 383732 265958 383744
rect 325694 383732 325700 383744
rect 325752 383732 325758 383784
rect 257338 383664 257344 383716
rect 257396 383704 257402 383716
rect 319070 383704 319076 383716
rect 257396 383676 319076 383704
rect 257396 383664 257402 383676
rect 319070 383664 319076 383676
rect 319128 383664 319134 383716
rect 313918 383596 313924 383648
rect 313976 383636 313982 383648
rect 314194 383636 314200 383648
rect 313976 383608 314200 383636
rect 313976 383596 313982 383608
rect 314194 383596 314200 383608
rect 314252 383596 314258 383648
rect 314838 383052 314844 383104
rect 314896 383092 314902 383104
rect 315482 383092 315488 383104
rect 314896 383064 315488 383092
rect 314896 383052 314902 383064
rect 315482 383052 315488 383064
rect 315540 383052 315546 383104
rect 318886 382984 318892 383036
rect 318944 383024 318950 383036
rect 319622 383024 319628 383036
rect 318944 382996 319628 383024
rect 318944 382984 318950 382996
rect 319622 382984 319628 382996
rect 319680 382984 319686 383036
rect 318978 382576 318984 382628
rect 319036 382616 319042 382628
rect 319530 382616 319536 382628
rect 319036 382588 319536 382616
rect 319036 382576 319042 382588
rect 319530 382576 319536 382588
rect 319588 382576 319594 382628
rect 272518 382508 272524 382560
rect 272576 382548 272582 382560
rect 321646 382548 321652 382560
rect 272576 382520 321652 382548
rect 272576 382508 272582 382520
rect 321646 382508 321652 382520
rect 321704 382548 321710 382560
rect 322382 382548 322388 382560
rect 321704 382520 322388 382548
rect 321704 382508 321710 382520
rect 322382 382508 322388 382520
rect 322440 382508 322446 382560
rect 265710 382440 265716 382492
rect 265768 382480 265774 382492
rect 318886 382480 318892 382492
rect 265768 382452 318892 382480
rect 265768 382440 265774 382452
rect 318886 382440 318892 382452
rect 318944 382440 318950 382492
rect 253198 382372 253204 382424
rect 253256 382412 253262 382424
rect 313458 382412 313464 382424
rect 253256 382384 313464 382412
rect 253256 382372 253262 382384
rect 313458 382372 313464 382384
rect 313516 382372 313522 382424
rect 258718 382304 258724 382356
rect 258776 382344 258782 382356
rect 318978 382344 318984 382356
rect 258776 382316 318984 382344
rect 258776 382304 258782 382316
rect 318978 382304 318984 382316
rect 319036 382304 319042 382356
rect 254578 382236 254584 382288
rect 254636 382276 254642 382288
rect 314838 382276 314844 382288
rect 254636 382248 314844 382276
rect 254636 382236 254642 382248
rect 314838 382236 314844 382248
rect 314896 382236 314902 382288
rect 324406 381964 324412 382016
rect 324464 382004 324470 382016
rect 324958 382004 324964 382016
rect 324464 381976 324964 382004
rect 324464 381964 324470 381976
rect 324958 381964 324964 381976
rect 325016 381964 325022 382016
rect 343266 381624 343272 381676
rect 343324 381664 343330 381676
rect 358998 381664 359004 381676
rect 343324 381636 359004 381664
rect 343324 381624 343330 381636
rect 358998 381624 359004 381636
rect 359056 381624 359062 381676
rect 345750 381556 345756 381608
rect 345808 381596 345814 381608
rect 368750 381596 368756 381608
rect 345808 381568 368756 381596
rect 345808 381556 345814 381568
rect 368750 381556 368756 381568
rect 368808 381556 368814 381608
rect 350166 381488 350172 381540
rect 350224 381528 350230 381540
rect 374270 381528 374276 381540
rect 350224 381500 374276 381528
rect 350224 381488 350230 381500
rect 374270 381488 374276 381500
rect 374328 381488 374334 381540
rect 279418 381148 279424 381200
rect 279476 381188 279482 381200
rect 317506 381188 317512 381200
rect 279476 381160 317512 381188
rect 279476 381148 279482 381160
rect 317506 381148 317512 381160
rect 317564 381188 317570 381200
rect 318242 381188 318248 381200
rect 317564 381160 318248 381188
rect 317564 381148 317570 381160
rect 318242 381148 318248 381160
rect 318300 381148 318306 381200
rect 261478 381080 261484 381132
rect 261536 381120 261542 381132
rect 311250 381120 311256 381132
rect 261536 381092 311256 381120
rect 261536 381080 261542 381092
rect 311250 381080 311256 381092
rect 311308 381080 311314 381132
rect 268378 381012 268384 381064
rect 268436 381052 268442 381064
rect 268436 381024 324636 381052
rect 268436 381012 268442 381024
rect 246298 380944 246304 380996
rect 246356 380984 246362 380996
rect 305086 380984 305092 380996
rect 246356 380956 305092 380984
rect 246356 380944 246362 380956
rect 305086 380944 305092 380956
rect 305144 380944 305150 380996
rect 324608 380928 324636 381024
rect 264330 380876 264336 380928
rect 264388 380916 264394 380928
rect 324406 380916 324412 380928
rect 264388 380888 324412 380916
rect 264388 380876 264394 380888
rect 324406 380876 324412 380888
rect 324464 380876 324470 380928
rect 324590 380876 324596 380928
rect 324648 380916 324654 380928
rect 325050 380916 325056 380928
rect 324648 380888 325056 380916
rect 324648 380876 324654 380888
rect 325050 380876 325056 380888
rect 325108 380876 325114 380928
rect 250530 379856 250536 379908
rect 250588 379896 250594 379908
rect 309134 379896 309140 379908
rect 250588 379868 309140 379896
rect 250588 379856 250594 379868
rect 309134 379856 309140 379868
rect 309192 379896 309198 379908
rect 309318 379896 309324 379908
rect 309192 379868 309324 379896
rect 309192 379856 309198 379868
rect 309318 379856 309324 379868
rect 309376 379856 309382 379908
rect 254762 379788 254768 379840
rect 254820 379828 254826 379840
rect 314746 379828 314752 379840
rect 254820 379800 314752 379828
rect 254820 379788 254826 379800
rect 314746 379788 314752 379800
rect 314804 379788 314810 379840
rect 246390 379720 246396 379772
rect 246448 379760 246454 379772
rect 306374 379760 306380 379772
rect 246448 379732 306380 379760
rect 246448 379720 246454 379732
rect 306374 379720 306380 379732
rect 306432 379760 306438 379772
rect 306558 379760 306564 379772
rect 306432 379732 306564 379760
rect 306432 379720 306438 379732
rect 306558 379720 306564 379732
rect 306616 379720 306622 379772
rect 255958 379652 255964 379704
rect 256016 379692 256022 379704
rect 316126 379692 316132 379704
rect 256016 379664 316132 379692
rect 256016 379652 256022 379664
rect 316126 379652 316132 379664
rect 316184 379652 316190 379704
rect 243538 379584 243544 379636
rect 243596 379624 243602 379636
rect 303614 379624 303620 379636
rect 243596 379596 303620 379624
rect 243596 379584 243602 379596
rect 303614 379584 303620 379596
rect 303672 379584 303678 379636
rect 259822 379516 259828 379568
rect 259880 379556 259886 379568
rect 320358 379556 320364 379568
rect 259880 379528 320364 379556
rect 259880 379516 259886 379528
rect 320358 379516 320364 379528
rect 320416 379556 320422 379568
rect 321002 379556 321008 379568
rect 320416 379528 321008 379556
rect 320416 379516 320422 379528
rect 321002 379516 321008 379528
rect 321060 379516 321066 379568
rect 335326 379052 345014 379080
rect 317598 378972 317604 379024
rect 317656 379012 317662 379024
rect 318150 379012 318156 379024
rect 317656 378984 318156 379012
rect 317656 378972 317662 378984
rect 318150 378972 318156 378984
rect 318208 378972 318214 379024
rect 286778 378836 286784 378888
rect 286836 378876 286842 378888
rect 335326 378876 335354 379052
rect 341978 378972 341984 379024
rect 342036 378972 342042 379024
rect 286836 378848 335354 378876
rect 286836 378836 286842 378848
rect 307662 378768 307668 378820
rect 307720 378808 307726 378820
rect 307720 378780 335354 378808
rect 307720 378768 307726 378780
rect 335326 378672 335354 378780
rect 341996 378740 342024 378972
rect 344986 378876 345014 379052
rect 345290 378876 345296 378888
rect 344986 378848 345296 378876
rect 345290 378836 345296 378848
rect 345348 378836 345354 378888
rect 367370 378808 367376 378820
rect 344986 378780 367376 378808
rect 342070 378740 342076 378752
rect 341996 378712 342076 378740
rect 342070 378700 342076 378712
rect 342128 378700 342134 378752
rect 344986 378672 345014 378780
rect 367370 378768 367376 378780
rect 367428 378768 367434 378820
rect 335326 378644 345014 378672
rect 317506 378360 317512 378412
rect 317564 378400 317570 378412
rect 317966 378400 317972 378412
rect 317564 378372 317972 378400
rect 317564 378360 317570 378372
rect 317966 378360 317972 378372
rect 318024 378360 318030 378412
rect 259178 378292 259184 378344
rect 259236 378332 259242 378344
rect 317598 378332 317604 378344
rect 259236 378304 317604 378332
rect 259236 378292 259242 378304
rect 317598 378292 317604 378304
rect 317656 378292 317662 378344
rect 253842 378224 253848 378276
rect 253900 378264 253906 378276
rect 314102 378264 314108 378276
rect 253900 378236 314108 378264
rect 253900 378224 253906 378236
rect 314102 378224 314108 378236
rect 314160 378224 314166 378276
rect 262214 378156 262220 378208
rect 262272 378196 262278 378208
rect 322934 378196 322940 378208
rect 262272 378168 322940 378196
rect 262272 378156 262278 378168
rect 322934 378156 322940 378168
rect 322992 378196 322998 378208
rect 323670 378196 323676 378208
rect 322992 378168 323676 378196
rect 322992 378156 322998 378168
rect 323670 378156 323676 378168
rect 323728 378156 323734 378208
rect 301958 377408 301964 377460
rect 302016 377448 302022 377460
rect 337286 377448 337292 377460
rect 302016 377420 337292 377448
rect 302016 377408 302022 377420
rect 337286 377408 337292 377420
rect 337344 377408 337350 377460
rect 351454 377408 351460 377460
rect 351512 377448 351518 377460
rect 359274 377448 359280 377460
rect 351512 377420 359280 377448
rect 351512 377408 351518 377420
rect 359274 377408 359280 377420
rect 359332 377408 359338 377460
rect 250438 376864 250444 376916
rect 250496 376904 250502 376916
rect 302602 376904 302608 376916
rect 250496 376876 302608 376904
rect 250496 376864 250502 376876
rect 302602 376864 302608 376876
rect 302660 376904 302666 376916
rect 302878 376904 302884 376916
rect 302660 376876 302884 376904
rect 302660 376864 302666 376876
rect 302878 376864 302884 376876
rect 302936 376864 302942 376916
rect 263042 376796 263048 376848
rect 263100 376836 263106 376848
rect 323578 376836 323584 376848
rect 263100 376808 323584 376836
rect 263100 376796 263106 376808
rect 323578 376796 323584 376808
rect 323636 376836 323642 376848
rect 323854 376836 323860 376848
rect 323636 376808 323860 376836
rect 323636 376796 323642 376808
rect 323854 376796 323860 376808
rect 323912 376796 323918 376848
rect 254670 376728 254676 376780
rect 254728 376768 254734 376780
rect 315390 376768 315396 376780
rect 254728 376740 315396 376768
rect 254728 376728 254734 376740
rect 315390 376728 315396 376740
rect 315448 376728 315454 376780
rect 261570 376048 261576 376100
rect 261628 376088 261634 376100
rect 300302 376088 300308 376100
rect 261628 376060 300308 376088
rect 261628 376048 261634 376060
rect 300302 376048 300308 376060
rect 300360 376048 300366 376100
rect 267182 375980 267188 376032
rect 267240 376020 267246 376032
rect 310882 376020 310888 376032
rect 267240 375992 310888 376020
rect 267240 375980 267246 375992
rect 310882 375980 310888 375992
rect 310940 375980 310946 376032
rect 267090 375912 267096 375964
rect 267148 375952 267154 375964
rect 312170 375952 312176 375964
rect 267148 375924 312176 375952
rect 267148 375912 267154 375924
rect 312170 375912 312176 375924
rect 312228 375912 312234 375964
rect 264238 375844 264244 375896
rect 264296 375884 264302 375896
rect 312814 375884 312820 375896
rect 264296 375856 312820 375884
rect 264296 375844 264302 375856
rect 312814 375844 312820 375856
rect 312872 375844 312878 375896
rect 232498 375776 232504 375828
rect 232556 375816 232562 375828
rect 291838 375816 291844 375828
rect 232556 375788 291844 375816
rect 232556 375776 232562 375788
rect 291838 375776 291844 375788
rect 291896 375816 291902 375828
rect 292298 375816 292304 375828
rect 291896 375788 292304 375816
rect 291896 375776 291902 375788
rect 292298 375776 292304 375788
rect 292356 375776 292362 375828
rect 235258 375708 235264 375760
rect 235316 375748 235322 375760
rect 294414 375748 294420 375760
rect 235316 375720 294420 375748
rect 235316 375708 235322 375720
rect 294414 375708 294420 375720
rect 294472 375748 294478 375760
rect 294690 375748 294696 375760
rect 294472 375720 294696 375748
rect 294472 375708 294478 375720
rect 294690 375708 294696 375720
rect 294748 375708 294754 375760
rect 237374 375640 237380 375692
rect 237432 375680 237438 375692
rect 297450 375680 297456 375692
rect 237432 375652 297456 375680
rect 237432 375640 237438 375652
rect 297450 375640 297456 375652
rect 297508 375640 297514 375692
rect 240134 375572 240140 375624
rect 240192 375612 240198 375624
rect 300394 375612 300400 375624
rect 240192 375584 300400 375612
rect 240192 375572 240198 375584
rect 300394 375572 300400 375584
rect 300452 375572 300458 375624
rect 261662 375504 261668 375556
rect 261720 375544 261726 375556
rect 321830 375544 321836 375556
rect 261720 375516 321836 375544
rect 261720 375504 261726 375516
rect 321830 375504 321836 375516
rect 321888 375544 321894 375556
rect 322198 375544 322204 375556
rect 321888 375516 322204 375544
rect 321888 375504 321894 375516
rect 322198 375504 322204 375516
rect 322256 375504 322262 375556
rect 236638 375436 236644 375488
rect 236696 375476 236702 375488
rect 297542 375476 297548 375488
rect 236696 375448 297548 375476
rect 236696 375436 236702 375448
rect 297542 375436 297548 375448
rect 297600 375436 297606 375488
rect 220722 375368 220728 375420
rect 220780 375408 220786 375420
rect 291746 375408 291752 375420
rect 220780 375380 291752 375408
rect 220780 375368 220786 375380
rect 291746 375368 291752 375380
rect 291804 375408 291810 375420
rect 291930 375408 291936 375420
rect 291804 375380 291936 375408
rect 291804 375368 291810 375380
rect 291930 375368 291936 375380
rect 291988 375368 291994 375420
rect 297450 375368 297456 375420
rect 297508 375408 297514 375420
rect 297726 375408 297732 375420
rect 297508 375380 297732 375408
rect 297508 375368 297514 375380
rect 297726 375368 297732 375380
rect 297784 375368 297790 375420
rect 281166 375300 281172 375352
rect 281224 375340 281230 375352
rect 281442 375340 281448 375352
rect 281224 375312 281448 375340
rect 281224 375300 281230 375312
rect 281442 375300 281448 375312
rect 281500 375300 281506 375352
rect 258810 374960 258816 375012
rect 258868 375000 258874 375012
rect 298370 375000 298376 375012
rect 258868 374972 298376 375000
rect 258868 374960 258874 374972
rect 298370 374960 298376 374972
rect 298428 374960 298434 375012
rect 259546 374892 259552 374944
rect 259604 374932 259610 374944
rect 319530 374932 319536 374944
rect 259604 374904 319536 374932
rect 259604 374892 259610 374904
rect 319530 374892 319536 374904
rect 319588 374892 319594 374944
rect 281166 374756 281172 374808
rect 281224 374796 281230 374808
rect 307294 374796 307300 374808
rect 281224 374768 307300 374796
rect 281224 374756 281230 374768
rect 307294 374756 307300 374768
rect 307352 374756 307358 374808
rect 275646 374688 275652 374740
rect 275704 374728 275710 374740
rect 300854 374728 300860 374740
rect 275704 374700 300860 374728
rect 275704 374688 275710 374700
rect 300854 374688 300860 374700
rect 300912 374728 300918 374740
rect 301590 374728 301596 374740
rect 300912 374700 301596 374728
rect 300912 374688 300918 374700
rect 301590 374688 301596 374700
rect 301648 374688 301654 374740
rect 220078 374620 220084 374672
rect 220136 374660 220142 374672
rect 281994 374660 282000 374672
rect 220136 374632 282000 374660
rect 220136 374620 220142 374632
rect 281994 374620 282000 374632
rect 282052 374620 282058 374672
rect 314746 374620 314752 374672
rect 314804 374660 314810 374672
rect 315390 374660 315396 374672
rect 314804 374632 315396 374660
rect 314804 374620 314810 374632
rect 315390 374620 315396 374632
rect 315448 374620 315454 374672
rect 321646 374620 321652 374672
rect 321704 374660 321710 374672
rect 322382 374660 322388 374672
rect 321704 374632 322388 374660
rect 321704 374620 321710 374632
rect 322382 374620 322388 374632
rect 322440 374620 322446 374672
rect 324406 374620 324412 374672
rect 324464 374660 324470 374672
rect 324958 374660 324964 374672
rect 324464 374632 324964 374660
rect 324464 374620 324470 374632
rect 324958 374620 324964 374632
rect 325016 374620 325022 374672
rect 273162 374552 273168 374604
rect 273220 374592 273226 374604
rect 301958 374592 301964 374604
rect 273220 374564 301964 374592
rect 273220 374552 273226 374564
rect 301958 374552 301964 374564
rect 302016 374552 302022 374604
rect 264606 374484 264612 374536
rect 264664 374524 264670 374536
rect 294782 374524 294788 374536
rect 264664 374496 294788 374524
rect 264664 374484 264670 374496
rect 294782 374484 294788 374496
rect 294840 374484 294846 374536
rect 305546 374484 305552 374536
rect 305604 374524 305610 374536
rect 305730 374524 305736 374536
rect 305604 374496 305736 374524
rect 305604 374484 305610 374496
rect 305730 374484 305736 374496
rect 305788 374484 305794 374536
rect 272794 374416 272800 374468
rect 272852 374456 272858 374468
rect 304350 374456 304356 374468
rect 272852 374428 304356 374456
rect 272852 374416 272858 374428
rect 304350 374416 304356 374428
rect 304408 374416 304414 374468
rect 264422 374348 264428 374400
rect 264480 374388 264486 374400
rect 297082 374388 297088 374400
rect 264480 374360 297088 374388
rect 264480 374348 264486 374360
rect 297082 374348 297088 374360
rect 297140 374348 297146 374400
rect 274542 374280 274548 374332
rect 274600 374320 274606 374332
rect 308398 374320 308404 374332
rect 274600 374292 308404 374320
rect 274600 374280 274606 374292
rect 308398 374280 308404 374292
rect 308456 374280 308462 374332
rect 272702 374212 272708 374264
rect 272760 374252 272766 374264
rect 307018 374252 307024 374264
rect 272760 374224 307024 374252
rect 272760 374212 272766 374224
rect 307018 374212 307024 374224
rect 307076 374212 307082 374264
rect 267274 374144 267280 374196
rect 267332 374184 267338 374196
rect 305546 374184 305552 374196
rect 267332 374156 305552 374184
rect 267332 374144 267338 374156
rect 305546 374144 305552 374156
rect 305604 374144 305610 374196
rect 290182 374116 290188 374128
rect 277366 374088 290188 374116
rect 277366 374060 277394 374088
rect 290182 374076 290188 374088
rect 290240 374076 290246 374128
rect 295518 374076 295524 374128
rect 295576 374116 295582 374128
rect 300118 374116 300124 374128
rect 295576 374088 300124 374116
rect 295576 374076 295582 374088
rect 300118 374076 300124 374088
rect 300176 374076 300182 374128
rect 277302 374008 277308 374060
rect 277360 374020 277394 374060
rect 277360 374008 277366 374020
rect 278498 374008 278504 374060
rect 278556 374048 278562 374060
rect 283558 374048 283564 374060
rect 278556 374020 283564 374048
rect 278556 374008 278562 374020
rect 283558 374008 283564 374020
rect 283616 374008 283622 374060
rect 153194 373940 153200 373992
rect 153252 373980 153258 373992
rect 282270 373980 282276 373992
rect 153252 373952 282276 373980
rect 153252 373940 153258 373952
rect 282270 373940 282276 373952
rect 282328 373940 282334 373992
rect 304810 373940 304816 373992
rect 304868 373980 304874 373992
rect 309778 373980 309784 373992
rect 304868 373952 309784 373980
rect 304868 373940 304874 373952
rect 309778 373940 309784 373952
rect 309836 373940 309842 373992
rect 277946 373464 277952 373516
rect 278004 373504 278010 373516
rect 281442 373504 281448 373516
rect 278004 373476 281448 373504
rect 278004 373464 278010 373476
rect 281442 373464 281448 373476
rect 281500 373464 281506 373516
rect 294322 373464 294328 373516
rect 294380 373504 294386 373516
rect 294782 373504 294788 373516
rect 294380 373476 294788 373504
rect 294380 373464 294386 373476
rect 294782 373464 294788 373476
rect 294840 373464 294846 373516
rect 278774 373396 278780 373448
rect 278832 373436 278838 373448
rect 278832 373408 289814 373436
rect 278832 373396 278838 373408
rect 278314 373328 278320 373380
rect 278372 373368 278378 373380
rect 287422 373368 287428 373380
rect 278372 373340 287428 373368
rect 278372 373328 278378 373340
rect 287422 373328 287428 373340
rect 287480 373328 287486 373380
rect 226978 373260 226984 373312
rect 227036 373300 227042 373312
rect 278590 373300 278596 373312
rect 227036 373272 278596 373300
rect 227036 373260 227042 373272
rect 278590 373260 278596 373272
rect 278648 373300 278654 373312
rect 288526 373300 288532 373312
rect 278648 373272 288532 373300
rect 278648 373260 278654 373272
rect 288526 373260 288532 373272
rect 288584 373260 288590 373312
rect 289786 373300 289814 373408
rect 298462 373396 298468 373448
rect 298520 373436 298526 373448
rect 337930 373436 337936 373448
rect 298520 373408 337936 373436
rect 298520 373396 298526 373408
rect 337930 373396 337936 373408
rect 337988 373396 337994 373448
rect 295610 373328 295616 373380
rect 295668 373368 295674 373380
rect 297542 373368 297548 373380
rect 295668 373340 297548 373368
rect 295668 373328 295674 373340
rect 297542 373328 297548 373340
rect 297600 373368 297606 373380
rect 340690 373368 340696 373380
rect 297600 373340 340696 373368
rect 297600 373328 297606 373340
rect 340690 373328 340696 373340
rect 340748 373328 340754 373380
rect 296622 373300 296628 373312
rect 289786 373272 296628 373300
rect 296622 373260 296628 373272
rect 296680 373300 296686 373312
rect 340046 373300 340052 373312
rect 296680 373272 340052 373300
rect 296680 373260 296686 373272
rect 340046 373260 340052 373272
rect 340104 373260 340110 373312
rect 220354 373192 220360 373244
rect 220412 373232 220418 373244
rect 282178 373232 282184 373244
rect 220412 373204 282184 373232
rect 220412 373192 220418 373204
rect 282178 373192 282184 373204
rect 282236 373232 282242 373244
rect 286502 373232 286508 373244
rect 282236 373204 286508 373232
rect 282236 373192 282242 373204
rect 286502 373192 286508 373204
rect 286560 373192 286566 373244
rect 278590 373124 278596 373176
rect 278648 373164 278654 373176
rect 278774 373164 278780 373176
rect 278648 373136 278780 373164
rect 278648 373124 278654 373136
rect 278774 373124 278780 373136
rect 278832 373124 278838 373176
rect 295518 373164 295524 373176
rect 281184 373136 295524 373164
rect 278130 373056 278136 373108
rect 278188 373096 278194 373108
rect 281184 373096 281212 373136
rect 295518 373124 295524 373136
rect 295576 373124 295582 373176
rect 278188 373068 281212 373096
rect 278188 373056 278194 373068
rect 281442 373056 281448 373108
rect 281500 373096 281506 373108
rect 298462 373096 298468 373108
rect 281500 373068 298468 373096
rect 281500 373056 281506 373068
rect 298462 373056 298468 373068
rect 298520 373056 298526 373108
rect 275830 372988 275836 373040
rect 275888 373028 275894 373040
rect 295610 373028 295616 373040
rect 275888 373000 295616 373028
rect 275888 372988 275894 373000
rect 295610 372988 295616 373000
rect 295668 372988 295674 373040
rect 275186 372920 275192 372972
rect 275244 372960 275250 372972
rect 300210 372960 300216 372972
rect 275244 372932 300216 372960
rect 275244 372920 275250 372932
rect 300210 372920 300216 372932
rect 300268 372920 300274 372972
rect 267458 372852 267464 372904
rect 267516 372892 267522 372904
rect 301314 372892 301320 372904
rect 267516 372864 301320 372892
rect 267516 372852 267522 372864
rect 301314 372852 301320 372864
rect 301372 372852 301378 372904
rect 244918 372784 244924 372836
rect 244976 372824 244982 372836
rect 304810 372824 304816 372836
rect 244976 372796 304816 372824
rect 244976 372784 244982 372796
rect 304810 372784 304816 372796
rect 304868 372784 304874 372836
rect 238110 372716 238116 372768
rect 238168 372756 238174 372768
rect 299198 372756 299204 372768
rect 238168 372728 299204 372756
rect 238168 372716 238174 372728
rect 299198 372716 299204 372728
rect 299256 372716 299262 372768
rect 273070 372648 273076 372700
rect 273128 372688 273134 372700
rect 303430 372688 303436 372700
rect 273128 372660 303436 372688
rect 273128 372648 273134 372660
rect 303430 372648 303436 372660
rect 303488 372648 303494 372700
rect 306926 372648 306932 372700
rect 306984 372688 306990 372700
rect 308490 372688 308496 372700
rect 306984 372660 308496 372688
rect 306984 372648 306990 372660
rect 308490 372648 308496 372660
rect 308548 372648 308554 372700
rect 219894 372580 219900 372632
rect 219952 372620 219958 372632
rect 293218 372620 293224 372632
rect 219952 372592 293224 372620
rect 219952 372580 219958 372592
rect 293218 372580 293224 372592
rect 293276 372620 293282 372632
rect 342070 372620 342076 372632
rect 293276 372592 342076 372620
rect 293276 372580 293282 372592
rect 342070 372580 342076 372592
rect 342128 372580 342134 372632
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 259178 372552 259184 372564
rect 3292 372524 259184 372552
rect 3292 372512 3298 372524
rect 259178 372512 259184 372524
rect 259236 372512 259242 372564
rect 303430 372512 303436 372564
rect 303488 372552 303494 372564
rect 337378 372552 337384 372564
rect 303488 372524 337384 372552
rect 303488 372512 303494 372524
rect 337378 372512 337384 372524
rect 337436 372512 337442 372564
rect 309502 372444 309508 372496
rect 309560 372484 309566 372496
rect 309962 372484 309968 372496
rect 309560 372456 309968 372484
rect 309560 372444 309566 372456
rect 309962 372444 309968 372456
rect 310020 372444 310026 372496
rect 315206 372444 315212 372496
rect 315264 372484 315270 372496
rect 315758 372484 315764 372496
rect 315264 372456 315764 372484
rect 315264 372444 315270 372456
rect 315758 372444 315764 372456
rect 315816 372444 315822 372496
rect 323762 372444 323768 372496
rect 323820 372484 323826 372496
rect 324314 372484 324320 372496
rect 323820 372456 324320 372484
rect 323820 372444 323826 372456
rect 324314 372444 324320 372456
rect 324372 372444 324378 372496
rect 279234 372376 279240 372428
rect 279292 372416 279298 372428
rect 320818 372416 320824 372428
rect 279292 372388 320824 372416
rect 279292 372376 279298 372388
rect 320818 372376 320824 372388
rect 320876 372416 320882 372428
rect 321462 372416 321468 372428
rect 320876 372388 321468 372416
rect 320876 372376 320882 372388
rect 321462 372376 321468 372388
rect 321520 372376 321526 372428
rect 291746 372308 291752 372360
rect 291804 372348 291810 372360
rect 327718 372348 327724 372360
rect 291804 372320 327724 372348
rect 291804 372308 291810 372320
rect 327718 372308 327724 372320
rect 327776 372308 327782 372360
rect 239398 372240 239404 372292
rect 239456 372280 239462 372292
rect 295242 372280 295248 372292
rect 239456 372252 295248 372280
rect 239456 372240 239462 372252
rect 295242 372240 295248 372252
rect 295300 372240 295306 372292
rect 316034 372240 316040 372292
rect 316092 372280 316098 372292
rect 316862 372280 316868 372292
rect 316092 372252 316868 372280
rect 316092 372240 316098 372252
rect 316862 372240 316868 372252
rect 316920 372240 316926 372292
rect 238018 372172 238024 372224
rect 238076 372212 238082 372224
rect 293034 372212 293040 372224
rect 238076 372184 293040 372212
rect 238076 372172 238082 372184
rect 293034 372172 293040 372184
rect 293092 372172 293098 372224
rect 293862 372104 293868 372156
rect 293920 372144 293926 372156
rect 329650 372144 329656 372156
rect 293920 372116 329656 372144
rect 293920 372104 293926 372116
rect 329650 372104 329656 372116
rect 329708 372104 329714 372156
rect 288250 372036 288256 372088
rect 288308 372076 288314 372088
rect 328362 372076 328368 372088
rect 288308 372048 328368 372076
rect 288308 372036 288314 372048
rect 328362 372036 328368 372048
rect 328420 372036 328426 372088
rect 332686 372036 332692 372088
rect 332744 372076 332750 372088
rect 333422 372076 333428 372088
rect 332744 372048 333428 372076
rect 332744 372036 332750 372048
rect 333422 372036 333428 372048
rect 333480 372036 333486 372088
rect 281994 371968 282000 372020
rect 282052 372008 282058 372020
rect 306926 372008 306932 372020
rect 282052 371980 306932 372008
rect 282052 371968 282058 371980
rect 306926 371968 306932 371980
rect 306984 371968 306990 372020
rect 331214 371968 331220 372020
rect 331272 372008 331278 372020
rect 347498 372008 347504 372020
rect 331272 371980 347504 372008
rect 331272 371968 331278 371980
rect 347498 371968 347504 371980
rect 347556 371968 347562 372020
rect 280614 371900 280620 371952
rect 280672 371940 280678 371952
rect 285214 371940 285220 371952
rect 280672 371912 285220 371940
rect 280672 371900 280678 371912
rect 285214 371900 285220 371912
rect 285272 371900 285278 371952
rect 304718 371900 304724 371952
rect 304776 371940 304782 371952
rect 332226 371940 332232 371952
rect 304776 371912 332232 371940
rect 304776 371900 304782 371912
rect 332226 371900 332232 371912
rect 332284 371900 332290 371952
rect 332594 371900 332600 371952
rect 332652 371940 332658 371952
rect 345566 371940 345572 371952
rect 332652 371912 345572 371940
rect 332652 371900 332658 371912
rect 345566 371900 345572 371912
rect 345624 371900 345630 371952
rect 275278 371832 275284 371884
rect 275336 371872 275342 371884
rect 290458 371872 290464 371884
rect 275336 371844 290464 371872
rect 275336 371832 275342 371844
rect 290458 371832 290464 371844
rect 290516 371832 290522 371884
rect 295242 371832 295248 371884
rect 295300 371872 295306 371884
rect 336458 371872 336464 371884
rect 295300 371844 336464 371872
rect 295300 371832 295306 371844
rect 336458 371832 336464 371844
rect 336516 371832 336522 371884
rect 282270 371764 282276 371816
rect 282328 371804 282334 371816
rect 282454 371804 282460 371816
rect 282328 371776 282460 371804
rect 282328 371764 282334 371776
rect 282454 371764 282460 371776
rect 282512 371804 282518 371816
rect 308306 371804 308312 371816
rect 282512 371776 308312 371804
rect 282512 371764 282518 371776
rect 308306 371764 308312 371776
rect 308364 371764 308370 371816
rect 280614 371696 280620 371748
rect 280672 371736 280678 371748
rect 302878 371736 302884 371748
rect 280672 371708 302884 371736
rect 280672 371696 280678 371708
rect 302878 371696 302884 371708
rect 302936 371696 302942 371748
rect 280522 371628 280528 371680
rect 280580 371668 280586 371680
rect 315758 371668 315764 371680
rect 280580 371640 315764 371668
rect 280580 371628 280586 371640
rect 315758 371628 315764 371640
rect 315816 371628 315822 371680
rect 280890 371560 280896 371612
rect 280948 371600 280954 371612
rect 316034 371600 316040 371612
rect 280948 371572 316040 371600
rect 280948 371560 280954 371572
rect 316034 371560 316040 371572
rect 316092 371560 316098 371612
rect 273806 371492 273812 371544
rect 273864 371532 273870 371544
rect 309502 371532 309508 371544
rect 273864 371504 309508 371532
rect 273864 371492 273870 371504
rect 309502 371492 309508 371504
rect 309560 371492 309566 371544
rect 276566 371424 276572 371476
rect 276624 371464 276630 371476
rect 276624 371436 277394 371464
rect 276624 371424 276630 371436
rect 277366 371396 277394 371436
rect 302878 371424 302884 371476
rect 302936 371464 302942 371476
rect 314010 371464 314016 371476
rect 302936 371436 314016 371464
rect 302936 371424 302942 371436
rect 314010 371424 314016 371436
rect 314068 371424 314074 371476
rect 293862 371396 293868 371408
rect 277366 371368 293868 371396
rect 293862 371356 293868 371368
rect 293920 371356 293926 371408
rect 303522 371356 303528 371408
rect 303580 371396 303586 371408
rect 303982 371396 303988 371408
rect 303580 371368 303988 371396
rect 303580 371356 303586 371368
rect 303982 371356 303988 371368
rect 304040 371356 304046 371408
rect 320266 371356 320272 371408
rect 320324 371396 320330 371408
rect 332686 371396 332692 371408
rect 320324 371368 332692 371396
rect 320324 371356 320330 371368
rect 332686 371356 332692 371368
rect 332744 371356 332750 371408
rect 325418 371288 325424 371340
rect 325476 371328 325482 371340
rect 332594 371328 332600 371340
rect 325476 371300 332600 371328
rect 325476 371288 325482 371300
rect 332594 371288 332600 371300
rect 332652 371328 332658 371340
rect 332962 371328 332968 371340
rect 332652 371300 332968 371328
rect 332652 371288 332658 371300
rect 332962 371288 332968 371300
rect 333020 371288 333026 371340
rect 259178 371220 259184 371272
rect 259236 371260 259242 371272
rect 259730 371260 259736 371272
rect 259236 371232 259736 371260
rect 259236 371220 259242 371232
rect 259730 371220 259736 371232
rect 259788 371220 259794 371272
rect 287790 371220 287796 371272
rect 287848 371260 287854 371272
rect 290734 371260 290740 371272
rect 287848 371232 290740 371260
rect 287848 371220 287854 371232
rect 290734 371220 290740 371232
rect 290792 371220 290798 371272
rect 291838 371260 291844 371272
rect 291120 371232 291844 371260
rect 281350 371152 281356 371204
rect 281408 371192 281414 371204
rect 291120 371192 291148 371232
rect 291838 371220 291844 371232
rect 291896 371220 291902 371272
rect 323578 371220 323584 371272
rect 323636 371260 323642 371272
rect 331214 371260 331220 371272
rect 323636 371232 331220 371260
rect 323636 371220 323642 371232
rect 331214 371220 331220 371232
rect 331272 371260 331278 371272
rect 331674 371260 331680 371272
rect 331272 371232 331680 371260
rect 331272 371220 331278 371232
rect 331674 371220 331680 371232
rect 331732 371220 331738 371272
rect 281408 371164 291148 371192
rect 281408 371152 281414 371164
rect 299198 371152 299204 371204
rect 299256 371192 299262 371204
rect 332042 371192 332048 371204
rect 299256 371164 332048 371192
rect 299256 371152 299262 371164
rect 332042 371152 332048 371164
rect 332100 371152 332106 371204
rect 318886 371084 318892 371136
rect 318944 371124 318950 371136
rect 319162 371124 319168 371136
rect 318944 371096 319168 371124
rect 318944 371084 318950 371096
rect 319162 371084 319168 371096
rect 319220 371084 319226 371136
rect 279878 370948 279884 371000
rect 279936 370988 279942 371000
rect 307754 370988 307760 371000
rect 279936 370960 307760 370988
rect 279936 370948 279942 370960
rect 307754 370948 307760 370960
rect 307812 370948 307818 371000
rect 301406 370880 301412 370932
rect 301464 370920 301470 370932
rect 333330 370920 333336 370932
rect 301464 370892 333336 370920
rect 301464 370880 301470 370892
rect 333330 370880 333336 370892
rect 333388 370880 333394 370932
rect 234614 370812 234620 370864
rect 234672 370852 234678 370864
rect 234672 370824 282914 370852
rect 234672 370812 234678 370824
rect 233142 370676 233148 370728
rect 233200 370716 233206 370728
rect 281350 370716 281356 370728
rect 233200 370688 281356 370716
rect 233200 370676 233206 370688
rect 281350 370676 281356 370688
rect 281408 370676 281414 370728
rect 231762 370608 231768 370660
rect 231820 370648 231826 370660
rect 280062 370648 280068 370660
rect 231820 370620 280068 370648
rect 231820 370608 231826 370620
rect 280062 370608 280068 370620
rect 280120 370608 280126 370660
rect 282886 370648 282914 370824
rect 303430 370812 303436 370864
rect 303488 370852 303494 370864
rect 335170 370852 335176 370864
rect 303488 370824 335176 370852
rect 303488 370812 303494 370824
rect 335170 370812 335176 370824
rect 335228 370812 335234 370864
rect 296346 370744 296352 370796
rect 296404 370784 296410 370796
rect 332134 370784 332140 370796
rect 296404 370756 332140 370784
rect 296404 370744 296410 370756
rect 332134 370744 332140 370756
rect 332192 370744 332198 370796
rect 298830 370676 298836 370728
rect 298888 370716 298894 370728
rect 335262 370716 335268 370728
rect 298888 370688 335268 370716
rect 298888 370676 298894 370688
rect 335262 370676 335268 370688
rect 335320 370676 335326 370728
rect 295978 370648 295984 370660
rect 282886 370620 295984 370648
rect 295978 370608 295984 370620
rect 296036 370648 296042 370660
rect 334618 370648 334624 370660
rect 296036 370620 334624 370648
rect 296036 370608 296042 370620
rect 334618 370608 334624 370620
rect 334676 370608 334682 370660
rect 339402 370608 339408 370660
rect 339460 370648 339466 370660
rect 523678 370648 523684 370660
rect 339460 370620 523684 370648
rect 339460 370608 339466 370620
rect 523678 370608 523684 370620
rect 523736 370608 523742 370660
rect 258902 370540 258908 370592
rect 258960 370580 258966 370592
rect 318058 370580 318064 370592
rect 258960 370552 318064 370580
rect 258960 370540 258966 370552
rect 318058 370540 318064 370552
rect 318116 370580 318122 370592
rect 318702 370580 318708 370592
rect 318116 370552 318708 370580
rect 318116 370540 318122 370552
rect 318702 370540 318708 370552
rect 318760 370540 318766 370592
rect 342070 370540 342076 370592
rect 342128 370580 342134 370592
rect 580718 370580 580724 370592
rect 342128 370552 580724 370580
rect 342128 370540 342134 370552
rect 580718 370540 580724 370552
rect 580776 370540 580782 370592
rect 228358 370472 228364 370524
rect 228416 370512 228422 370524
rect 278314 370512 278320 370524
rect 228416 370484 278320 370512
rect 228416 370472 228422 370484
rect 278314 370472 278320 370484
rect 278372 370472 278378 370524
rect 290458 370472 290464 370524
rect 290516 370512 290522 370524
rect 294598 370512 294604 370524
rect 290516 370484 294604 370512
rect 290516 370472 290522 370484
rect 294598 370472 294604 370484
rect 294656 370512 294662 370524
rect 580350 370512 580356 370524
rect 294656 370484 580356 370512
rect 294656 370472 294662 370484
rect 580350 370472 580356 370484
rect 580408 370472 580414 370524
rect 271322 370404 271328 370456
rect 271380 370444 271386 370456
rect 301406 370444 301412 370456
rect 271380 370416 301412 370444
rect 271380 370404 271386 370416
rect 301406 370404 301412 370416
rect 301464 370404 301470 370456
rect 282270 370336 282276 370388
rect 282328 370376 282334 370388
rect 312078 370376 312084 370388
rect 282328 370348 312084 370376
rect 282328 370336 282334 370348
rect 312078 370336 312084 370348
rect 312136 370336 312142 370388
rect 265986 370268 265992 370320
rect 266044 370308 266050 370320
rect 298830 370308 298836 370320
rect 266044 370280 298836 370308
rect 266044 370268 266050 370280
rect 298830 370268 298836 370280
rect 298888 370268 298894 370320
rect 281442 370200 281448 370252
rect 281500 370240 281506 370252
rect 314194 370240 314200 370252
rect 281500 370212 314200 370240
rect 281500 370200 281506 370212
rect 314194 370200 314200 370212
rect 314252 370200 314258 370252
rect 235350 370132 235356 370184
rect 235408 370172 235414 370184
rect 296346 370172 296352 370184
rect 235408 370144 296352 370172
rect 235408 370132 235414 370144
rect 296346 370132 296352 370144
rect 296404 370132 296410 370184
rect 242158 370064 242164 370116
rect 242216 370104 242222 370116
rect 302372 370104 302378 370116
rect 242216 370076 302378 370104
rect 242216 370064 242222 370076
rect 302372 370064 302378 370076
rect 302430 370104 302436 370116
rect 303430 370104 303436 370116
rect 302430 370076 303436 370104
rect 302430 370064 302436 370076
rect 303430 370064 303436 370076
rect 303488 370064 303494 370116
rect 306420 370064 306426 370116
rect 306478 370104 306484 370116
rect 307018 370104 307024 370116
rect 306478 370076 307024 370104
rect 306478 370064 306484 370076
rect 307018 370064 307024 370076
rect 307076 370064 307082 370116
rect 312078 370064 312084 370116
rect 312136 370104 312142 370116
rect 312676 370104 312682 370116
rect 312136 370076 312682 370104
rect 312136 370064 312142 370076
rect 312676 370064 312682 370076
rect 312734 370064 312740 370116
rect 314194 370064 314200 370116
rect 314252 370104 314258 370116
rect 314516 370104 314522 370116
rect 314252 370076 314522 370104
rect 314252 370064 314258 370076
rect 314516 370064 314522 370076
rect 314574 370064 314580 370116
rect 318978 370064 318984 370116
rect 319036 370104 319042 370116
rect 320036 370104 320042 370116
rect 319036 370076 320042 370104
rect 319036 370064 319042 370076
rect 320036 370064 320042 370076
rect 320094 370064 320100 370116
rect 322290 370064 322296 370116
rect 322348 370104 322354 370116
rect 323348 370104 323354 370116
rect 322348 370076 323354 370104
rect 322348 370064 322354 370076
rect 323348 370064 323354 370076
rect 323406 370064 323412 370116
rect 280798 369996 280804 370048
rect 280856 370036 280862 370048
rect 317690 370036 317696 370048
rect 280856 370008 317696 370036
rect 280856 369996 280862 370008
rect 317690 369996 317696 370008
rect 317748 369996 317754 370048
rect 279326 369928 279332 369980
rect 279384 369968 279390 369980
rect 279878 369968 279884 369980
rect 279384 369940 279884 369968
rect 279384 369928 279390 369940
rect 279878 369928 279884 369940
rect 279936 369928 279942 369980
rect 293034 369928 293040 369980
rect 293092 369968 293098 369980
rect 339402 369968 339408 369980
rect 293092 369940 339408 369968
rect 293092 369928 293098 369940
rect 339402 369928 339408 369940
rect 339460 369928 339466 369980
rect 245010 369860 245016 369912
rect 245068 369900 245074 369912
rect 304350 369900 304356 369912
rect 245068 369872 304356 369900
rect 245068 369860 245074 369872
rect 304350 369860 304356 369872
rect 304408 369860 304414 369912
rect 340874 369832 340880 369844
rect 291580 369804 340880 369832
rect 291580 369776 291608 369804
rect 340874 369792 340880 369804
rect 340932 369792 340938 369844
rect 291562 369724 291568 369776
rect 291620 369724 291626 369776
rect 292546 369532 311894 369560
rect 291102 369424 291108 369436
rect 282886 369396 291108 369424
rect 233878 369180 233884 369232
rect 233936 369220 233942 369232
rect 279142 369220 279148 369232
rect 233936 369192 279148 369220
rect 233936 369180 233942 369192
rect 279142 369180 279148 369192
rect 279200 369180 279206 369232
rect 231118 369112 231124 369164
rect 231176 369152 231182 369164
rect 282886 369152 282914 369396
rect 291102 369384 291108 369396
rect 291160 369384 291166 369436
rect 292298 369384 292304 369436
rect 292356 369424 292362 369436
rect 292546 369424 292574 369532
rect 305086 369492 305092 369504
rect 292356 369396 292574 369424
rect 297376 369464 305092 369492
rect 292356 369384 292362 369396
rect 231176 369124 282914 369152
rect 231176 369112 231182 369124
rect 245654 368636 245660 368688
rect 245712 368676 245718 368688
rect 297376 368676 297404 369464
rect 305086 369452 305092 369464
rect 305144 369492 305150 369504
rect 305454 369492 305460 369504
rect 305144 369464 305460 369492
rect 305144 369452 305150 369464
rect 305454 369452 305460 369464
rect 305512 369452 305518 369504
rect 303982 369424 303988 369436
rect 245712 368648 297404 368676
rect 299446 369396 303988 369424
rect 245712 368636 245718 368648
rect 243262 368568 243268 368620
rect 243320 368608 243326 368620
rect 299446 368608 299474 369396
rect 303982 369384 303988 369396
rect 304040 369384 304046 369436
rect 243320 368580 299474 368608
rect 243320 368568 243326 368580
rect 228450 368500 228456 368552
rect 228508 368540 228514 368552
rect 276014 368540 276020 368552
rect 228508 368512 276020 368540
rect 228508 368500 228514 368512
rect 276014 368500 276020 368512
rect 276072 368500 276078 368552
rect 311866 368540 311894 369532
rect 340874 369112 340880 369164
rect 340932 369152 340938 369164
rect 341978 369152 341984 369164
rect 340932 369124 341984 369152
rect 340932 369112 340938 369124
rect 341978 369112 341984 369124
rect 342036 369152 342042 369164
rect 580626 369152 580632 369164
rect 342036 369124 580632 369152
rect 342036 369112 342042 369124
rect 580626 369112 580632 369124
rect 580684 369112 580690 369164
rect 333882 368976 333888 369028
rect 333940 369016 333946 369028
rect 334618 369016 334624 369028
rect 333940 368988 334624 369016
rect 333940 368976 333946 368988
rect 334618 368976 334624 368988
rect 334676 368976 334682 369028
rect 388438 368540 388444 368552
rect 311866 368512 388444 368540
rect 388438 368500 388444 368512
rect 388496 368500 388502 368552
rect 329742 367752 329748 367804
rect 329800 367792 329806 367804
rect 384298 367792 384304 367804
rect 329800 367764 384304 367792
rect 329800 367752 329806 367764
rect 384298 367752 384304 367764
rect 384356 367752 384362 367804
rect 329650 365644 329656 365696
rect 329708 365684 329714 365696
rect 342162 365684 342168 365696
rect 329708 365656 342168 365684
rect 329708 365644 329714 365656
rect 342162 365644 342168 365656
rect 342220 365684 342226 365696
rect 580166 365684 580172 365696
rect 342220 365656 580172 365684
rect 342220 365644 342226 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 249058 363604 249064 363656
rect 249116 363644 249122 363656
rect 274542 363644 274548 363656
rect 249116 363616 274548 363644
rect 249116 363604 249122 363616
rect 274542 363604 274548 363616
rect 274600 363604 274606 363656
rect 329098 363604 329104 363656
rect 329156 363644 329162 363656
rect 382642 363644 382648 363656
rect 329156 363616 382648 363644
rect 329156 363604 329162 363616
rect 382642 363604 382648 363616
rect 382700 363604 382706 363656
rect 256050 362176 256056 362228
rect 256108 362216 256114 362228
rect 280522 362216 280528 362228
rect 256108 362188 280528 362216
rect 256108 362176 256114 362188
rect 280522 362176 280528 362188
rect 280580 362176 280586 362228
rect 224218 361564 224224 361616
rect 224276 361604 224282 361616
rect 279878 361604 279884 361616
rect 224276 361576 279884 361604
rect 224276 361564 224282 361576
rect 279878 361564 279884 361576
rect 279936 361604 279942 361616
rect 280062 361604 280068 361616
rect 279936 361576 280068 361604
rect 279936 361564 279942 361576
rect 280062 361564 280068 361576
rect 280120 361564 280126 361616
rect 253290 359456 253296 359508
rect 253348 359496 253354 359508
rect 280614 359496 280620 359508
rect 253348 359468 280620 359496
rect 253348 359456 253354 359468
rect 280614 359456 280620 359468
rect 280672 359456 280678 359508
rect 331122 359456 331128 359508
rect 331180 359496 331186 359508
rect 375834 359496 375840 359508
rect 331180 359468 375840 359496
rect 331180 359456 331186 359468
rect 375834 359456 375840 359468
rect 375892 359456 375898 359508
rect 268562 358028 268568 358080
rect 268620 358068 268626 358080
rect 279418 358068 279424 358080
rect 268620 358040 279424 358068
rect 268620 358028 268626 358040
rect 279418 358028 279424 358040
rect 279476 358028 279482 358080
rect 333330 358028 333336 358080
rect 333388 358068 333394 358080
rect 352190 358068 352196 358080
rect 333388 358040 352196 358068
rect 333388 358028 333394 358040
rect 352190 358028 352196 358040
rect 352248 358028 352254 358080
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 268562 357456 268568 357468
rect 3200 357428 268568 357456
rect 3200 357416 3206 357428
rect 268562 357416 268568 357428
rect 268620 357416 268626 357468
rect 335170 356668 335176 356720
rect 335228 356708 335234 356720
rect 345382 356708 345388 356720
rect 335228 356680 345388 356708
rect 335228 356668 335234 356680
rect 345382 356668 345388 356680
rect 345440 356668 345446 356720
rect 333422 355308 333428 355360
rect 333480 355348 333486 355360
rect 350626 355348 350632 355360
rect 333480 355320 350632 355348
rect 333480 355308 333486 355320
rect 350626 355308 350632 355320
rect 350684 355308 350690 355360
rect 229830 353948 229836 354000
rect 229888 353988 229894 354000
rect 276014 353988 276020 354000
rect 229888 353960 276020 353988
rect 229888 353948 229894 353960
rect 276014 353948 276020 353960
rect 276072 353948 276078 354000
rect 330386 353948 330392 354000
rect 330444 353988 330450 354000
rect 375742 353988 375748 354000
rect 330444 353960 375748 353988
rect 330444 353948 330450 353960
rect 375742 353948 375748 353960
rect 375800 353948 375806 354000
rect 276014 353268 276020 353320
rect 276072 353308 276078 353320
rect 277302 353308 277308 353320
rect 276072 353280 277308 353308
rect 276072 353268 276078 353280
rect 277302 353268 277308 353280
rect 277360 353308 277366 353320
rect 278038 353308 278044 353320
rect 277360 353280 278044 353308
rect 277360 353268 277366 353280
rect 278038 353268 278044 353280
rect 278096 353268 278102 353320
rect 257430 351160 257436 351212
rect 257488 351200 257494 351212
rect 280890 351200 280896 351212
rect 257488 351172 280896 351200
rect 257488 351160 257494 351172
rect 280890 351160 280896 351172
rect 280948 351160 280954 351212
rect 261754 349800 261760 349852
rect 261812 349840 261818 349852
rect 279234 349840 279240 349852
rect 261812 349812 279240 349840
rect 261812 349800 261818 349812
rect 279234 349800 279240 349812
rect 279292 349800 279298 349852
rect 332042 349800 332048 349852
rect 332100 349840 332106 349852
rect 351638 349840 351644 349852
rect 332100 349812 351644 349840
rect 332100 349800 332106 349812
rect 351638 349800 351644 349812
rect 351696 349800 351702 349852
rect 332134 348372 332140 348424
rect 332192 348412 332198 348424
rect 349246 348412 349252 348424
rect 332192 348384 349252 348412
rect 332192 348372 332198 348384
rect 349246 348372 349252 348384
rect 349304 348372 349310 348424
rect 256694 345652 256700 345704
rect 256752 345692 256758 345704
rect 280798 345692 280804 345704
rect 256752 345664 280804 345692
rect 256752 345652 256758 345664
rect 280798 345652 280804 345664
rect 280856 345652 280862 345704
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 256694 345080 256700 345092
rect 3384 345052 256700 345080
rect 3384 345040 3390 345052
rect 256694 345040 256700 345052
rect 256752 345040 256758 345092
rect 332226 342864 332232 342916
rect 332284 342904 332290 342916
rect 349614 342904 349620 342916
rect 332284 342876 349620 342904
rect 332284 342864 332290 342876
rect 349614 342864 349620 342876
rect 349672 342864 349678 342916
rect 329558 334568 329564 334620
rect 329616 334608 329622 334620
rect 385678 334608 385684 334620
rect 329616 334580 385684 334608
rect 329616 334568 329622 334580
rect 385678 334568 385684 334580
rect 385736 334568 385742 334620
rect 380158 333956 380164 334008
rect 380216 333996 380222 334008
rect 380802 333996 380808 334008
rect 380216 333968 380808 333996
rect 380216 333956 380222 333968
rect 380802 333956 380808 333968
rect 380860 333996 380866 334008
rect 498194 333996 498200 334008
rect 380860 333968 498200 333996
rect 380860 333956 380866 333968
rect 498194 333956 498200 333968
rect 498252 333956 498258 334008
rect 333698 333208 333704 333260
rect 333756 333248 333762 333260
rect 389634 333248 389640 333260
rect 333756 333220 389640 333248
rect 333756 333208 333762 333220
rect 389634 333208 389640 333220
rect 389692 333208 389698 333260
rect 379882 332596 379888 332648
rect 379940 332636 379946 332648
rect 484394 332636 484400 332648
rect 379940 332608 484400 332636
rect 379940 332596 379946 332608
rect 484394 332596 484400 332608
rect 484452 332596 484458 332648
rect 335906 331848 335912 331900
rect 335964 331888 335970 331900
rect 379882 331888 379888 331900
rect 335964 331860 379888 331888
rect 335964 331848 335970 331860
rect 379882 331848 379888 331860
rect 379940 331848 379946 331900
rect 385310 330488 385316 330540
rect 385368 330528 385374 330540
rect 385770 330528 385776 330540
rect 385368 330500 385776 330528
rect 385368 330488 385374 330500
rect 385770 330488 385776 330500
rect 385828 330488 385834 330540
rect 386966 329808 386972 329860
rect 387024 329848 387030 329860
rect 569954 329848 569960 329860
rect 387024 329820 569960 329848
rect 387024 329808 387030 329820
rect 569954 329808 569960 329820
rect 570012 329808 570018 329860
rect 329006 329060 329012 329112
rect 329064 329100 329070 329112
rect 384206 329100 384212 329112
rect 329064 329072 384212 329100
rect 329064 329060 329070 329072
rect 384206 329060 384212 329072
rect 384264 329060 384270 329112
rect 385310 327020 385316 327072
rect 385368 327060 385374 327072
rect 385586 327060 385592 327072
rect 385368 327032 385592 327060
rect 385368 327020 385374 327032
rect 385586 327020 385592 327032
rect 385644 327020 385650 327072
rect 280982 326544 280988 326596
rect 281040 326544 281046 326596
rect 281000 326392 281028 326544
rect 337286 326408 337292 326460
rect 337344 326448 337350 326460
rect 378594 326448 378600 326460
rect 337344 326420 378600 326448
rect 337344 326408 337350 326420
rect 378594 326408 378600 326420
rect 378652 326408 378658 326460
rect 233970 326340 233976 326392
rect 234028 326380 234034 326392
rect 276566 326380 276572 326392
rect 234028 326352 276572 326380
rect 234028 326340 234034 326352
rect 276566 326340 276572 326352
rect 276624 326340 276630 326392
rect 280982 326340 280988 326392
rect 281040 326340 281046 326392
rect 329650 326340 329656 326392
rect 329708 326380 329714 326392
rect 372982 326380 372988 326392
rect 329708 326352 372988 326380
rect 329708 326340 329714 326352
rect 372982 326340 372988 326352
rect 373040 326340 373046 326392
rect 385310 325728 385316 325780
rect 385368 325768 385374 325780
rect 547874 325768 547880 325780
rect 385368 325740 547880 325768
rect 385368 325728 385374 325740
rect 547874 325728 547880 325740
rect 547932 325728 547938 325780
rect 385678 325660 385684 325712
rect 385736 325700 385742 325712
rect 563054 325700 563060 325712
rect 385736 325672 563060 325700
rect 385736 325660 385742 325672
rect 563054 325660 563060 325672
rect 563112 325660 563118 325712
rect 388438 325592 388444 325644
rect 388496 325632 388502 325644
rect 579982 325632 579988 325644
rect 388496 325604 579988 325632
rect 388496 325592 388502 325604
rect 579982 325592 579988 325604
rect 580040 325592 580046 325644
rect 333974 325048 333980 325100
rect 334032 325088 334038 325100
rect 378502 325088 378508 325100
rect 334032 325060 378508 325088
rect 334032 325048 334038 325060
rect 378502 325048 378508 325060
rect 378560 325048 378566 325100
rect 337194 324980 337200 325032
rect 337252 325020 337258 325032
rect 377214 325020 377220 325032
rect 337252 324992 377220 325020
rect 337252 324980 337258 324992
rect 377214 324980 377220 324992
rect 377272 324980 377278 325032
rect 231210 324912 231216 324964
rect 231268 324952 231274 324964
rect 275278 324952 275284 324964
rect 231268 324924 275284 324952
rect 231268 324912 231274 324924
rect 275278 324912 275284 324924
rect 275336 324912 275342 324964
rect 372614 324912 372620 324964
rect 372672 324952 372678 324964
rect 384482 324952 384488 324964
rect 372672 324924 384488 324952
rect 372672 324912 372678 324924
rect 384482 324912 384488 324924
rect 384540 324952 384546 324964
rect 396074 324952 396080 324964
rect 384540 324924 396080 324952
rect 384540 324912 384546 324924
rect 396074 324912 396080 324924
rect 396132 324912 396138 324964
rect 340782 323688 340788 323740
rect 340840 323728 340846 323740
rect 372614 323728 372620 323740
rect 340840 323700 372620 323728
rect 340840 323688 340846 323700
rect 372614 323688 372620 323700
rect 372672 323688 372678 323740
rect 342254 323620 342260 323672
rect 342312 323660 342318 323672
rect 385402 323660 385408 323672
rect 342312 323632 385408 323660
rect 342312 323620 342318 323632
rect 385402 323620 385408 323632
rect 385460 323620 385466 323672
rect 331214 323552 331220 323604
rect 331272 323592 331278 323604
rect 331766 323592 331772 323604
rect 331272 323564 331772 323592
rect 331272 323552 331278 323564
rect 331766 323552 331772 323564
rect 331824 323592 331830 323604
rect 384114 323592 384120 323604
rect 331824 323564 384120 323592
rect 331824 323552 331830 323564
rect 384114 323552 384120 323564
rect 384172 323552 384178 323604
rect 263318 322940 263324 322992
rect 263376 322980 263382 322992
rect 280982 322980 280988 322992
rect 263376 322952 280988 322980
rect 263376 322940 263382 322952
rect 280982 322940 280988 322952
rect 281040 322940 281046 322992
rect 330386 322872 330392 322924
rect 330444 322912 330450 322924
rect 384022 322912 384028 322924
rect 330444 322884 384028 322912
rect 330444 322872 330450 322884
rect 384022 322872 384028 322884
rect 384080 322872 384086 322924
rect 331306 322804 331312 322856
rect 331364 322844 331370 322856
rect 338022 322844 338028 322856
rect 331364 322816 338028 322844
rect 331364 322804 331370 322816
rect 338022 322804 338028 322816
rect 338080 322804 338086 322856
rect 209682 322260 209688 322312
rect 209740 322300 209746 322312
rect 260466 322300 260472 322312
rect 209740 322272 260472 322300
rect 209740 322260 209746 322272
rect 260466 322260 260472 322272
rect 260524 322260 260530 322312
rect 385770 322300 385776 322312
rect 373966 322272 385776 322300
rect 212442 322192 212448 322244
rect 212500 322232 212506 322244
rect 263318 322232 263324 322244
rect 212500 322204 263324 322232
rect 212500 322192 212506 322204
rect 263318 322192 263324 322204
rect 263376 322192 263382 322244
rect 332686 322192 332692 322244
rect 332744 322232 332750 322244
rect 373966 322232 373994 322272
rect 385770 322260 385776 322272
rect 385828 322260 385834 322312
rect 332744 322204 373994 322232
rect 332744 322192 332750 322204
rect 327442 321852 327448 321904
rect 327500 321892 327506 321904
rect 327626 321892 327632 321904
rect 327500 321864 327632 321892
rect 327500 321852 327506 321864
rect 327626 321852 327632 321864
rect 327684 321852 327690 321904
rect 216582 321648 216588 321700
rect 216640 321688 216646 321700
rect 265802 321688 265808 321700
rect 216640 321660 265808 321688
rect 216640 321648 216646 321660
rect 265802 321648 265808 321660
rect 265860 321648 265866 321700
rect 204070 321580 204076 321632
rect 204128 321620 204134 321632
rect 273898 321620 273904 321632
rect 204128 321592 273904 321620
rect 204128 321580 204134 321592
rect 273898 321580 273904 321592
rect 273956 321580 273962 321632
rect 378042 321580 378048 321632
rect 378100 321620 378106 321632
rect 378410 321620 378416 321632
rect 378100 321592 378416 321620
rect 378100 321580 378106 321592
rect 378410 321580 378416 321592
rect 378468 321580 378474 321632
rect 327810 321512 327816 321564
rect 327868 321552 327874 321564
rect 328086 321552 328092 321564
rect 327868 321524 328092 321552
rect 327868 321512 327874 321524
rect 328086 321512 328092 321524
rect 328144 321512 328150 321564
rect 275278 321376 275284 321428
rect 275336 321416 275342 321428
rect 279510 321416 279516 321428
rect 275336 321388 279516 321416
rect 275336 321376 275342 321388
rect 279510 321376 279516 321388
rect 279568 321416 279574 321428
rect 281994 321416 282000 321428
rect 279568 321388 282000 321416
rect 279568 321376 279574 321388
rect 281994 321376 282000 321388
rect 282052 321376 282058 321428
rect 291166 321388 306374 321416
rect 249150 321104 249156 321156
rect 249208 321144 249214 321156
rect 273806 321144 273812 321156
rect 249208 321116 273812 321144
rect 249208 321104 249214 321116
rect 273806 321104 273812 321116
rect 273864 321104 273870 321156
rect 287532 321116 287928 321144
rect 268654 321076 268660 321088
rect 258046 321048 268660 321076
rect 208302 320900 208308 320952
rect 208360 320940 208366 320952
rect 258046 320940 258074 321048
rect 268654 321036 268660 321048
rect 268712 321076 268718 321088
rect 287532 321076 287560 321116
rect 268712 321048 287560 321076
rect 287900 321076 287928 321116
rect 287900 321048 290044 321076
rect 268712 321036 268718 321048
rect 277854 320968 277860 321020
rect 277912 320968 277918 321020
rect 208360 320912 258074 320940
rect 208360 320900 208366 320912
rect 209498 320832 209504 320884
rect 209556 320872 209562 320884
rect 277872 320872 277900 320968
rect 280890 320872 280896 320884
rect 209556 320844 280896 320872
rect 209556 320832 209562 320844
rect 280890 320832 280896 320844
rect 280948 320832 280954 320884
rect 282086 320696 282092 320748
rect 282144 320736 282150 320748
rect 285904 320736 285910 320748
rect 282144 320708 285910 320736
rect 282144 320696 282150 320708
rect 285904 320696 285910 320708
rect 285962 320696 285968 320748
rect 290016 320736 290044 321048
rect 290228 320736 290234 320748
rect 290016 320708 290234 320736
rect 290228 320696 290234 320708
rect 290286 320696 290292 320748
rect 274358 320628 274364 320680
rect 274416 320668 274422 320680
rect 280614 320668 280620 320680
rect 274416 320640 280620 320668
rect 274416 320628 274422 320640
rect 280614 320628 280620 320640
rect 280672 320628 280678 320680
rect 280706 320532 280712 320544
rect 278746 320504 280712 320532
rect 273530 320356 273536 320408
rect 273588 320396 273594 320408
rect 278746 320396 278774 320504
rect 280706 320492 280712 320504
rect 280764 320532 280770 320544
rect 281350 320532 281356 320544
rect 280764 320504 281356 320532
rect 280764 320492 280770 320504
rect 281350 320492 281356 320504
rect 281408 320492 281414 320544
rect 273588 320368 278774 320396
rect 273588 320356 273594 320368
rect 271046 320288 271052 320340
rect 271104 320328 271110 320340
rect 282178 320328 282184 320340
rect 271104 320300 282184 320328
rect 271104 320288 271110 320300
rect 282178 320288 282184 320300
rect 282236 320288 282242 320340
rect 216398 320152 216404 320204
rect 216456 320192 216462 320204
rect 216456 320164 291102 320192
rect 216456 320152 216462 320164
rect 272426 320084 272432 320136
rect 272484 320124 272490 320136
rect 272610 320124 272616 320136
rect 272484 320096 272616 320124
rect 272484 320084 272490 320096
rect 272610 320084 272616 320096
rect 272668 320084 272674 320136
rect 282178 320084 282184 320136
rect 282236 320124 282242 320136
rect 282236 320096 291010 320124
rect 282236 320084 282242 320096
rect 281994 320016 282000 320068
rect 282052 320056 282058 320068
rect 282052 320028 286134 320056
rect 282052 320016 282058 320028
rect 281902 319948 281908 320000
rect 281960 319988 281966 320000
rect 281960 319960 284800 319988
rect 281960 319948 281966 319960
rect 273990 319880 273996 319932
rect 274048 319920 274054 319932
rect 284772 319920 284800 319960
rect 286106 319932 286134 320028
rect 290384 319960 290918 319988
rect 284846 319920 284852 319932
rect 274048 319892 284708 319920
rect 284772 319892 284852 319920
rect 274048 319880 274054 319892
rect 216490 319812 216496 319864
rect 216548 319852 216554 319864
rect 276934 319852 276940 319864
rect 216548 319824 276940 319852
rect 216548 319812 216554 319824
rect 276934 319812 276940 319824
rect 276992 319812 276998 319864
rect 282592 319812 282598 319864
rect 282650 319812 282656 319864
rect 284680 319852 284708 319892
rect 284846 319880 284852 319892
rect 284904 319880 284910 319932
rect 286088 319880 286094 319932
rect 286146 319880 286152 319932
rect 289952 319880 289958 319932
rect 290010 319920 290016 319932
rect 290010 319880 290044 319920
rect 290136 319880 290142 319932
rect 290194 319920 290200 319932
rect 290274 319920 290280 319932
rect 290194 319892 290280 319920
rect 290194 319880 290200 319892
rect 290274 319880 290280 319892
rect 290332 319880 290338 319932
rect 289262 319852 289268 319864
rect 284680 319824 289268 319852
rect 289262 319812 289268 319824
rect 289320 319812 289326 319864
rect 213086 319744 213092 319796
rect 213144 319784 213150 319796
rect 269482 319784 269488 319796
rect 213144 319756 269488 319784
rect 213144 319744 213150 319756
rect 269482 319744 269488 319756
rect 269540 319744 269546 319796
rect 281718 319784 281724 319796
rect 273226 319756 281724 319784
rect 217962 319608 217968 319660
rect 218020 319648 218026 319660
rect 273226 319648 273254 319756
rect 281718 319744 281724 319756
rect 281776 319784 281782 319796
rect 282610 319784 282638 319812
rect 281776 319756 282638 319784
rect 281776 319744 281782 319756
rect 282822 319744 282828 319796
rect 282880 319784 282886 319796
rect 284846 319784 284852 319796
rect 282880 319756 284852 319784
rect 282880 319744 282886 319756
rect 284846 319744 284852 319756
rect 284904 319744 284910 319796
rect 285600 319756 285812 319784
rect 280890 319676 280896 319728
rect 280948 319716 280954 319728
rect 285600 319716 285628 319756
rect 280948 319688 285628 319716
rect 285784 319716 285812 319756
rect 290016 319716 290044 319880
rect 290384 319852 290412 319960
rect 290890 319932 290918 319960
rect 290872 319880 290878 319932
rect 290930 319880 290936 319932
rect 290688 319852 290694 319864
rect 290200 319824 290412 319852
rect 290476 319824 290694 319852
rect 290200 319796 290228 319824
rect 290182 319744 290188 319796
rect 290240 319744 290246 319796
rect 285784 319688 290044 319716
rect 280948 319676 280954 319688
rect 218020 319620 273254 319648
rect 218020 319608 218026 319620
rect 279970 319608 279976 319660
rect 280028 319648 280034 319660
rect 280522 319648 280528 319660
rect 280028 319620 280528 319648
rect 280028 319608 280034 319620
rect 280522 319608 280528 319620
rect 280580 319648 280586 319660
rect 280580 319620 285076 319648
rect 280580 319608 280586 319620
rect 216306 319540 216312 319592
rect 216364 319580 216370 319592
rect 277118 319580 277124 319592
rect 216364 319552 277124 319580
rect 216364 319540 216370 319552
rect 277118 319540 277124 319552
rect 277176 319580 277182 319592
rect 277176 319552 284984 319580
rect 277176 319540 277182 319552
rect 213730 319472 213736 319524
rect 213788 319512 213794 319524
rect 274174 319512 274180 319524
rect 213788 319484 274180 319512
rect 213788 319472 213794 319484
rect 274174 319472 274180 319484
rect 274232 319512 274238 319524
rect 282822 319512 282828 319524
rect 274232 319484 282828 319512
rect 274232 319472 274238 319484
rect 282822 319472 282828 319484
rect 282880 319472 282886 319524
rect 283558 319512 283564 319524
rect 283484 319484 283564 319512
rect 3418 319404 3424 319456
rect 3476 319444 3482 319456
rect 258350 319444 258356 319456
rect 3476 319416 258356 319444
rect 3476 319404 3482 319416
rect 258350 319404 258356 319416
rect 258408 319444 258414 319456
rect 258902 319444 258908 319456
rect 258408 319416 258908 319444
rect 258408 319404 258414 319416
rect 258902 319404 258908 319416
rect 258960 319404 258966 319456
rect 276934 319404 276940 319456
rect 276992 319444 276998 319456
rect 281994 319444 282000 319456
rect 276992 319416 282000 319444
rect 276992 319404 276998 319416
rect 281994 319404 282000 319416
rect 282052 319404 282058 319456
rect 283282 319336 283288 319388
rect 283340 319376 283346 319388
rect 283484 319376 283512 319484
rect 283558 319472 283564 319484
rect 283616 319472 283622 319524
rect 284956 319444 284984 319552
rect 285048 319512 285076 319620
rect 286594 319540 286600 319592
rect 286652 319580 286658 319592
rect 287606 319580 287612 319592
rect 286652 319552 287612 319580
rect 286652 319540 286658 319552
rect 287606 319540 287612 319552
rect 287664 319580 287670 319592
rect 289078 319580 289084 319592
rect 287664 319552 289084 319580
rect 287664 319540 287670 319552
rect 289078 319540 289084 319552
rect 289136 319540 289142 319592
rect 290476 319580 290504 319824
rect 290688 319812 290694 319824
rect 290746 319812 290752 319864
rect 290780 319812 290786 319864
rect 290838 319812 290844 319864
rect 290982 319852 291010 320096
rect 290890 319824 291010 319852
rect 291074 319852 291102 320164
rect 291166 319932 291194 321388
rect 306346 321144 306374 321388
rect 327902 321376 327908 321428
rect 327960 321416 327966 321428
rect 328270 321416 328276 321428
rect 327960 321388 328276 321416
rect 327960 321376 327966 321388
rect 328270 321376 328276 321388
rect 328328 321376 328334 321428
rect 332686 321240 332692 321292
rect 332744 321280 332750 321292
rect 370590 321280 370596 321292
rect 332744 321252 370596 321280
rect 332744 321240 332750 321252
rect 370590 321240 370596 321252
rect 370648 321240 370654 321292
rect 327718 321172 327724 321224
rect 327776 321212 327782 321224
rect 361022 321212 361028 321224
rect 327776 321184 361028 321212
rect 327776 321172 327782 321184
rect 361022 321172 361028 321184
rect 361080 321172 361086 321224
rect 344738 321144 344744 321156
rect 306346 321116 344744 321144
rect 344738 321104 344744 321116
rect 344796 321104 344802 321156
rect 357986 321076 357992 321088
rect 298618 321048 357992 321076
rect 292086 319960 296944 319988
rect 291148 319880 291154 319932
rect 291206 319880 291212 319932
rect 292086 319852 292114 319960
rect 292160 319880 292166 319932
rect 292218 319880 292224 319932
rect 291074 319824 292114 319852
rect 290798 319784 290826 319812
rect 290752 319756 290826 319784
rect 290550 319580 290556 319592
rect 290476 319552 290556 319580
rect 290550 319540 290556 319552
rect 290608 319540 290614 319592
rect 285048 319484 287744 319512
rect 287606 319444 287612 319456
rect 284956 319416 287612 319444
rect 287606 319404 287612 319416
rect 287664 319404 287670 319456
rect 283340 319348 283512 319376
rect 283340 319336 283346 319348
rect 283558 319336 283564 319388
rect 283616 319376 283622 319388
rect 283742 319376 283748 319388
rect 283616 319348 283748 319376
rect 283616 319336 283622 319348
rect 283742 319336 283748 319348
rect 283800 319336 283806 319388
rect 287716 319376 287744 319484
rect 289998 319472 290004 319524
rect 290056 319512 290062 319524
rect 290752 319512 290780 319756
rect 290890 319648 290918 319824
rect 291838 319744 291844 319796
rect 291896 319784 291902 319796
rect 292178 319784 292206 319880
rect 294138 319784 294144 319796
rect 291896 319756 292206 319784
rect 292270 319756 294144 319784
rect 291896 319744 291902 319756
rect 292270 319716 292298 319756
rect 294138 319744 294144 319756
rect 294196 319744 294202 319796
rect 295426 319716 295432 319728
rect 291120 319688 292298 319716
rect 292454 319688 295432 319716
rect 291120 319648 291148 319688
rect 290890 319620 291148 319648
rect 291194 319608 291200 319660
rect 291252 319648 291258 319660
rect 292454 319648 292482 319688
rect 295426 319676 295432 319688
rect 295484 319676 295490 319728
rect 295656 319676 295662 319728
rect 295714 319716 295720 319728
rect 296346 319716 296352 319728
rect 295714 319688 296352 319716
rect 295714 319676 295720 319688
rect 296346 319676 296352 319688
rect 296404 319676 296410 319728
rect 291252 319620 292482 319648
rect 291252 319608 291258 319620
rect 293954 319608 293960 319660
rect 294012 319648 294018 319660
rect 295794 319648 295800 319660
rect 294012 319620 295800 319648
rect 294012 319608 294018 319620
rect 295794 319608 295800 319620
rect 295852 319608 295858 319660
rect 296916 319648 296944 319960
rect 298618 319716 298646 321048
rect 357986 321036 357992 321048
rect 358044 321036 358050 321088
rect 358170 321008 358176 321020
rect 298710 320980 358176 321008
rect 298710 319988 298738 320980
rect 358170 320968 358176 320980
rect 358228 320968 358234 321020
rect 368014 320940 368020 320952
rect 307634 320912 368020 320940
rect 307634 320612 307662 320912
rect 368014 320900 368020 320912
rect 368072 320900 368078 320952
rect 354306 320872 354312 320884
rect 307864 320844 354312 320872
rect 307616 320560 307622 320612
rect 307674 320560 307680 320612
rect 307864 320532 307892 320844
rect 354306 320832 354312 320844
rect 354364 320832 354370 320884
rect 314792 320696 314798 320748
rect 314850 320736 314856 320748
rect 327718 320736 327724 320748
rect 314850 320708 327724 320736
rect 314850 320696 314856 320708
rect 327718 320696 327724 320708
rect 327776 320696 327782 320748
rect 307726 320504 307892 320532
rect 307726 320464 307754 320504
rect 302758 320436 307754 320464
rect 302758 320124 302786 320436
rect 327810 320260 327816 320272
rect 308002 320232 309134 320260
rect 308002 320192 308030 320232
rect 302942 320164 308030 320192
rect 302758 320096 302832 320124
rect 298848 320028 302694 320056
rect 298710 319960 298784 319988
rect 298756 319864 298784 319960
rect 298738 319812 298744 319864
rect 298796 319812 298802 319864
rect 298848 319728 298876 320028
rect 299906 319960 302602 319988
rect 299906 319932 299934 319960
rect 299888 319920 299894 319932
rect 299032 319892 299894 319920
rect 299032 319796 299060 319892
rect 299888 319880 299894 319892
rect 299946 319880 299952 319932
rect 301176 319920 301182 319932
rect 301148 319880 301182 319920
rect 301234 319880 301240 319932
rect 301636 319880 301642 319932
rect 301694 319880 301700 319932
rect 302188 319880 302194 319932
rect 302246 319880 302252 319932
rect 299014 319744 299020 319796
rect 299072 319744 299078 319796
rect 298738 319716 298744 319728
rect 298618 319688 298744 319716
rect 298738 319676 298744 319688
rect 298796 319676 298802 319728
rect 298830 319676 298836 319728
rect 298888 319676 298894 319728
rect 301148 319660 301176 319880
rect 301654 319716 301682 319880
rect 302206 319728 302234 319880
rect 301332 319688 301682 319716
rect 301332 319660 301360 319688
rect 302142 319676 302148 319728
rect 302200 319688 302234 319728
rect 302574 319716 302602 319960
rect 302666 319932 302694 320028
rect 302804 319932 302832 320096
rect 302648 319880 302654 319932
rect 302706 319880 302712 319932
rect 302786 319880 302792 319932
rect 302844 319880 302850 319932
rect 302942 319716 302970 320164
rect 309106 320124 309134 320232
rect 318766 320232 327816 320260
rect 318766 320124 318794 320232
rect 327810 320220 327816 320232
rect 327868 320220 327874 320272
rect 304414 320096 307754 320124
rect 309106 320096 318794 320124
rect 323596 320164 327856 320192
rect 303200 319880 303206 319932
rect 303258 319880 303264 319932
rect 303292 319880 303298 319932
rect 303350 319880 303356 319932
rect 303476 319880 303482 319932
rect 303534 319880 303540 319932
rect 304120 319920 304126 319932
rect 303908 319892 304126 319920
rect 302574 319688 302970 319716
rect 302200 319676 302206 319688
rect 298646 319648 298652 319660
rect 296916 319620 298652 319648
rect 298646 319608 298652 319620
rect 298704 319608 298710 319660
rect 301130 319608 301136 319660
rect 301188 319608 301194 319660
rect 301314 319608 301320 319660
rect 301372 319608 301378 319660
rect 302694 319608 302700 319660
rect 302752 319648 302758 319660
rect 303218 319648 303246 319880
rect 302752 319620 303246 319648
rect 302752 319608 302758 319620
rect 291562 319540 291568 319592
rect 291620 319580 291626 319592
rect 291930 319580 291936 319592
rect 291620 319552 291936 319580
rect 291620 319540 291626 319552
rect 291930 319540 291936 319552
rect 291988 319540 291994 319592
rect 292574 319540 292580 319592
rect 292632 319580 292638 319592
rect 294966 319580 294972 319592
rect 292632 319552 294972 319580
rect 292632 319540 292638 319552
rect 294966 319540 294972 319552
rect 295024 319540 295030 319592
rect 295702 319540 295708 319592
rect 295760 319580 295766 319592
rect 295760 319552 296576 319580
rect 295760 319540 295766 319552
rect 290056 319484 290780 319512
rect 290056 319472 290062 319484
rect 291378 319472 291384 319524
rect 291436 319512 291442 319524
rect 294230 319512 294236 319524
rect 291436 319484 294236 319512
rect 291436 319472 291442 319484
rect 294230 319472 294236 319484
rect 294288 319472 294294 319524
rect 295610 319472 295616 319524
rect 295668 319512 295674 319524
rect 296438 319512 296444 319524
rect 295668 319484 296444 319512
rect 295668 319472 295674 319484
rect 296438 319472 296444 319484
rect 296496 319472 296502 319524
rect 296548 319512 296576 319552
rect 297266 319540 297272 319592
rect 297324 319580 297330 319592
rect 297450 319580 297456 319592
rect 297324 319552 297456 319580
rect 297324 319540 297330 319552
rect 297450 319540 297456 319552
rect 297508 319540 297514 319592
rect 299474 319540 299480 319592
rect 299532 319580 299538 319592
rect 299658 319580 299664 319592
rect 299532 319552 299664 319580
rect 299532 319540 299538 319552
rect 299658 319540 299664 319552
rect 299716 319540 299722 319592
rect 303062 319540 303068 319592
rect 303120 319580 303126 319592
rect 303310 319580 303338 319880
rect 303494 319728 303522 319880
rect 303908 319728 303936 319892
rect 304120 319880 304126 319892
rect 304178 319880 304184 319932
rect 304304 319852 304310 319864
rect 304092 319824 304310 319852
rect 304092 319796 304120 319824
rect 304304 319812 304310 319824
rect 304362 319812 304368 319864
rect 304074 319744 304080 319796
rect 304132 319744 304138 319796
rect 303430 319676 303436 319728
rect 303488 319688 303522 319728
rect 303488 319676 303494 319688
rect 303890 319676 303896 319728
rect 303948 319676 303954 319728
rect 303120 319552 303338 319580
rect 303120 319540 303126 319552
rect 304414 319512 304442 320096
rect 307726 319988 307754 320096
rect 308508 320028 311894 320056
rect 308508 319988 308536 320028
rect 305702 319960 307616 319988
rect 307726 319960 308536 319988
rect 311866 319988 311894 320028
rect 323596 319988 323624 320164
rect 327718 320124 327724 320136
rect 311866 319960 323624 319988
rect 325114 320096 327724 320124
rect 305702 319932 305730 319960
rect 304672 319920 304678 319932
rect 304644 319880 304678 319920
rect 304730 319880 304736 319932
rect 305684 319880 305690 319932
rect 305742 319880 305748 319932
rect 306512 319880 306518 319932
rect 306570 319880 306576 319932
rect 306788 319880 306794 319932
rect 306846 319920 306852 319932
rect 307018 319920 307024 319932
rect 306846 319892 307024 319920
rect 306846 319880 306852 319892
rect 307018 319880 307024 319892
rect 307076 319880 307082 319932
rect 304644 319796 304672 319880
rect 304626 319744 304632 319796
rect 304684 319744 304690 319796
rect 306530 319716 306558 319880
rect 307478 319716 307484 319728
rect 306530 319688 307484 319716
rect 307478 319676 307484 319688
rect 307536 319676 307542 319728
rect 307588 319716 307616 319960
rect 325114 319932 325142 320096
rect 327718 320084 327724 320096
rect 327776 320084 327782 320136
rect 327534 320056 327540 320068
rect 327138 320028 327540 320056
rect 327138 319932 327166 320028
rect 327534 320016 327540 320028
rect 327592 320016 327598 320068
rect 327828 320056 327856 320164
rect 328362 320152 328368 320204
rect 328420 320192 328426 320204
rect 332686 320192 332692 320204
rect 328420 320164 332692 320192
rect 328420 320152 328426 320164
rect 332686 320152 332692 320164
rect 332744 320152 332750 320204
rect 327828 320028 328454 320056
rect 307726 319892 308490 319920
rect 307726 319716 307754 319892
rect 308462 319852 308490 319892
rect 308904 319880 308910 319932
rect 308962 319880 308968 319932
rect 309272 319880 309278 319932
rect 309330 319920 309336 319932
rect 310100 319920 310106 319932
rect 309330 319892 309456 319920
rect 309330 319880 309336 319892
rect 308462 319824 308812 319852
rect 307588 319688 307754 319716
rect 306098 319608 306104 319660
rect 306156 319648 306162 319660
rect 307938 319648 307944 319660
rect 306156 319620 307944 319648
rect 306156 319608 306162 319620
rect 307938 319608 307944 319620
rect 307996 319608 308002 319660
rect 308784 319648 308812 319824
rect 308922 319728 308950 319880
rect 309428 319728 309456 319892
rect 309520 319892 310106 319920
rect 309520 319864 309548 319892
rect 310100 319880 310106 319892
rect 310158 319880 310164 319932
rect 310744 319880 310750 319932
rect 310802 319920 310808 319932
rect 310802 319880 310836 319920
rect 312308 319880 312314 319932
rect 312366 319880 312372 319932
rect 313044 319920 313050 319932
rect 312924 319892 313050 319920
rect 309502 319812 309508 319864
rect 309560 319812 309566 319864
rect 310652 319812 310658 319864
rect 310710 319852 310716 319864
rect 310710 319812 310744 319852
rect 310716 319728 310744 319812
rect 310808 319796 310836 319880
rect 311940 319812 311946 319864
rect 311998 319812 312004 319864
rect 310790 319744 310796 319796
rect 310848 319744 310854 319796
rect 308858 319676 308864 319728
rect 308916 319688 308950 319728
rect 308916 319676 308922 319688
rect 309410 319676 309416 319728
rect 309468 319676 309474 319728
rect 310698 319676 310704 319728
rect 310756 319676 310762 319728
rect 311958 319660 311986 319812
rect 308784 319620 309088 319648
rect 307110 319540 307116 319592
rect 307168 319580 307174 319592
rect 307294 319580 307300 319592
rect 307168 319552 307300 319580
rect 307168 319540 307174 319552
rect 307294 319540 307300 319552
rect 307352 319540 307358 319592
rect 307662 319540 307668 319592
rect 307720 319580 307726 319592
rect 307846 319580 307852 319592
rect 307720 319552 307852 319580
rect 307720 319540 307726 319552
rect 307846 319540 307852 319552
rect 307904 319540 307910 319592
rect 308674 319540 308680 319592
rect 308732 319580 308738 319592
rect 308950 319580 308956 319592
rect 308732 319552 308956 319580
rect 308732 319540 308738 319552
rect 308950 319540 308956 319552
rect 309008 319540 309014 319592
rect 309060 319580 309088 319620
rect 310882 319608 310888 319660
rect 310940 319648 310946 319660
rect 311342 319648 311348 319660
rect 310940 319620 311348 319648
rect 310940 319608 310946 319620
rect 311342 319608 311348 319620
rect 311400 319608 311406 319660
rect 311894 319608 311900 319660
rect 311952 319620 311986 319660
rect 312326 319648 312354 319880
rect 312924 319660 312952 319892
rect 313044 319880 313050 319892
rect 313102 319880 313108 319932
rect 314240 319920 314246 319932
rect 313568 319892 314246 319920
rect 313568 319728 313596 319892
rect 314240 319880 314246 319892
rect 314298 319880 314304 319932
rect 314516 319880 314522 319932
rect 314574 319880 314580 319932
rect 315252 319880 315258 319932
rect 315310 319920 315316 319932
rect 315310 319892 315758 319920
rect 315310 319880 315316 319892
rect 313550 319676 313556 319728
rect 313608 319676 313614 319728
rect 313826 319676 313832 319728
rect 313884 319716 313890 319728
rect 314534 319716 314562 319880
rect 314608 319812 314614 319864
rect 314666 319812 314672 319864
rect 313884 319688 314562 319716
rect 313884 319676 313890 319688
rect 312446 319648 312452 319660
rect 312326 319620 312452 319648
rect 311952 319608 311958 319620
rect 312446 319608 312452 319620
rect 312504 319608 312510 319660
rect 312906 319608 312912 319660
rect 312964 319608 312970 319660
rect 314378 319608 314384 319660
rect 314436 319648 314442 319660
rect 314626 319648 314654 319812
rect 315730 319660 315758 319892
rect 316080 319880 316086 319932
rect 316138 319880 316144 319932
rect 317368 319880 317374 319932
rect 317426 319880 317432 319932
rect 317552 319880 317558 319932
rect 317610 319920 317616 319932
rect 317610 319892 317736 319920
rect 317610 319880 317616 319892
rect 316098 319784 316126 319880
rect 314436 319620 314654 319648
rect 314436 319608 314442 319620
rect 315666 319608 315672 319660
rect 315724 319620 315758 319660
rect 316052 319756 316126 319784
rect 316052 319648 316080 319756
rect 316862 319648 316868 319660
rect 316052 319620 316868 319648
rect 315724 319608 315730 319620
rect 316862 319608 316868 319620
rect 316920 319608 316926 319660
rect 317230 319608 317236 319660
rect 317288 319648 317294 319660
rect 317386 319648 317414 319880
rect 317708 319660 317736 319892
rect 318656 319880 318662 319932
rect 318714 319920 318720 319932
rect 318714 319880 318748 319920
rect 319208 319880 319214 319932
rect 319266 319880 319272 319932
rect 319392 319880 319398 319932
rect 319450 319880 319456 319932
rect 320312 319880 320318 319932
rect 320370 319880 320376 319932
rect 320542 319880 320548 319932
rect 320600 319880 320606 319932
rect 321140 319880 321146 319932
rect 321198 319920 321204 319932
rect 321198 319892 321324 319920
rect 321198 319880 321204 319892
rect 318720 319660 318748 319880
rect 318840 319852 318846 319864
rect 318812 319812 318846 319852
rect 318898 319812 318904 319864
rect 318812 319660 318840 319812
rect 319226 319660 319254 319880
rect 319410 319660 319438 319880
rect 319944 319812 319950 319864
rect 320002 319812 320008 319864
rect 319962 319660 319990 319812
rect 320330 319728 320358 319880
rect 320560 319796 320588 319880
rect 320542 319744 320548 319796
rect 320600 319744 320606 319796
rect 320330 319688 320364 319728
rect 320358 319676 320364 319688
rect 320416 319676 320422 319728
rect 321296 319660 321324 319892
rect 324038 319880 324044 319932
rect 324096 319880 324102 319932
rect 325096 319880 325102 319932
rect 325154 319880 325160 319932
rect 325648 319880 325654 319932
rect 325706 319880 325712 319932
rect 327120 319880 327126 319932
rect 327178 319880 327184 319932
rect 322152 319812 322158 319864
rect 322210 319812 322216 319864
rect 322170 319728 322198 319812
rect 322170 319688 322204 319728
rect 322198 319676 322204 319688
rect 322256 319676 322262 319728
rect 323026 319676 323032 319728
rect 323084 319716 323090 319728
rect 323210 319716 323216 319728
rect 323084 319688 323216 319716
rect 323084 319676 323090 319688
rect 323210 319676 323216 319688
rect 323268 319676 323274 319728
rect 323946 319676 323952 319728
rect 324004 319716 324010 319728
rect 324056 319716 324084 319880
rect 324544 319852 324550 319864
rect 324332 319824 324550 319852
rect 324332 319796 324360 319824
rect 324544 319812 324550 319824
rect 324602 319812 324608 319864
rect 325666 319852 325694 319880
rect 325160 319824 325694 319852
rect 324314 319744 324320 319796
rect 324372 319744 324378 319796
rect 325160 319728 325188 319824
rect 325740 319812 325746 319864
rect 325798 319852 325804 319864
rect 327626 319852 327632 319864
rect 325798 319824 327632 319852
rect 325798 319812 325804 319824
rect 327626 319812 327632 319824
rect 327684 319812 327690 319864
rect 328426 319784 328454 320028
rect 346578 319784 346584 319796
rect 328426 319756 346584 319784
rect 346578 319744 346584 319756
rect 346636 319744 346642 319796
rect 324004 319688 324084 319716
rect 324004 319676 324010 319688
rect 325142 319676 325148 319728
rect 325200 319676 325206 319728
rect 328362 319716 328368 319728
rect 325620 319688 328368 319716
rect 317288 319620 317414 319648
rect 317288 319608 317294 319620
rect 317690 319608 317696 319660
rect 317748 319608 317754 319660
rect 318702 319608 318708 319660
rect 318760 319608 318766 319660
rect 318794 319608 318800 319660
rect 318852 319608 318858 319660
rect 319226 319620 319260 319660
rect 319254 319608 319260 319620
rect 319312 319608 319318 319660
rect 319346 319608 319352 319660
rect 319404 319620 319438 319660
rect 319404 319608 319410 319620
rect 319898 319608 319904 319660
rect 319956 319620 319990 319660
rect 319956 319608 319962 319620
rect 321278 319608 321284 319660
rect 321336 319608 321342 319660
rect 322842 319608 322848 319660
rect 322900 319648 322906 319660
rect 325620 319648 325648 319688
rect 328362 319676 328368 319688
rect 328420 319676 328426 319728
rect 322900 319620 325648 319648
rect 322900 319608 322906 319620
rect 326522 319608 326528 319660
rect 326580 319648 326586 319660
rect 326706 319648 326712 319660
rect 326580 319620 326712 319648
rect 326580 319608 326586 319620
rect 326706 319608 326712 319620
rect 326764 319608 326770 319660
rect 327810 319608 327816 319660
rect 327868 319648 327874 319660
rect 359182 319648 359188 319660
rect 327868 319620 359188 319648
rect 327868 319608 327874 319620
rect 359182 319608 359188 319620
rect 359240 319608 359246 319660
rect 330754 319580 330760 319592
rect 309060 319552 330760 319580
rect 330754 319540 330760 319552
rect 330812 319540 330818 319592
rect 296548 319484 304442 319512
rect 304534 319472 304540 319524
rect 304592 319512 304598 319524
rect 304718 319512 304724 319524
rect 304592 319484 304724 319512
rect 304592 319472 304598 319484
rect 304718 319472 304724 319484
rect 304776 319472 304782 319524
rect 306466 319472 306472 319524
rect 306524 319512 306530 319524
rect 330846 319512 330852 319524
rect 306524 319484 330852 319512
rect 306524 319472 306530 319484
rect 330846 319472 330852 319484
rect 330904 319472 330910 319524
rect 288250 319404 288256 319456
rect 288308 319444 288314 319456
rect 288526 319444 288532 319456
rect 288308 319416 288532 319444
rect 288308 319404 288314 319416
rect 288526 319404 288532 319416
rect 288584 319404 288590 319456
rect 289262 319404 289268 319456
rect 289320 319444 289326 319456
rect 294966 319444 294972 319456
rect 289320 319416 294972 319444
rect 289320 319404 289326 319416
rect 294966 319404 294972 319416
rect 295024 319404 295030 319456
rect 295426 319404 295432 319456
rect 295484 319444 295490 319456
rect 343634 319444 343640 319456
rect 295484 319416 343640 319444
rect 295484 319404 295490 319416
rect 343634 319404 343640 319416
rect 343692 319404 343698 319456
rect 291194 319376 291200 319388
rect 287716 319348 291200 319376
rect 291194 319336 291200 319348
rect 291252 319336 291258 319388
rect 291562 319336 291568 319388
rect 291620 319376 291626 319388
rect 292298 319376 292304 319388
rect 291620 319348 292304 319376
rect 291620 319336 291626 319348
rect 292298 319336 292304 319348
rect 292356 319336 292362 319388
rect 293678 319336 293684 319388
rect 293736 319376 293742 319388
rect 352466 319376 352472 319388
rect 293736 319348 352472 319376
rect 293736 319336 293742 319348
rect 352466 319336 352472 319348
rect 352524 319336 352530 319388
rect 278498 319268 278504 319320
rect 278556 319308 278562 319320
rect 292114 319308 292120 319320
rect 278556 319280 292120 319308
rect 278556 319268 278562 319280
rect 292114 319268 292120 319280
rect 292172 319268 292178 319320
rect 295242 319268 295248 319320
rect 295300 319308 295306 319320
rect 295794 319308 295800 319320
rect 295300 319280 295800 319308
rect 295300 319268 295306 319280
rect 295794 319268 295800 319280
rect 295852 319308 295858 319320
rect 354398 319308 354404 319320
rect 295852 319280 354404 319308
rect 295852 319268 295858 319280
rect 354398 319268 354404 319280
rect 354456 319268 354462 319320
rect 269758 319200 269764 319252
rect 269816 319240 269822 319252
rect 271506 319240 271512 319252
rect 269816 319212 271512 319240
rect 269816 319200 269822 319212
rect 271506 319200 271512 319212
rect 271564 319240 271570 319252
rect 292942 319240 292948 319252
rect 271564 319212 292948 319240
rect 271564 319200 271570 319212
rect 292942 319200 292948 319212
rect 293000 319200 293006 319252
rect 294322 319200 294328 319252
rect 294380 319240 294386 319252
rect 353386 319240 353392 319252
rect 294380 319212 353392 319240
rect 294380 319200 294386 319212
rect 353386 319200 353392 319212
rect 353444 319200 353450 319252
rect 282914 319132 282920 319184
rect 282972 319172 282978 319184
rect 284202 319172 284208 319184
rect 282972 319144 284208 319172
rect 282972 319132 282978 319144
rect 284202 319132 284208 319144
rect 284260 319132 284266 319184
rect 284754 319132 284760 319184
rect 284812 319172 284818 319184
rect 344094 319172 344100 319184
rect 284812 319144 344100 319172
rect 284812 319132 284818 319144
rect 344094 319132 344100 319144
rect 344152 319132 344158 319184
rect 295886 319104 295892 319116
rect 273226 319076 295892 319104
rect 272426 318996 272432 319048
rect 272484 319036 272490 319048
rect 273226 319036 273254 319076
rect 295886 319064 295892 319076
rect 295944 319064 295950 319116
rect 295978 319064 295984 319116
rect 296036 319104 296042 319116
rect 352098 319104 352104 319116
rect 296036 319076 352104 319104
rect 296036 319064 296042 319076
rect 352098 319064 352104 319076
rect 352156 319064 352162 319116
rect 272484 319008 273254 319036
rect 272484 318996 272490 319008
rect 275462 318996 275468 319048
rect 275520 319036 275526 319048
rect 282914 319036 282920 319048
rect 275520 319008 282920 319036
rect 275520 318996 275526 319008
rect 282914 318996 282920 319008
rect 282972 318996 282978 319048
rect 283742 318996 283748 319048
rect 283800 319036 283806 319048
rect 299566 319036 299572 319048
rect 283800 319008 299572 319036
rect 283800 318996 283806 319008
rect 299566 318996 299572 319008
rect 299624 318996 299630 319048
rect 300210 318996 300216 319048
rect 300268 319036 300274 319048
rect 308950 319036 308956 319048
rect 300268 319008 308956 319036
rect 300268 318996 300274 319008
rect 308950 318996 308956 319008
rect 309008 318996 309014 319048
rect 309686 318996 309692 319048
rect 309744 319036 309750 319048
rect 359734 319036 359740 319048
rect 309744 319008 359740 319036
rect 309744 318996 309750 319008
rect 359734 318996 359740 319008
rect 359792 318996 359798 319048
rect 287054 318968 287060 318980
rect 273226 318940 287060 318968
rect 208210 318860 208216 318912
rect 208268 318900 208274 318912
rect 273226 318900 273254 318940
rect 287054 318928 287060 318940
rect 287112 318968 287118 318980
rect 288342 318968 288348 318980
rect 287112 318940 288348 318968
rect 287112 318928 287118 318940
rect 288342 318928 288348 318940
rect 288400 318928 288406 318980
rect 288526 318928 288532 318980
rect 288584 318968 288590 318980
rect 289446 318968 289452 318980
rect 288584 318940 289452 318968
rect 288584 318928 288590 318940
rect 289446 318928 289452 318940
rect 289504 318968 289510 318980
rect 348786 318968 348792 318980
rect 289504 318940 348792 318968
rect 289504 318928 289510 318940
rect 348786 318928 348792 318940
rect 348844 318928 348850 318980
rect 208268 318872 273254 318900
rect 208268 318860 208274 318872
rect 274266 318860 274272 318912
rect 274324 318900 274330 318912
rect 280522 318900 280528 318912
rect 274324 318872 280528 318900
rect 274324 318860 274330 318872
rect 280522 318860 280528 318872
rect 280580 318860 280586 318912
rect 280890 318860 280896 318912
rect 280948 318900 280954 318912
rect 294322 318900 294328 318912
rect 280948 318872 294328 318900
rect 280948 318860 280954 318872
rect 294322 318860 294328 318872
rect 294380 318860 294386 318912
rect 294966 318860 294972 318912
rect 295024 318900 295030 318912
rect 301682 318900 301688 318912
rect 295024 318872 301688 318900
rect 295024 318860 295030 318872
rect 301682 318860 301688 318872
rect 301740 318860 301746 318912
rect 306466 318900 306472 318912
rect 306346 318872 306472 318900
rect 276658 318792 276664 318844
rect 276716 318832 276722 318844
rect 278498 318832 278504 318844
rect 276716 318804 278504 318832
rect 276716 318792 276722 318804
rect 278498 318792 278504 318804
rect 278556 318792 278562 318844
rect 280706 318792 280712 318844
rect 280764 318832 280770 318844
rect 283742 318832 283748 318844
rect 280764 318804 283748 318832
rect 280764 318792 280770 318804
rect 283742 318792 283748 318804
rect 283800 318792 283806 318844
rect 283834 318792 283840 318844
rect 283892 318832 283898 318844
rect 289446 318832 289452 318844
rect 283892 318804 289452 318832
rect 283892 318792 283898 318804
rect 289446 318792 289452 318804
rect 289504 318792 289510 318844
rect 290182 318792 290188 318844
rect 290240 318832 290246 318844
rect 295426 318832 295432 318844
rect 290240 318804 295432 318832
rect 290240 318792 290246 318804
rect 295426 318792 295432 318804
rect 295484 318792 295490 318844
rect 296438 318792 296444 318844
rect 296496 318832 296502 318844
rect 296622 318832 296628 318844
rect 296496 318804 296628 318832
rect 296496 318792 296502 318804
rect 296622 318792 296628 318804
rect 296680 318792 296686 318844
rect 298922 318792 298928 318844
rect 298980 318832 298986 318844
rect 299106 318832 299112 318844
rect 298980 318804 299112 318832
rect 298980 318792 298986 318804
rect 299106 318792 299112 318804
rect 299164 318792 299170 318844
rect 299658 318792 299664 318844
rect 299716 318832 299722 318844
rect 306346 318832 306374 318872
rect 306466 318860 306472 318872
rect 306524 318860 306530 318912
rect 307846 318860 307852 318912
rect 307904 318900 307910 318912
rect 308490 318900 308496 318912
rect 307904 318872 308496 318900
rect 307904 318860 307910 318872
rect 308490 318860 308496 318872
rect 308548 318860 308554 318912
rect 308950 318860 308956 318912
rect 309008 318900 309014 318912
rect 361482 318900 361488 318912
rect 309008 318872 361488 318900
rect 309008 318860 309014 318872
rect 361482 318860 361488 318872
rect 361540 318860 361546 318912
rect 299716 318804 306374 318832
rect 299716 318792 299722 318804
rect 310882 318792 310888 318844
rect 310940 318832 310946 318844
rect 311250 318832 311256 318844
rect 310940 318804 311256 318832
rect 310940 318792 310946 318804
rect 311250 318792 311256 318804
rect 311308 318792 311314 318844
rect 320174 318792 320180 318844
rect 320232 318832 320238 318844
rect 320542 318832 320548 318844
rect 320232 318804 320548 318832
rect 320232 318792 320238 318804
rect 320542 318792 320548 318804
rect 320600 318792 320606 318844
rect 324222 318792 324228 318844
rect 324280 318832 324286 318844
rect 330938 318832 330944 318844
rect 324280 318804 330944 318832
rect 324280 318792 324286 318804
rect 330938 318792 330944 318804
rect 330996 318792 331002 318844
rect 253750 318724 253756 318776
rect 253808 318764 253814 318776
rect 256602 318764 256608 318776
rect 253808 318736 256608 318764
rect 253808 318724 253814 318736
rect 256602 318724 256608 318736
rect 256660 318764 256666 318776
rect 283374 318764 283380 318776
rect 256660 318736 283380 318764
rect 256660 318724 256666 318736
rect 283374 318724 283380 318736
rect 283432 318724 283438 318776
rect 284846 318724 284852 318776
rect 284904 318764 284910 318776
rect 284904 318736 285996 318764
rect 284904 318724 284910 318736
rect 280982 318656 280988 318708
rect 281040 318696 281046 318708
rect 285766 318696 285772 318708
rect 281040 318668 285772 318696
rect 281040 318656 281046 318668
rect 285766 318656 285772 318668
rect 285824 318656 285830 318708
rect 272610 318588 272616 318640
rect 272668 318628 272674 318640
rect 272978 318628 272984 318640
rect 272668 318600 272984 318628
rect 272668 318588 272674 318600
rect 272978 318588 272984 318600
rect 273036 318628 273042 318640
rect 285858 318628 285864 318640
rect 273036 318600 285864 318628
rect 273036 318588 273042 318600
rect 285858 318588 285864 318600
rect 285916 318588 285922 318640
rect 285968 318628 285996 318736
rect 287054 318724 287060 318776
rect 287112 318764 287118 318776
rect 287238 318764 287244 318776
rect 287112 318736 287244 318764
rect 287112 318724 287118 318736
rect 287238 318724 287244 318736
rect 287296 318724 287302 318776
rect 287698 318724 287704 318776
rect 287756 318764 287762 318776
rect 287882 318764 287888 318776
rect 287756 318736 287888 318764
rect 287756 318724 287762 318736
rect 287882 318724 287888 318736
rect 287940 318724 287946 318776
rect 290366 318724 290372 318776
rect 290424 318764 290430 318776
rect 290424 318736 292068 318764
rect 290424 318724 290430 318736
rect 287606 318656 287612 318708
rect 287664 318696 287670 318708
rect 291838 318696 291844 318708
rect 287664 318668 291844 318696
rect 287664 318656 287670 318668
rect 291838 318656 291844 318668
rect 291896 318656 291902 318708
rect 292040 318696 292068 318736
rect 292574 318724 292580 318776
rect 292632 318764 292638 318776
rect 295978 318764 295984 318776
rect 292632 318736 295984 318764
rect 292632 318724 292638 318736
rect 295978 318724 295984 318736
rect 296036 318724 296042 318776
rect 296990 318724 296996 318776
rect 297048 318764 297054 318776
rect 302326 318764 302332 318776
rect 297048 318736 302332 318764
rect 297048 318724 297054 318736
rect 302326 318724 302332 318736
rect 302384 318724 302390 318776
rect 306650 318724 306656 318776
rect 306708 318764 306714 318776
rect 310698 318764 310704 318776
rect 306708 318736 310704 318764
rect 306708 318724 306714 318736
rect 310698 318724 310704 318736
rect 310756 318724 310762 318776
rect 310974 318724 310980 318776
rect 311032 318764 311038 318776
rect 311032 318736 311894 318764
rect 311032 318724 311038 318736
rect 297266 318696 297272 318708
rect 292040 318668 297272 318696
rect 297266 318656 297272 318668
rect 297324 318656 297330 318708
rect 298002 318656 298008 318708
rect 298060 318696 298066 318708
rect 298922 318696 298928 318708
rect 298060 318668 298928 318696
rect 298060 318656 298066 318668
rect 298922 318656 298928 318668
rect 298980 318656 298986 318708
rect 304442 318656 304448 318708
rect 304500 318696 304506 318708
rect 307662 318696 307668 318708
rect 304500 318668 307668 318696
rect 304500 318656 304506 318668
rect 307662 318656 307668 318668
rect 307720 318656 307726 318708
rect 311866 318696 311894 318736
rect 316126 318724 316132 318776
rect 316184 318764 316190 318776
rect 316184 318736 324544 318764
rect 316184 318724 316190 318736
rect 322842 318696 322848 318708
rect 311866 318668 322848 318696
rect 322842 318656 322848 318668
rect 322900 318656 322906 318708
rect 324222 318696 324228 318708
rect 323136 318668 324228 318696
rect 291378 318628 291384 318640
rect 285968 318600 291384 318628
rect 291378 318588 291384 318600
rect 291436 318588 291442 318640
rect 292206 318588 292212 318640
rect 292264 318628 292270 318640
rect 292264 318600 302234 318628
rect 292264 318588 292270 318600
rect 269022 318520 269028 318572
rect 269080 318560 269086 318572
rect 269080 318532 273254 318560
rect 269080 318520 269086 318532
rect 273226 318424 273254 318532
rect 280798 318520 280804 318572
rect 280856 318560 280862 318572
rect 286594 318560 286600 318572
rect 280856 318532 286600 318560
rect 280856 318520 280862 318532
rect 286594 318520 286600 318532
rect 286652 318520 286658 318572
rect 287698 318520 287704 318572
rect 287756 318560 287762 318572
rect 296254 318560 296260 318572
rect 287756 318532 296260 318560
rect 287756 318520 287762 318532
rect 296254 318520 296260 318532
rect 296312 318520 296318 318572
rect 299658 318520 299664 318572
rect 299716 318560 299722 318572
rect 300210 318560 300216 318572
rect 299716 318532 300216 318560
rect 299716 318520 299722 318532
rect 300210 318520 300216 318532
rect 300268 318520 300274 318572
rect 302206 318560 302234 318600
rect 311158 318588 311164 318640
rect 311216 318628 311222 318640
rect 323136 318628 323164 318668
rect 324222 318656 324228 318668
rect 324280 318656 324286 318708
rect 311216 318600 323164 318628
rect 311216 318588 311222 318600
rect 323210 318588 323216 318640
rect 323268 318628 323274 318640
rect 324406 318628 324412 318640
rect 323268 318600 324412 318628
rect 323268 318588 323274 318600
rect 324406 318588 324412 318600
rect 324464 318588 324470 318640
rect 324516 318628 324544 318736
rect 324590 318724 324596 318776
rect 324648 318764 324654 318776
rect 329006 318764 329012 318776
rect 324648 318736 329012 318764
rect 324648 318724 324654 318736
rect 329006 318724 329012 318736
rect 329064 318724 329070 318776
rect 329834 318724 329840 318776
rect 329892 318764 329898 318776
rect 330202 318764 330208 318776
rect 329892 318736 330208 318764
rect 329892 318724 329898 318736
rect 330202 318724 330208 318736
rect 330260 318764 330266 318776
rect 331214 318764 331220 318776
rect 330260 318736 331220 318764
rect 330260 318724 330266 318736
rect 331214 318724 331220 318736
rect 331272 318724 331278 318776
rect 324682 318656 324688 318708
rect 324740 318696 324746 318708
rect 329742 318696 329748 318708
rect 324740 318668 329748 318696
rect 324740 318656 324746 318668
rect 329742 318656 329748 318668
rect 329800 318696 329806 318708
rect 331490 318696 331496 318708
rect 329800 318668 331496 318696
rect 329800 318656 329806 318668
rect 331490 318656 331496 318668
rect 331548 318656 331554 318708
rect 329834 318628 329840 318640
rect 324516 318600 329840 318628
rect 329834 318588 329840 318600
rect 329892 318588 329898 318640
rect 330018 318588 330024 318640
rect 330076 318628 330082 318640
rect 331122 318628 331128 318640
rect 330076 318600 331128 318628
rect 330076 318588 330082 318600
rect 331122 318588 331128 318600
rect 331180 318628 331186 318640
rect 333054 318628 333060 318640
rect 331180 318600 333060 318628
rect 331180 318588 331186 318600
rect 333054 318588 333060 318600
rect 333112 318588 333118 318640
rect 333330 318560 333336 318572
rect 302206 318532 333336 318560
rect 333330 318520 333336 318532
rect 333388 318520 333394 318572
rect 277210 318452 277216 318504
rect 277268 318492 277274 318504
rect 296530 318492 296536 318504
rect 277268 318464 296536 318492
rect 277268 318452 277274 318464
rect 296530 318452 296536 318464
rect 296588 318452 296594 318504
rect 298002 318452 298008 318504
rect 298060 318492 298066 318504
rect 305638 318492 305644 318504
rect 298060 318464 305644 318492
rect 298060 318452 298066 318464
rect 305638 318452 305644 318464
rect 305696 318452 305702 318504
rect 309134 318452 309140 318504
rect 309192 318492 309198 318504
rect 317506 318492 317512 318504
rect 309192 318464 317512 318492
rect 309192 318452 309198 318464
rect 317506 318452 317512 318464
rect 317564 318452 317570 318504
rect 320542 318452 320548 318504
rect 320600 318492 320606 318504
rect 320726 318492 320732 318504
rect 320600 318464 320732 318492
rect 320600 318452 320606 318464
rect 320726 318452 320732 318464
rect 320784 318452 320790 318504
rect 323854 318452 323860 318504
rect 323912 318492 323918 318504
rect 324038 318492 324044 318504
rect 323912 318464 324044 318492
rect 323912 318452 323918 318464
rect 324038 318452 324044 318464
rect 324096 318452 324102 318504
rect 288434 318424 288440 318436
rect 273226 318396 288440 318424
rect 288434 318384 288440 318396
rect 288492 318384 288498 318436
rect 290734 318384 290740 318436
rect 290792 318424 290798 318436
rect 291010 318424 291016 318436
rect 290792 318396 291016 318424
rect 290792 318384 290798 318396
rect 291010 318384 291016 318396
rect 291068 318384 291074 318436
rect 292482 318384 292488 318436
rect 292540 318424 292546 318436
rect 332042 318424 332048 318436
rect 292540 318396 332048 318424
rect 292540 318384 292546 318396
rect 332042 318384 332048 318396
rect 332100 318384 332106 318436
rect 256786 318316 256792 318368
rect 256844 318356 256850 318368
rect 257798 318356 257804 318368
rect 256844 318328 257804 318356
rect 256844 318316 256850 318328
rect 257798 318316 257804 318328
rect 257856 318356 257862 318368
rect 283650 318356 283656 318368
rect 257856 318328 283656 318356
rect 257856 318316 257862 318328
rect 283650 318316 283656 318328
rect 283708 318316 283714 318368
rect 284202 318316 284208 318368
rect 284260 318356 284266 318368
rect 290458 318356 290464 318368
rect 284260 318328 290464 318356
rect 284260 318316 284266 318328
rect 290458 318316 290464 318328
rect 290516 318316 290522 318368
rect 290918 318316 290924 318368
rect 290976 318356 290982 318368
rect 327902 318356 327908 318368
rect 290976 318328 327908 318356
rect 290976 318316 290982 318328
rect 327902 318316 327908 318328
rect 327960 318316 327966 318368
rect 328730 318316 328736 318368
rect 328788 318356 328794 318368
rect 365990 318356 365996 318368
rect 328788 318328 365996 318356
rect 328788 318316 328794 318328
rect 365990 318316 365996 318328
rect 366048 318316 366054 318368
rect 244274 318248 244280 318300
rect 244332 318288 244338 318300
rect 281534 318288 281540 318300
rect 244332 318260 281540 318288
rect 244332 318248 244338 318260
rect 281534 318248 281540 318260
rect 281592 318288 281598 318300
rect 282730 318288 282736 318300
rect 281592 318260 282736 318288
rect 281592 318248 281598 318260
rect 282730 318248 282736 318260
rect 282788 318248 282794 318300
rect 283190 318248 283196 318300
rect 283248 318288 283254 318300
rect 284018 318288 284024 318300
rect 283248 318260 284024 318288
rect 283248 318248 283254 318260
rect 284018 318248 284024 318260
rect 284076 318248 284082 318300
rect 285858 318248 285864 318300
rect 285916 318288 285922 318300
rect 286686 318288 286692 318300
rect 285916 318260 286692 318288
rect 285916 318248 285922 318260
rect 286686 318248 286692 318260
rect 286744 318248 286750 318300
rect 288434 318248 288440 318300
rect 288492 318288 288498 318300
rect 297082 318288 297088 318300
rect 288492 318260 297088 318288
rect 288492 318248 288498 318260
rect 297082 318248 297088 318260
rect 297140 318248 297146 318300
rect 315022 318248 315028 318300
rect 315080 318288 315086 318300
rect 315080 318260 327580 318288
rect 315080 318248 315086 318260
rect 327552 318232 327580 318260
rect 328546 318248 328552 318300
rect 328604 318288 328610 318300
rect 365898 318288 365904 318300
rect 328604 318260 365904 318288
rect 328604 318248 328610 318260
rect 365898 318248 365904 318260
rect 365956 318248 365962 318300
rect 247034 318180 247040 318232
rect 247092 318220 247098 318232
rect 256786 318220 256792 318232
rect 247092 318192 256792 318220
rect 247092 318180 247098 318192
rect 256786 318180 256792 318192
rect 256844 318180 256850 318232
rect 272426 318180 272432 318232
rect 272484 318220 272490 318232
rect 272610 318220 272616 318232
rect 272484 318192 272616 318220
rect 272484 318180 272490 318192
rect 272610 318180 272616 318192
rect 272668 318180 272674 318232
rect 281350 318180 281356 318232
rect 281408 318220 281414 318232
rect 281408 318192 281764 318220
rect 281408 318180 281414 318192
rect 242434 318112 242440 318164
rect 242492 318152 242498 318164
rect 281626 318152 281632 318164
rect 242492 318124 281632 318152
rect 242492 318112 242498 318124
rect 281626 318112 281632 318124
rect 281684 318112 281690 318164
rect 281736 318152 281764 318192
rect 282178 318180 282184 318232
rect 282236 318220 282242 318232
rect 291470 318220 291476 318232
rect 282236 318192 291476 318220
rect 282236 318180 282242 318192
rect 291470 318180 291476 318192
rect 291528 318180 291534 318232
rect 291838 318180 291844 318232
rect 291896 318220 291902 318232
rect 293954 318220 293960 318232
rect 291896 318192 293960 318220
rect 291896 318180 291902 318192
rect 293954 318180 293960 318192
rect 294012 318180 294018 318232
rect 294138 318180 294144 318232
rect 294196 318220 294202 318232
rect 295334 318220 295340 318232
rect 294196 318192 295340 318220
rect 294196 318180 294202 318192
rect 295334 318180 295340 318192
rect 295392 318180 295398 318232
rect 313458 318180 313464 318232
rect 313516 318220 313522 318232
rect 324222 318220 324228 318232
rect 313516 318192 324228 318220
rect 313516 318180 313522 318192
rect 324222 318180 324228 318192
rect 324280 318180 324286 318232
rect 327534 318180 327540 318232
rect 327592 318220 327598 318232
rect 328270 318220 328276 318232
rect 327592 318192 328276 318220
rect 327592 318180 327598 318192
rect 328270 318180 328276 318192
rect 328328 318180 328334 318232
rect 328454 318180 328460 318232
rect 328512 318220 328518 318232
rect 368658 318220 368664 318232
rect 328512 318192 368664 318220
rect 328512 318180 328518 318192
rect 368658 318180 368664 318192
rect 368716 318180 368722 318232
rect 281736 318124 284064 318152
rect 206830 318044 206836 318096
rect 206888 318084 206894 318096
rect 269022 318084 269028 318096
rect 206888 318056 269028 318084
rect 206888 318044 206894 318056
rect 269022 318044 269028 318056
rect 269080 318044 269086 318096
rect 271230 318044 271236 318096
rect 271288 318084 271294 318096
rect 271288 318056 273254 318084
rect 271288 318044 271294 318056
rect 273226 317948 273254 318056
rect 283190 318044 283196 318096
rect 283248 318084 283254 318096
rect 283926 318084 283932 318096
rect 283248 318056 283932 318084
rect 283248 318044 283254 318056
rect 283926 318044 283932 318056
rect 283984 318044 283990 318096
rect 284036 318084 284064 318124
rect 285306 318112 285312 318164
rect 285364 318152 285370 318164
rect 299934 318152 299940 318164
rect 285364 318124 299940 318152
rect 285364 318112 285370 318124
rect 299934 318112 299940 318124
rect 299992 318112 299998 318164
rect 316494 318112 316500 318164
rect 316552 318152 316558 318164
rect 316552 318124 328592 318152
rect 316552 318112 316558 318124
rect 286594 318084 286600 318096
rect 284036 318056 286600 318084
rect 286594 318044 286600 318056
rect 286652 318044 286658 318096
rect 286686 318044 286692 318096
rect 286744 318084 286750 318096
rect 298002 318084 298008 318096
rect 286744 318056 298008 318084
rect 286744 318044 286750 318056
rect 298002 318044 298008 318056
rect 298060 318044 298066 318096
rect 328564 318084 328592 318124
rect 328638 318112 328644 318164
rect 328696 318152 328702 318164
rect 371510 318152 371516 318164
rect 328696 318124 371516 318152
rect 328696 318112 328702 318124
rect 371510 318112 371516 318124
rect 371568 318112 371574 318164
rect 330018 318084 330024 318096
rect 328564 318056 330024 318084
rect 330018 318044 330024 318056
rect 330076 318044 330082 318096
rect 330754 318044 330760 318096
rect 330812 318084 330818 318096
rect 381262 318084 381268 318096
rect 330812 318056 381268 318084
rect 330812 318044 330818 318056
rect 381262 318044 381268 318056
rect 381320 318044 381326 318096
rect 277026 317976 277032 318028
rect 277084 318016 277090 318028
rect 287698 318016 287704 318028
rect 277084 317988 287704 318016
rect 277084 317976 277090 317988
rect 287698 317976 287704 317988
rect 287756 317976 287762 318028
rect 289446 317976 289452 318028
rect 289504 318016 289510 318028
rect 289504 317988 290688 318016
rect 289504 317976 289510 317988
rect 281258 317948 281264 317960
rect 273226 317920 281264 317948
rect 281258 317908 281264 317920
rect 281316 317948 281322 317960
rect 289814 317948 289820 317960
rect 281316 317920 289820 317948
rect 281316 317908 281322 317920
rect 289814 317908 289820 317920
rect 289872 317908 289878 317960
rect 290660 317948 290688 317988
rect 292758 317976 292764 318028
rect 292816 318016 292822 318028
rect 293034 318016 293040 318028
rect 292816 317988 293040 318016
rect 292816 317976 292822 317988
rect 293034 317976 293040 317988
rect 293092 317976 293098 318028
rect 297450 318016 297456 318028
rect 293144 317988 297456 318016
rect 293144 317948 293172 317988
rect 297450 317976 297456 317988
rect 297508 317976 297514 318028
rect 303338 317976 303344 318028
rect 303396 318016 303402 318028
rect 303982 318016 303988 318028
rect 303396 317988 303988 318016
rect 303396 317976 303402 317988
rect 303982 317976 303988 317988
rect 304040 317976 304046 318028
rect 331398 317976 331404 318028
rect 331456 318016 331462 318028
rect 354214 318016 354220 318028
rect 331456 317988 354220 318016
rect 331456 317976 331462 317988
rect 354214 317976 354220 317988
rect 354272 317976 354278 318028
rect 290660 317920 293172 317948
rect 293678 317908 293684 317960
rect 293736 317948 293742 317960
rect 346026 317948 346032 317960
rect 293736 317920 346032 317948
rect 293736 317908 293742 317920
rect 346026 317908 346032 317920
rect 346084 317908 346090 317960
rect 257062 317840 257068 317892
rect 257120 317880 257126 317892
rect 257982 317880 257988 317892
rect 257120 317852 257988 317880
rect 257120 317840 257126 317852
rect 257982 317840 257988 317852
rect 258040 317880 258046 317892
rect 285122 317880 285128 317892
rect 258040 317852 285128 317880
rect 258040 317840 258046 317852
rect 285122 317840 285128 317852
rect 285180 317840 285186 317892
rect 286594 317840 286600 317892
rect 286652 317880 286658 317892
rect 296990 317880 296996 317892
rect 286652 317852 296996 317880
rect 286652 317840 286658 317852
rect 296990 317840 296996 317852
rect 297048 317840 297054 317892
rect 297266 317840 297272 317892
rect 297324 317880 297330 317892
rect 332134 317880 332140 317892
rect 297324 317852 332140 317880
rect 297324 317840 297330 317852
rect 332134 317840 332140 317852
rect 332192 317840 332198 317892
rect 265802 317772 265808 317824
rect 265860 317812 265866 317824
rect 283006 317812 283012 317824
rect 265860 317784 283012 317812
rect 265860 317772 265866 317784
rect 283006 317772 283012 317784
rect 283064 317772 283070 317824
rect 290274 317772 290280 317824
rect 290332 317812 290338 317824
rect 332226 317812 332232 317824
rect 290332 317784 332232 317812
rect 290332 317772 290338 317784
rect 332226 317772 332232 317784
rect 332284 317772 332290 317824
rect 270034 317704 270040 317756
rect 270092 317744 270098 317756
rect 275554 317744 275560 317756
rect 270092 317716 275560 317744
rect 270092 317704 270098 317716
rect 275554 317704 275560 317716
rect 275612 317744 275618 317756
rect 293862 317744 293868 317756
rect 275612 317716 293868 317744
rect 275612 317704 275618 317716
rect 293862 317704 293868 317716
rect 293920 317704 293926 317756
rect 299566 317704 299572 317756
rect 299624 317744 299630 317756
rect 300946 317744 300952 317756
rect 299624 317716 300952 317744
rect 299624 317704 299630 317716
rect 300946 317704 300952 317716
rect 301004 317704 301010 317756
rect 303982 317704 303988 317756
rect 304040 317744 304046 317756
rect 307478 317744 307484 317756
rect 304040 317716 307484 317744
rect 304040 317704 304046 317716
rect 307478 317704 307484 317716
rect 307536 317744 307542 317756
rect 311250 317744 311256 317756
rect 307536 317716 311256 317744
rect 307536 317704 307542 317716
rect 311250 317704 311256 317716
rect 311308 317704 311314 317756
rect 324590 317704 324596 317756
rect 324648 317744 324654 317756
rect 324958 317744 324964 317756
rect 324648 317716 324964 317744
rect 324648 317704 324654 317716
rect 324958 317704 324964 317716
rect 325016 317704 325022 317756
rect 284846 317636 284852 317688
rect 284904 317676 284910 317688
rect 285030 317676 285036 317688
rect 284904 317648 285036 317676
rect 284904 317636 284910 317648
rect 285030 317636 285036 317648
rect 285088 317636 285094 317688
rect 286042 317636 286048 317688
rect 286100 317676 286106 317688
rect 287330 317676 287336 317688
rect 286100 317648 287336 317676
rect 286100 317636 286106 317648
rect 287330 317636 287336 317648
rect 287388 317636 287394 317688
rect 291930 317636 291936 317688
rect 291988 317676 291994 317688
rect 292298 317676 292304 317688
rect 291988 317648 292304 317676
rect 291988 317636 291994 317648
rect 292298 317636 292304 317648
rect 292356 317676 292362 317688
rect 333422 317676 333428 317688
rect 292356 317648 333428 317676
rect 292356 317636 292362 317648
rect 333422 317636 333428 317648
rect 333480 317636 333486 317688
rect 282822 317568 282828 317620
rect 282880 317608 282886 317620
rect 288802 317608 288808 317620
rect 282880 317580 288808 317608
rect 282880 317568 282886 317580
rect 288802 317568 288808 317580
rect 288860 317568 288866 317620
rect 296254 317608 296260 317620
rect 292132 317580 296260 317608
rect 279878 317500 279884 317552
rect 279936 317540 279942 317552
rect 292132 317540 292160 317580
rect 296254 317568 296260 317580
rect 296312 317608 296318 317620
rect 296714 317608 296720 317620
rect 296312 317580 296720 317608
rect 296312 317568 296318 317580
rect 296714 317568 296720 317580
rect 296772 317568 296778 317620
rect 299842 317568 299848 317620
rect 299900 317608 299906 317620
rect 300578 317608 300584 317620
rect 299900 317580 300584 317608
rect 299900 317568 299906 317580
rect 300578 317568 300584 317580
rect 300636 317568 300642 317620
rect 300946 317568 300952 317620
rect 301004 317608 301010 317620
rect 302142 317608 302148 317620
rect 301004 317580 302148 317608
rect 301004 317568 301010 317580
rect 302142 317568 302148 317580
rect 302200 317568 302206 317620
rect 314102 317568 314108 317620
rect 314160 317608 314166 317620
rect 314562 317608 314568 317620
rect 314160 317580 314568 317608
rect 314160 317568 314166 317580
rect 314562 317568 314568 317580
rect 314620 317568 314626 317620
rect 325786 317568 325792 317620
rect 325844 317608 325850 317620
rect 326522 317608 326528 317620
rect 325844 317580 326528 317608
rect 325844 317568 325850 317580
rect 326522 317568 326528 317580
rect 326580 317568 326586 317620
rect 327442 317568 327448 317620
rect 327500 317608 327506 317620
rect 329098 317608 329104 317620
rect 327500 317580 329104 317608
rect 327500 317568 327506 317580
rect 329098 317568 329104 317580
rect 329156 317568 329162 317620
rect 279936 317512 292160 317540
rect 279936 317500 279942 317512
rect 295978 317500 295984 317552
rect 296036 317540 296042 317552
rect 299658 317540 299664 317552
rect 296036 317512 299664 317540
rect 296036 317500 296042 317512
rect 299658 317500 299664 317512
rect 299716 317500 299722 317552
rect 314010 317500 314016 317552
rect 314068 317540 314074 317552
rect 317322 317540 317328 317552
rect 314068 317512 317328 317540
rect 314068 317500 314074 317512
rect 317322 317500 317328 317512
rect 317380 317500 317386 317552
rect 321922 317500 321928 317552
rect 321980 317540 321986 317552
rect 328822 317540 328828 317552
rect 321980 317512 328828 317540
rect 321980 317500 321986 317512
rect 328822 317500 328828 317512
rect 328880 317500 328886 317552
rect 276842 317432 276848 317484
rect 276900 317472 276906 317484
rect 277210 317472 277216 317484
rect 276900 317444 277216 317472
rect 276900 317432 276906 317444
rect 277210 317432 277216 317444
rect 277268 317432 277274 317484
rect 280614 317432 280620 317484
rect 280672 317472 280678 317484
rect 280672 317444 284340 317472
rect 280672 317432 280678 317444
rect 268838 317364 268844 317416
rect 268896 317404 268902 317416
rect 269574 317404 269580 317416
rect 268896 317376 269580 317404
rect 268896 317364 268902 317376
rect 269574 317364 269580 317376
rect 269632 317364 269638 317416
rect 281074 317364 281080 317416
rect 281132 317404 281138 317416
rect 283374 317404 283380 317416
rect 281132 317376 283380 317404
rect 281132 317364 281138 317376
rect 283374 317364 283380 317376
rect 283432 317404 283438 317416
rect 284202 317404 284208 317416
rect 283432 317376 284208 317404
rect 283432 317364 283438 317376
rect 284202 317364 284208 317376
rect 284260 317364 284266 317416
rect 284312 317404 284340 317444
rect 285398 317432 285404 317484
rect 285456 317472 285462 317484
rect 286870 317472 286876 317484
rect 285456 317444 286876 317472
rect 285456 317432 285462 317444
rect 286870 317432 286876 317444
rect 286928 317432 286934 317484
rect 286980 317444 288480 317472
rect 286980 317404 287008 317444
rect 284312 317376 287008 317404
rect 287146 317364 287152 317416
rect 287204 317404 287210 317416
rect 288342 317404 288348 317416
rect 287204 317376 288348 317404
rect 287204 317364 287210 317376
rect 288342 317364 288348 317376
rect 288400 317364 288406 317416
rect 288452 317404 288480 317444
rect 290274 317432 290280 317484
rect 290332 317472 290338 317484
rect 290458 317472 290464 317484
rect 290332 317444 290464 317472
rect 290332 317432 290338 317444
rect 290458 317432 290464 317444
rect 290516 317432 290522 317484
rect 297910 317432 297916 317484
rect 297968 317472 297974 317484
rect 298370 317472 298376 317484
rect 297968 317444 298376 317472
rect 297968 317432 297974 317444
rect 298370 317432 298376 317444
rect 298428 317432 298434 317484
rect 302142 317432 302148 317484
rect 302200 317472 302206 317484
rect 304718 317472 304724 317484
rect 302200 317444 304724 317472
rect 302200 317432 302206 317444
rect 304718 317432 304724 317444
rect 304776 317432 304782 317484
rect 307570 317432 307576 317484
rect 307628 317472 307634 317484
rect 307938 317472 307944 317484
rect 307628 317444 307944 317472
rect 307628 317432 307634 317444
rect 307938 317432 307944 317444
rect 307996 317432 308002 317484
rect 313182 317432 313188 317484
rect 313240 317472 313246 317484
rect 314102 317472 314108 317484
rect 313240 317444 314108 317472
rect 313240 317432 313246 317444
rect 314102 317432 314108 317444
rect 314160 317432 314166 317484
rect 320634 317432 320640 317484
rect 320692 317472 320698 317484
rect 327810 317472 327816 317484
rect 320692 317444 327816 317472
rect 320692 317432 320698 317444
rect 327810 317432 327816 317444
rect 327868 317432 327874 317484
rect 298830 317404 298836 317416
rect 288452 317376 298836 317404
rect 298830 317364 298836 317376
rect 298888 317364 298894 317416
rect 325602 317364 325608 317416
rect 325660 317404 325666 317416
rect 394878 317404 394884 317416
rect 325660 317376 394884 317404
rect 325660 317364 325666 317376
rect 394878 317364 394884 317376
rect 394936 317404 394942 317416
rect 395982 317404 395988 317416
rect 394936 317376 395988 317404
rect 394936 317364 394942 317376
rect 395982 317364 395988 317376
rect 396040 317364 396046 317416
rect 270126 317296 270132 317348
rect 270184 317336 270190 317348
rect 297542 317336 297548 317348
rect 270184 317308 297548 317336
rect 270184 317296 270190 317308
rect 297542 317296 297548 317308
rect 297600 317296 297606 317348
rect 322474 317296 322480 317348
rect 322532 317336 322538 317348
rect 322658 317336 322664 317348
rect 322532 317308 322664 317336
rect 322532 317296 322538 317308
rect 322658 317296 322664 317308
rect 322716 317296 322722 317348
rect 329098 317296 329104 317348
rect 329156 317336 329162 317348
rect 330110 317336 330116 317348
rect 329156 317308 330116 317336
rect 329156 317296 329162 317308
rect 330110 317296 330116 317308
rect 330168 317336 330174 317348
rect 389542 317336 389548 317348
rect 330168 317308 389548 317336
rect 330168 317296 330174 317308
rect 389542 317296 389548 317308
rect 389600 317296 389606 317348
rect 278682 317228 278688 317280
rect 278740 317268 278746 317280
rect 298186 317268 298192 317280
rect 278740 317240 298192 317268
rect 278740 317228 278746 317240
rect 298186 317228 298192 317240
rect 298244 317228 298250 317280
rect 323578 317228 323584 317280
rect 323636 317268 323642 317280
rect 324130 317268 324136 317280
rect 323636 317240 324136 317268
rect 323636 317228 323642 317240
rect 324130 317228 324136 317240
rect 324188 317228 324194 317280
rect 326154 317228 326160 317280
rect 326212 317268 326218 317280
rect 332870 317268 332876 317280
rect 326212 317240 332876 317268
rect 326212 317228 326218 317240
rect 332870 317228 332876 317240
rect 332928 317268 332934 317280
rect 333698 317268 333704 317280
rect 332928 317240 333704 317268
rect 332928 317228 332934 317240
rect 333698 317228 333704 317240
rect 333756 317228 333762 317280
rect 340874 317228 340880 317280
rect 340932 317268 340938 317280
rect 341978 317268 341984 317280
rect 340932 317240 341984 317268
rect 340932 317228 340938 317240
rect 341978 317228 341984 317240
rect 342036 317228 342042 317280
rect 279602 317160 279608 317212
rect 279660 317200 279666 317212
rect 299014 317200 299020 317212
rect 279660 317172 299020 317200
rect 279660 317160 279666 317172
rect 299014 317160 299020 317172
rect 299072 317160 299078 317212
rect 309134 317160 309140 317212
rect 309192 317200 309198 317212
rect 309410 317200 309416 317212
rect 309192 317172 309416 317200
rect 309192 317160 309198 317172
rect 309410 317160 309416 317172
rect 309468 317200 309474 317212
rect 328454 317200 328460 317212
rect 309468 317172 328460 317200
rect 309468 317160 309474 317172
rect 328454 317160 328460 317172
rect 328512 317160 328518 317212
rect 291286 317092 291292 317144
rect 291344 317132 291350 317144
rect 292206 317132 292212 317144
rect 291344 317104 292212 317132
rect 291344 317092 291350 317104
rect 292206 317092 292212 317104
rect 292264 317132 292270 317144
rect 293678 317132 293684 317144
rect 292264 317104 293684 317132
rect 292264 317092 292270 317104
rect 293678 317092 293684 317104
rect 293736 317092 293742 317144
rect 299474 317092 299480 317144
rect 299532 317132 299538 317144
rect 307018 317132 307024 317144
rect 299532 317104 307024 317132
rect 299532 317092 299538 317104
rect 307018 317092 307024 317104
rect 307076 317132 307082 317144
rect 328546 317132 328552 317144
rect 307076 317104 328552 317132
rect 307076 317092 307082 317104
rect 328546 317092 328552 317104
rect 328604 317092 328610 317144
rect 328822 317092 328828 317144
rect 328880 317132 328886 317144
rect 329742 317132 329748 317144
rect 328880 317104 329748 317132
rect 328880 317092 328886 317104
rect 329742 317092 329748 317104
rect 329800 317132 329806 317144
rect 339310 317132 339316 317144
rect 329800 317104 339316 317132
rect 329800 317092 329806 317104
rect 339310 317092 339316 317104
rect 339368 317092 339374 317144
rect 277026 317024 277032 317076
rect 277084 317064 277090 317076
rect 303338 317064 303344 317076
rect 277084 317036 303344 317064
rect 277084 317024 277090 317036
rect 303338 317024 303344 317036
rect 303396 317024 303402 317076
rect 317322 317024 317328 317076
rect 317380 317064 317386 317076
rect 340966 317064 340972 317076
rect 317380 317036 340972 317064
rect 317380 317024 317386 317036
rect 340966 317024 340972 317036
rect 341024 317024 341030 317076
rect 277762 316956 277768 317008
rect 277820 316996 277826 317008
rect 278682 316996 278688 317008
rect 277820 316968 278688 316996
rect 277820 316956 277826 316968
rect 278682 316956 278688 316968
rect 278740 316956 278746 317008
rect 279234 316956 279240 317008
rect 279292 316996 279298 317008
rect 309134 316996 309140 317008
rect 279292 316968 309140 316996
rect 279292 316956 279298 316968
rect 309134 316956 309140 316968
rect 309192 316956 309198 317008
rect 317506 316956 317512 317008
rect 317564 316996 317570 317008
rect 340874 316996 340880 317008
rect 317564 316968 340880 316996
rect 317564 316956 317570 316968
rect 340874 316956 340880 316968
rect 340932 316956 340938 317008
rect 275370 316888 275376 316940
rect 275428 316928 275434 316940
rect 309410 316928 309416 316940
rect 275428 316900 309416 316928
rect 275428 316888 275434 316900
rect 309410 316888 309416 316900
rect 309468 316888 309474 316940
rect 321094 316888 321100 316940
rect 321152 316928 321158 316940
rect 321278 316928 321284 316940
rect 321152 316900 321284 316928
rect 321152 316888 321158 316900
rect 321278 316888 321284 316900
rect 321336 316888 321342 316940
rect 324222 316888 324228 316940
rect 324280 316928 324286 316940
rect 328546 316928 328552 316940
rect 324280 316900 328552 316928
rect 324280 316888 324286 316900
rect 328546 316888 328552 316900
rect 328604 316928 328610 316940
rect 329650 316928 329656 316940
rect 328604 316900 329656 316928
rect 328604 316888 328610 316900
rect 329650 316888 329656 316900
rect 329708 316888 329714 316940
rect 213546 316820 213552 316872
rect 213604 316860 213610 316872
rect 270126 316860 270132 316872
rect 213604 316832 270132 316860
rect 213604 316820 213610 316832
rect 270126 316820 270132 316832
rect 270184 316820 270190 316872
rect 273898 316820 273904 316872
rect 273956 316860 273962 316872
rect 311986 316860 311992 316872
rect 273956 316832 311992 316860
rect 273956 316820 273962 316832
rect 311986 316820 311992 316832
rect 312044 316860 312050 316872
rect 324130 316860 324136 316872
rect 312044 316832 324136 316860
rect 312044 316820 312050 316832
rect 324130 316820 324136 316832
rect 324188 316820 324194 316872
rect 328270 316820 328276 316872
rect 328328 316860 328334 316872
rect 341334 316860 341340 316872
rect 328328 316832 341340 316860
rect 328328 316820 328334 316832
rect 341334 316820 341340 316832
rect 341392 316820 341398 316872
rect 347498 316820 347504 316872
rect 347556 316860 347562 316872
rect 362310 316860 362316 316872
rect 347556 316832 362316 316860
rect 347556 316820 347562 316832
rect 362310 316820 362316 316832
rect 362368 316820 362374 316872
rect 212166 316752 212172 316804
rect 212224 316792 212230 316804
rect 280154 316792 280160 316804
rect 212224 316764 280160 316792
rect 212224 316752 212230 316764
rect 280154 316752 280160 316764
rect 280212 316752 280218 316804
rect 309410 316752 309416 316804
rect 309468 316792 309474 316804
rect 309594 316792 309600 316804
rect 309468 316764 309600 316792
rect 309468 316752 309474 316764
rect 309594 316752 309600 316764
rect 309652 316792 309658 316804
rect 324222 316792 324228 316804
rect 309652 316764 324228 316792
rect 309652 316752 309658 316764
rect 324222 316752 324228 316764
rect 324280 316752 324286 316804
rect 325970 316752 325976 316804
rect 326028 316792 326034 316804
rect 326028 316764 348832 316792
rect 326028 316752 326034 316764
rect 348804 316736 348832 316764
rect 212350 316684 212356 316736
rect 212408 316724 212414 316736
rect 296070 316724 296076 316736
rect 212408 316696 296076 316724
rect 212408 316684 212414 316696
rect 296070 316684 296076 316696
rect 296128 316724 296134 316736
rect 296530 316724 296536 316736
rect 296128 316696 296536 316724
rect 296128 316684 296134 316696
rect 296530 316684 296536 316696
rect 296588 316684 296594 316736
rect 312722 316684 312728 316736
rect 312780 316724 312786 316736
rect 347498 316724 347504 316736
rect 312780 316696 347504 316724
rect 312780 316684 312786 316696
rect 347498 316684 347504 316696
rect 347556 316684 347562 316736
rect 348786 316684 348792 316736
rect 348844 316724 348850 316736
rect 385218 316724 385224 316736
rect 348844 316696 385224 316724
rect 348844 316684 348850 316696
rect 385218 316684 385224 316696
rect 385276 316684 385282 316736
rect 395982 316684 395988 316736
rect 396040 316724 396046 316736
rect 527818 316724 527824 316736
rect 396040 316696 527824 316724
rect 396040 316684 396046 316696
rect 527818 316684 527824 316696
rect 527876 316684 527882 316736
rect 275738 316616 275744 316668
rect 275796 316656 275802 316668
rect 276382 316656 276388 316668
rect 275796 316628 276388 316656
rect 275796 316616 275802 316628
rect 276382 316616 276388 316628
rect 276440 316656 276446 316668
rect 295058 316656 295064 316668
rect 276440 316628 295064 316656
rect 276440 316616 276446 316628
rect 295058 316616 295064 316628
rect 295116 316616 295122 316668
rect 298278 316616 298284 316668
rect 298336 316656 298342 316668
rect 299290 316656 299296 316668
rect 298336 316628 299296 316656
rect 298336 316616 298342 316628
rect 299290 316616 299296 316628
rect 299348 316616 299354 316668
rect 304718 316616 304724 316668
rect 304776 316656 304782 316668
rect 336642 316656 336648 316668
rect 304776 316628 336648 316656
rect 304776 316616 304782 316628
rect 336642 316616 336648 316628
rect 336700 316616 336706 316668
rect 272886 316548 272892 316600
rect 272944 316588 272950 316600
rect 276290 316588 276296 316600
rect 272944 316560 276296 316588
rect 272944 316548 272950 316560
rect 276290 316548 276296 316560
rect 276348 316588 276354 316600
rect 304442 316588 304448 316600
rect 276348 316560 304448 316588
rect 276348 316548 276354 316560
rect 304442 316548 304448 316560
rect 304500 316548 304506 316600
rect 317506 316548 317512 316600
rect 317564 316588 317570 316600
rect 317690 316588 317696 316600
rect 317564 316560 317696 316588
rect 317564 316548 317570 316560
rect 317690 316548 317696 316560
rect 317748 316548 317754 316600
rect 319438 316548 319444 316600
rect 319496 316588 319502 316600
rect 320082 316588 320088 316600
rect 319496 316560 320088 316588
rect 319496 316548 319502 316560
rect 320082 316548 320088 316560
rect 320140 316588 320146 316600
rect 378318 316588 378324 316600
rect 320140 316560 378324 316588
rect 320140 316548 320146 316560
rect 378318 316548 378324 316560
rect 378376 316548 378382 316600
rect 296530 316480 296536 316532
rect 296588 316520 296594 316532
rect 355042 316520 355048 316532
rect 296588 316492 355048 316520
rect 296588 316480 296594 316492
rect 355042 316480 355048 316492
rect 355100 316480 355106 316532
rect 303338 316412 303344 316464
rect 303396 316452 303402 316464
rect 305270 316452 305276 316464
rect 303396 316424 305276 316452
rect 303396 316412 303402 316424
rect 305270 316412 305276 316424
rect 305328 316452 305334 316464
rect 329374 316452 329380 316464
rect 305328 316424 329380 316452
rect 305328 316412 305334 316424
rect 329374 316412 329380 316424
rect 329432 316412 329438 316464
rect 278498 316344 278504 316396
rect 278556 316384 278562 316396
rect 303706 316384 303712 316396
rect 278556 316356 303712 316384
rect 278556 316344 278562 316356
rect 303706 316344 303712 316356
rect 303764 316384 303770 316396
rect 304718 316384 304724 316396
rect 303764 316356 304724 316384
rect 303764 316344 303770 316356
rect 304718 316344 304724 316356
rect 304776 316344 304782 316396
rect 316678 316344 316684 316396
rect 316736 316384 316742 316396
rect 329466 316384 329472 316396
rect 316736 316356 329472 316384
rect 316736 316344 316742 316356
rect 329466 316344 329472 316356
rect 329524 316344 329530 316396
rect 304442 316316 304448 316328
rect 299446 316288 304448 316316
rect 294506 316208 294512 316260
rect 294564 316248 294570 316260
rect 294966 316248 294972 316260
rect 294564 316220 294972 316248
rect 294564 316208 294570 316220
rect 294966 316208 294972 316220
rect 295024 316208 295030 316260
rect 298830 316208 298836 316260
rect 298888 316248 298894 316260
rect 299446 316248 299474 316288
rect 304442 316276 304448 316288
rect 304500 316276 304506 316328
rect 312998 316276 313004 316328
rect 313056 316316 313062 316328
rect 313182 316316 313188 316328
rect 313056 316288 313188 316316
rect 313056 316276 313062 316288
rect 313182 316276 313188 316288
rect 313240 316276 313246 316328
rect 321278 316276 321284 316328
rect 321336 316316 321342 316328
rect 321462 316316 321468 316328
rect 321336 316288 321468 316316
rect 321336 316276 321342 316288
rect 321462 316276 321468 316288
rect 321520 316276 321526 316328
rect 324866 316276 324872 316328
rect 324924 316316 324930 316328
rect 325602 316316 325608 316328
rect 324924 316288 325608 316316
rect 324924 316276 324930 316288
rect 325602 316276 325608 316288
rect 325660 316276 325666 316328
rect 298888 316220 299474 316248
rect 299584 316220 299888 316248
rect 298888 316208 298894 316220
rect 272978 316140 272984 316192
rect 273036 316180 273042 316192
rect 299584 316180 299612 316220
rect 273036 316152 299612 316180
rect 299860 316180 299888 316220
rect 300854 316208 300860 316260
rect 300912 316248 300918 316260
rect 301130 316248 301136 316260
rect 300912 316220 301136 316248
rect 300912 316208 300918 316220
rect 301130 316208 301136 316220
rect 301188 316208 301194 316260
rect 304166 316208 304172 316260
rect 304224 316248 304230 316260
rect 304718 316248 304724 316260
rect 304224 316220 304724 316248
rect 304224 316208 304230 316220
rect 304718 316208 304724 316220
rect 304776 316208 304782 316260
rect 306650 316208 306656 316260
rect 306708 316248 306714 316260
rect 307110 316248 307116 316260
rect 306708 316220 307116 316248
rect 306708 316208 306714 316220
rect 307110 316208 307116 316220
rect 307168 316208 307174 316260
rect 311434 316208 311440 316260
rect 311492 316248 311498 316260
rect 311618 316248 311624 316260
rect 311492 316220 311624 316248
rect 311492 316208 311498 316220
rect 311618 316208 311624 316220
rect 311676 316208 311682 316260
rect 313734 316248 313740 316260
rect 312004 316220 313740 316248
rect 312004 316192 312032 316220
rect 313734 316208 313740 316220
rect 313792 316208 313798 316260
rect 316126 316208 316132 316260
rect 316184 316248 316190 316260
rect 316402 316248 316408 316260
rect 316184 316220 316408 316248
rect 316184 316208 316190 316220
rect 316402 316208 316408 316220
rect 316460 316208 316466 316260
rect 311986 316180 311992 316192
rect 299860 316152 311992 316180
rect 273036 316140 273042 316152
rect 311986 316140 311992 316152
rect 312044 316140 312050 316192
rect 312170 316140 312176 316192
rect 312228 316180 312234 316192
rect 312998 316180 313004 316192
rect 312228 316152 313004 316180
rect 312228 316140 312234 316152
rect 312998 316140 313004 316152
rect 313056 316140 313062 316192
rect 313550 316140 313556 316192
rect 313608 316180 313614 316192
rect 314286 316180 314292 316192
rect 313608 316152 314292 316180
rect 313608 316140 313614 316152
rect 314286 316140 314292 316152
rect 314344 316140 314350 316192
rect 315022 316140 315028 316192
rect 315080 316180 315086 316192
rect 315482 316180 315488 316192
rect 315080 316152 315488 316180
rect 315080 316140 315086 316152
rect 315482 316140 315488 316152
rect 315540 316140 315546 316192
rect 320450 316140 320456 316192
rect 320508 316180 320514 316192
rect 321462 316180 321468 316192
rect 320508 316152 321468 316180
rect 320508 316140 320514 316152
rect 321462 316140 321468 316152
rect 321520 316140 321526 316192
rect 321830 316140 321836 316192
rect 321888 316180 321894 316192
rect 322566 316180 322572 316192
rect 321888 316152 322572 316180
rect 321888 316140 321894 316152
rect 322566 316140 322572 316152
rect 322624 316140 322630 316192
rect 285674 316072 285680 316124
rect 285732 316112 285738 316124
rect 286134 316112 286140 316124
rect 285732 316084 286140 316112
rect 285732 316072 285738 316084
rect 286134 316072 286140 316084
rect 286192 316072 286198 316124
rect 303982 316112 303988 316124
rect 292546 316084 299474 316112
rect 282546 316004 282552 316056
rect 282604 316044 282610 316056
rect 292546 316044 292574 316084
rect 282604 316016 292574 316044
rect 282604 316004 282610 316016
rect 294782 316004 294788 316056
rect 294840 316044 294846 316056
rect 295058 316044 295064 316056
rect 294840 316016 295064 316044
rect 294840 316004 294846 316016
rect 295058 316004 295064 316016
rect 295116 316004 295122 316056
rect 299446 316044 299474 316084
rect 299860 316084 303988 316112
rect 299860 316044 299888 316084
rect 303982 316072 303988 316084
rect 304040 316072 304046 316124
rect 304442 316072 304448 316124
rect 304500 316112 304506 316124
rect 323486 316112 323492 316124
rect 304500 316084 323492 316112
rect 304500 316072 304506 316084
rect 323486 316072 323492 316084
rect 323544 316112 323550 316124
rect 323670 316112 323676 316124
rect 323544 316084 323676 316112
rect 323544 316072 323550 316084
rect 323670 316072 323676 316084
rect 323728 316072 323734 316124
rect 299446 316016 299888 316044
rect 299934 316004 299940 316056
rect 299992 316044 299998 316056
rect 300670 316044 300676 316056
rect 299992 316016 300676 316044
rect 299992 316004 299998 316016
rect 300670 316004 300676 316016
rect 300728 316004 300734 316056
rect 302786 316004 302792 316056
rect 302844 316044 302850 316056
rect 303430 316044 303436 316056
rect 302844 316016 303436 316044
rect 302844 316004 302850 316016
rect 303430 316004 303436 316016
rect 303488 316004 303494 316056
rect 304166 316004 304172 316056
rect 304224 316044 304230 316056
rect 304810 316044 304816 316056
rect 304224 316016 304816 316044
rect 304224 316004 304230 316016
rect 304810 316004 304816 316016
rect 304868 316004 304874 316056
rect 305270 316004 305276 316056
rect 305328 316044 305334 316056
rect 305914 316044 305920 316056
rect 305328 316016 305920 316044
rect 305328 316004 305334 316016
rect 305914 316004 305920 316016
rect 305972 316004 305978 316056
rect 306834 316004 306840 316056
rect 306892 316044 306898 316056
rect 307294 316044 307300 316056
rect 306892 316016 307300 316044
rect 306892 316004 306898 316016
rect 307294 316004 307300 316016
rect 307352 316004 307358 316056
rect 308306 316004 308312 316056
rect 308364 316044 308370 316056
rect 309042 316044 309048 316056
rect 308364 316016 309048 316044
rect 308364 316004 308370 316016
rect 309042 316004 309048 316016
rect 309100 316004 309106 316056
rect 310698 316004 310704 316056
rect 310756 316044 310762 316056
rect 311710 316044 311716 316056
rect 310756 316016 311716 316044
rect 310756 316004 310762 316016
rect 311710 316004 311716 316016
rect 311768 316004 311774 316056
rect 312078 316004 312084 316056
rect 312136 316044 312142 316056
rect 312906 316044 312912 316056
rect 312136 316016 312912 316044
rect 312136 316004 312142 316016
rect 312906 316004 312912 316016
rect 312964 316004 312970 316056
rect 313366 316004 313372 316056
rect 313424 316044 313430 316056
rect 314286 316044 314292 316056
rect 313424 316016 314292 316044
rect 313424 316004 313430 316016
rect 314286 316004 314292 316016
rect 314344 316004 314350 316056
rect 314838 316004 314844 316056
rect 314896 316044 314902 316056
rect 315850 316044 315856 316056
rect 314896 316016 315856 316044
rect 314896 316004 314902 316016
rect 315850 316004 315856 316016
rect 315908 316004 315914 316056
rect 316218 316004 316224 316056
rect 316276 316044 316282 316056
rect 316954 316044 316960 316056
rect 316276 316016 316960 316044
rect 316276 316004 316282 316016
rect 316954 316004 316960 316016
rect 317012 316004 317018 316056
rect 324590 316004 324596 316056
rect 324648 316044 324654 316056
rect 325142 316044 325148 316056
rect 324648 316016 325148 316044
rect 324648 316004 324654 316016
rect 325142 316004 325148 316016
rect 325200 316004 325206 316056
rect 264790 315936 264796 315988
rect 264848 315976 264854 315988
rect 283466 315976 283472 315988
rect 264848 315948 283472 315976
rect 264848 315936 264854 315948
rect 283466 315936 283472 315948
rect 283524 315936 283530 315988
rect 284478 315936 284484 315988
rect 284536 315976 284542 315988
rect 285582 315976 285588 315988
rect 284536 315948 285588 315976
rect 284536 315936 284542 315948
rect 285582 315936 285588 315948
rect 285640 315936 285646 315988
rect 285950 315936 285956 315988
rect 286008 315976 286014 315988
rect 286962 315976 286968 315988
rect 286008 315948 286968 315976
rect 286008 315936 286014 315948
rect 286962 315936 286968 315948
rect 287020 315936 287026 315988
rect 287146 315936 287152 315988
rect 287204 315976 287210 315988
rect 287790 315976 287796 315988
rect 287204 315948 287796 315976
rect 287204 315936 287210 315948
rect 287790 315936 287796 315948
rect 287848 315936 287854 315988
rect 288802 315936 288808 315988
rect 288860 315976 288866 315988
rect 289354 315976 289360 315988
rect 288860 315948 289360 315976
rect 288860 315936 288866 315948
rect 289354 315936 289360 315948
rect 289412 315936 289418 315988
rect 291378 315936 291384 315988
rect 291436 315976 291442 315988
rect 292390 315976 292396 315988
rect 291436 315948 292396 315976
rect 291436 315936 291442 315948
rect 292390 315936 292396 315948
rect 292448 315936 292454 315988
rect 292850 315936 292856 315988
rect 292908 315976 292914 315988
rect 293494 315976 293500 315988
rect 292908 315948 293500 315976
rect 292908 315936 292914 315948
rect 293494 315936 293500 315948
rect 293552 315936 293558 315988
rect 294506 315936 294512 315988
rect 294564 315976 294570 315988
rect 295150 315976 295156 315988
rect 294564 315948 295156 315976
rect 294564 315936 294570 315948
rect 295150 315936 295156 315948
rect 295208 315936 295214 315988
rect 295518 315936 295524 315988
rect 295576 315976 295582 315988
rect 296162 315976 296168 315988
rect 295576 315948 296168 315976
rect 295576 315936 295582 315948
rect 296162 315936 296168 315948
rect 296220 315936 296226 315988
rect 296806 315936 296812 315988
rect 296864 315976 296870 315988
rect 297542 315976 297548 315988
rect 296864 315948 297548 315976
rect 296864 315936 296870 315948
rect 297542 315936 297548 315948
rect 297600 315936 297606 315988
rect 299842 315936 299848 315988
rect 299900 315976 299906 315988
rect 300394 315976 300400 315988
rect 299900 315948 300400 315976
rect 299900 315936 299906 315948
rect 300394 315936 300400 315948
rect 300452 315936 300458 315988
rect 302510 315936 302516 315988
rect 302568 315976 302574 315988
rect 302878 315976 302884 315988
rect 302568 315948 302884 315976
rect 302568 315936 302574 315948
rect 302878 315936 302884 315948
rect 302936 315936 302942 315988
rect 303982 315936 303988 315988
rect 304040 315976 304046 315988
rect 304350 315976 304356 315988
rect 304040 315948 304356 315976
rect 304040 315936 304046 315948
rect 304350 315936 304356 315948
rect 304408 315936 304414 315988
rect 307110 315936 307116 315988
rect 307168 315976 307174 315988
rect 307386 315976 307392 315988
rect 307168 315948 307392 315976
rect 307168 315936 307174 315948
rect 307386 315936 307392 315948
rect 307444 315936 307450 315988
rect 308582 315936 308588 315988
rect 308640 315976 308646 315988
rect 308858 315976 308864 315988
rect 308640 315948 308864 315976
rect 308640 315936 308646 315948
rect 308858 315936 308864 315948
rect 308916 315936 308922 315988
rect 309410 315936 309416 315988
rect 309468 315976 309474 315988
rect 310422 315976 310428 315988
rect 309468 315948 310428 315976
rect 309468 315936 309474 315948
rect 310422 315936 310428 315948
rect 310480 315936 310486 315988
rect 310790 315936 310796 315988
rect 310848 315976 310854 315988
rect 311066 315976 311072 315988
rect 310848 315948 311072 315976
rect 310848 315936 310854 315948
rect 311066 315936 311072 315948
rect 311124 315936 311130 315988
rect 312170 315936 312176 315988
rect 312228 315976 312234 315988
rect 312814 315976 312820 315988
rect 312228 315948 312820 315976
rect 312228 315936 312234 315948
rect 312814 315936 312820 315948
rect 312872 315936 312878 315988
rect 314930 315936 314936 315988
rect 314988 315976 314994 315988
rect 315942 315976 315948 315988
rect 314988 315948 315948 315976
rect 314988 315936 314994 315948
rect 315942 315936 315948 315948
rect 316000 315936 316006 315988
rect 316310 315936 316316 315988
rect 316368 315976 316374 315988
rect 316770 315976 316776 315988
rect 316368 315948 316776 315976
rect 316368 315936 316374 315948
rect 316770 315936 316776 315948
rect 316828 315936 316834 315988
rect 317690 315936 317696 315988
rect 317748 315976 317754 315988
rect 318426 315976 318432 315988
rect 317748 315948 318432 315976
rect 317748 315936 317754 315948
rect 318426 315936 318432 315948
rect 318484 315936 318490 315988
rect 320450 315936 320456 315988
rect 320508 315976 320514 315988
rect 321370 315976 321376 315988
rect 320508 315948 321376 315976
rect 320508 315936 320514 315948
rect 321370 315936 321376 315948
rect 321428 315936 321434 315988
rect 323026 315936 323032 315988
rect 323084 315976 323090 315988
rect 323394 315976 323400 315988
rect 323084 315948 323400 315976
rect 323084 315936 323090 315948
rect 323394 315936 323400 315948
rect 323452 315936 323458 315988
rect 324406 315936 324412 315988
rect 324464 315976 324470 315988
rect 324774 315976 324780 315988
rect 324464 315948 324780 315976
rect 324464 315936 324470 315948
rect 324774 315936 324780 315948
rect 324832 315936 324838 315988
rect 288526 315868 288532 315920
rect 288584 315908 288590 315920
rect 288894 315908 288900 315920
rect 288584 315880 288900 315908
rect 288584 315868 288590 315880
rect 288894 315868 288900 315880
rect 288952 315868 288958 315920
rect 288986 315868 288992 315920
rect 289044 315908 289050 315920
rect 289630 315908 289636 315920
rect 289044 315880 289636 315908
rect 289044 315868 289050 315880
rect 289630 315868 289636 315880
rect 289688 315868 289694 315920
rect 299658 315868 299664 315920
rect 299716 315908 299722 315920
rect 300762 315908 300768 315920
rect 299716 315880 300768 315908
rect 299716 315868 299722 315880
rect 300762 315868 300768 315880
rect 300820 315868 300826 315920
rect 303798 315868 303804 315920
rect 303856 315908 303862 315920
rect 304902 315908 304908 315920
rect 303856 315880 304908 315908
rect 303856 315868 303862 315880
rect 304902 315868 304908 315880
rect 304960 315868 304966 315920
rect 309594 315868 309600 315920
rect 309652 315908 309658 315920
rect 310330 315908 310336 315920
rect 309652 315880 310336 315908
rect 309652 315868 309658 315880
rect 310330 315868 310336 315880
rect 310388 315868 310394 315920
rect 310606 315868 310612 315920
rect 310664 315908 310670 315920
rect 311710 315908 311716 315920
rect 310664 315880 311716 315908
rect 310664 315868 310670 315880
rect 311710 315868 311716 315880
rect 311768 315868 311774 315920
rect 312354 315868 312360 315920
rect 312412 315908 312418 315920
rect 313090 315908 313096 315920
rect 312412 315880 313096 315908
rect 312412 315868 312418 315880
rect 313090 315868 313096 315880
rect 313148 315868 313154 315920
rect 314746 315868 314752 315920
rect 314804 315908 314810 315920
rect 315574 315908 315580 315920
rect 314804 315880 315580 315908
rect 314804 315868 314810 315880
rect 315574 315868 315580 315880
rect 315632 315868 315638 315920
rect 318058 315868 318064 315920
rect 318116 315908 318122 315920
rect 318518 315908 318524 315920
rect 318116 315880 318524 315908
rect 318116 315868 318122 315880
rect 318518 315868 318524 315880
rect 318576 315868 318582 315920
rect 324130 315868 324136 315920
rect 324188 315908 324194 315920
rect 328638 315908 328644 315920
rect 324188 315880 328644 315908
rect 324188 315868 324194 315880
rect 328638 315868 328644 315880
rect 328696 315868 328702 315920
rect 285398 315800 285404 315852
rect 285456 315840 285462 315852
rect 285582 315840 285588 315852
rect 285456 315812 285588 315840
rect 285456 315800 285462 315812
rect 285582 315800 285588 315812
rect 285640 315800 285646 315852
rect 287238 315800 287244 315852
rect 287296 315840 287302 315852
rect 288250 315840 288256 315852
rect 287296 315812 288256 315840
rect 287296 315800 287302 315812
rect 288250 315800 288256 315812
rect 288308 315800 288314 315852
rect 288618 315800 288624 315852
rect 288676 315840 288682 315852
rect 289354 315840 289360 315852
rect 288676 315812 289360 315840
rect 288676 315800 288682 315812
rect 289354 315800 289360 315812
rect 289412 315800 289418 315852
rect 310514 315840 310520 315852
rect 292546 315812 310520 315840
rect 278222 315664 278228 315716
rect 278280 315704 278286 315716
rect 292546 315704 292574 315812
rect 310514 315800 310520 315812
rect 310572 315800 310578 315852
rect 310790 315800 310796 315852
rect 310848 315840 310854 315852
rect 311802 315840 311808 315852
rect 310848 315812 311808 315840
rect 310848 315800 310854 315812
rect 311802 315800 311808 315812
rect 311860 315800 311866 315852
rect 312078 315800 312084 315852
rect 312136 315840 312142 315852
rect 312538 315840 312544 315852
rect 312136 315812 312544 315840
rect 312136 315800 312142 315812
rect 312538 315800 312544 315812
rect 312596 315800 312602 315852
rect 319806 315840 319812 315852
rect 315684 315812 319812 315840
rect 296806 315732 296812 315784
rect 296864 315772 296870 315784
rect 297726 315772 297732 315784
rect 296864 315744 297732 315772
rect 296864 315732 296870 315744
rect 297726 315732 297732 315744
rect 297784 315732 297790 315784
rect 302418 315732 302424 315784
rect 302476 315772 302482 315784
rect 302970 315772 302976 315784
rect 302476 315744 302976 315772
rect 302476 315732 302482 315744
rect 302970 315732 302976 315744
rect 303028 315732 303034 315784
rect 309134 315732 309140 315784
rect 309192 315772 309198 315784
rect 310238 315772 310244 315784
rect 309192 315744 310244 315772
rect 309192 315732 309198 315744
rect 310238 315732 310244 315744
rect 310296 315732 310302 315784
rect 315684 315772 315712 315812
rect 319806 315800 319812 315812
rect 319864 315840 319870 315852
rect 328178 315840 328184 315852
rect 319864 315812 328184 315840
rect 319864 315800 319870 315812
rect 328178 315800 328184 315812
rect 328236 315800 328242 315852
rect 311866 315744 315712 315772
rect 278280 315676 292574 315704
rect 278280 315664 278286 315676
rect 302326 315664 302332 315716
rect 302384 315704 302390 315716
rect 303062 315704 303068 315716
rect 302384 315676 303068 315704
rect 302384 315664 302390 315676
rect 303062 315664 303068 315676
rect 303120 315664 303126 315716
rect 281350 315596 281356 315648
rect 281408 315636 281414 315648
rect 311866 315636 311894 315744
rect 315758 315732 315764 315784
rect 315816 315772 315822 315784
rect 375650 315772 375656 315784
rect 315816 315744 375656 315772
rect 315816 315732 315822 315744
rect 375650 315732 375656 315744
rect 375708 315732 375714 315784
rect 314378 315664 314384 315716
rect 314436 315704 314442 315716
rect 375006 315704 375012 315716
rect 314436 315676 375012 315704
rect 314436 315664 314442 315676
rect 375006 315664 375012 315676
rect 375064 315664 375070 315716
rect 319714 315636 319720 315648
rect 281408 315608 311894 315636
rect 316328 315608 319720 315636
rect 281408 315596 281414 315608
rect 281258 315528 281264 315580
rect 281316 315568 281322 315580
rect 316328 315568 316356 315608
rect 319714 315596 319720 315608
rect 319772 315636 319778 315648
rect 319772 315608 321554 315636
rect 319772 315596 319778 315608
rect 281316 315540 316356 315568
rect 281316 315528 281322 315540
rect 316402 315528 316408 315580
rect 316460 315568 316466 315580
rect 317322 315568 317328 315580
rect 316460 315540 317328 315568
rect 316460 315528 316466 315540
rect 317322 315528 317328 315540
rect 317380 315528 317386 315580
rect 321526 315568 321554 315608
rect 337746 315568 337752 315580
rect 321526 315540 337752 315568
rect 337746 315528 337752 315540
rect 337804 315528 337810 315580
rect 213638 315460 213644 315512
rect 213696 315500 213702 315512
rect 272610 315500 272616 315512
rect 213696 315472 272616 315500
rect 213696 315460 213702 315472
rect 272610 315460 272616 315472
rect 272668 315460 272674 315512
rect 275554 315460 275560 315512
rect 275612 315500 275618 315512
rect 320726 315500 320732 315512
rect 275612 315472 320732 315500
rect 275612 315460 275618 315472
rect 320726 315460 320732 315472
rect 320784 315460 320790 315512
rect 246942 315392 246948 315444
rect 247000 315432 247006 315444
rect 302234 315432 302240 315444
rect 247000 315404 302240 315432
rect 247000 315392 247006 315404
rect 302234 315392 302240 315404
rect 302292 315392 302298 315444
rect 302510 315392 302516 315444
rect 302568 315432 302574 315444
rect 303522 315432 303528 315444
rect 302568 315404 303528 315432
rect 302568 315392 302574 315404
rect 303522 315392 303528 315404
rect 303580 315392 303586 315444
rect 307018 315392 307024 315444
rect 307076 315432 307082 315444
rect 307478 315432 307484 315444
rect 307076 315404 307484 315432
rect 307076 315392 307082 315404
rect 307478 315392 307484 315404
rect 307536 315392 307542 315444
rect 312446 315432 312452 315444
rect 311866 315404 312452 315432
rect 213454 315324 213460 315376
rect 213512 315364 213518 315376
rect 283834 315364 283840 315376
rect 213512 315336 283840 315364
rect 213512 315324 213518 315336
rect 283834 315324 283840 315336
rect 283892 315324 283898 315376
rect 285122 315324 285128 315376
rect 285180 315364 285186 315376
rect 311866 315364 311894 315404
rect 312446 315392 312452 315404
rect 312504 315432 312510 315444
rect 336550 315432 336556 315444
rect 312504 315404 336556 315432
rect 312504 315392 312510 315404
rect 336550 315392 336556 315404
rect 336608 315392 336614 315444
rect 285180 315336 311894 315364
rect 285180 315324 285186 315336
rect 321002 315324 321008 315376
rect 321060 315364 321066 315376
rect 331582 315364 331588 315376
rect 321060 315336 331588 315364
rect 321060 315324 321066 315336
rect 331582 315324 331588 315336
rect 331640 315364 331646 315376
rect 334986 315364 334992 315376
rect 331640 315336 334992 315364
rect 331640 315324 331646 315336
rect 334986 315324 334992 315336
rect 335044 315324 335050 315376
rect 219710 315256 219716 315308
rect 219768 315296 219774 315308
rect 313642 315296 313648 315308
rect 219768 315268 313648 315296
rect 219768 315256 219774 315268
rect 313642 315256 313648 315268
rect 313700 315256 313706 315308
rect 328454 315256 328460 315308
rect 328512 315296 328518 315308
rect 328822 315296 328828 315308
rect 328512 315268 328828 315296
rect 328512 315256 328518 315268
rect 328822 315256 328828 315268
rect 328880 315296 328886 315308
rect 385034 315296 385040 315308
rect 328880 315268 385040 315296
rect 328880 315256 328886 315268
rect 385034 315256 385040 315268
rect 385092 315256 385098 315308
rect 291930 315188 291936 315240
rect 291988 315228 291994 315240
rect 317506 315228 317512 315240
rect 291988 315200 317512 315228
rect 291988 315188 291994 315200
rect 317506 315188 317512 315200
rect 317564 315188 317570 315240
rect 291654 315120 291660 315172
rect 291712 315160 291718 315172
rect 292206 315160 292212 315172
rect 291712 315132 292212 315160
rect 291712 315120 291718 315132
rect 292206 315120 292212 315132
rect 292264 315120 292270 315172
rect 308766 315120 308772 315172
rect 308824 315160 308830 315172
rect 327718 315160 327724 315172
rect 308824 315132 327724 315160
rect 308824 315120 308830 315132
rect 327718 315120 327724 315132
rect 327776 315120 327782 315172
rect 327810 315120 327816 315172
rect 327868 315160 327874 315172
rect 328638 315160 328644 315172
rect 327868 315132 328644 315160
rect 327868 315120 327874 315132
rect 328638 315120 328644 315132
rect 328696 315160 328702 315172
rect 337838 315160 337844 315172
rect 328696 315132 337844 315160
rect 328696 315120 328702 315132
rect 337838 315120 337844 315132
rect 337896 315120 337902 315172
rect 314562 315052 314568 315104
rect 314620 315092 314626 315104
rect 382734 315092 382740 315104
rect 314620 315064 382740 315092
rect 314620 315052 314626 315064
rect 382734 315052 382740 315064
rect 382792 315052 382798 315104
rect 317230 314984 317236 315036
rect 317288 315024 317294 315036
rect 377122 315024 377128 315036
rect 317288 314996 377128 315024
rect 317288 314984 317294 314996
rect 377122 314984 377128 314996
rect 377180 314984 377186 315036
rect 313182 314916 313188 314968
rect 313240 314956 313246 314968
rect 372890 314956 372896 314968
rect 313240 314928 372896 314956
rect 313240 314916 313246 314928
rect 372890 314916 372896 314928
rect 372948 314916 372954 314968
rect 287330 314848 287336 314900
rect 287388 314888 287394 314900
rect 288158 314888 288164 314900
rect 287388 314860 288164 314888
rect 287388 314848 287394 314860
rect 288158 314848 288164 314860
rect 288216 314848 288222 314900
rect 292942 314848 292948 314900
rect 293000 314888 293006 314900
rect 293586 314888 293592 314900
rect 293000 314860 293592 314888
rect 293000 314848 293006 314860
rect 293586 314848 293592 314860
rect 293644 314848 293650 314900
rect 317506 314848 317512 314900
rect 317564 314888 317570 314900
rect 332410 314888 332416 314900
rect 317564 314860 332416 314888
rect 317564 314848 317570 314860
rect 332410 314848 332416 314860
rect 332468 314848 332474 314900
rect 317322 314780 317328 314832
rect 317380 314820 317386 314832
rect 352650 314820 352656 314832
rect 317380 314792 352656 314820
rect 317380 314780 317386 314792
rect 352650 314780 352656 314792
rect 352708 314780 352714 314832
rect 302234 314712 302240 314764
rect 302292 314752 302298 314764
rect 306466 314752 306472 314764
rect 302292 314724 306472 314752
rect 302292 314712 302298 314724
rect 306466 314712 306472 314724
rect 306524 314752 306530 314764
rect 328730 314752 328736 314764
rect 306524 314724 328736 314752
rect 306524 314712 306530 314724
rect 328730 314712 328736 314724
rect 328788 314712 328794 314764
rect 248138 314644 248144 314696
rect 248196 314684 248202 314696
rect 307018 314684 307024 314696
rect 248196 314656 307024 314684
rect 248196 314644 248202 314656
rect 307018 314644 307024 314656
rect 307076 314644 307082 314696
rect 327810 314644 327816 314696
rect 327868 314684 327874 314696
rect 328270 314684 328276 314696
rect 327868 314656 328276 314684
rect 327868 314644 327874 314656
rect 328270 314644 328276 314656
rect 328328 314644 328334 314696
rect 274542 314576 274548 314628
rect 274600 314616 274606 314628
rect 306374 314616 306380 314628
rect 274600 314588 306380 314616
rect 274600 314576 274606 314588
rect 306374 314576 306380 314588
rect 306432 314576 306438 314628
rect 308398 314576 308404 314628
rect 308456 314616 308462 314628
rect 329282 314616 329288 314628
rect 308456 314588 329288 314616
rect 308456 314576 308462 314588
rect 329282 314576 329288 314588
rect 329340 314576 329346 314628
rect 275922 314508 275928 314560
rect 275980 314548 275986 314560
rect 304994 314548 305000 314560
rect 275980 314520 305000 314548
rect 275980 314508 275986 314520
rect 304994 314508 305000 314520
rect 305052 314508 305058 314560
rect 317874 314508 317880 314560
rect 317932 314548 317938 314560
rect 318426 314548 318432 314560
rect 317932 314520 318432 314548
rect 317932 314508 317938 314520
rect 318426 314508 318432 314520
rect 318484 314508 318490 314560
rect 333606 314548 333612 314560
rect 318536 314520 333612 314548
rect 284294 314440 284300 314492
rect 284352 314480 284358 314492
rect 285214 314480 285220 314492
rect 284352 314452 285220 314480
rect 284352 314440 284358 314452
rect 285214 314440 285220 314452
rect 285272 314440 285278 314492
rect 297634 314440 297640 314492
rect 297692 314480 297698 314492
rect 298002 314480 298008 314492
rect 297692 314452 298008 314480
rect 297692 314440 297698 314452
rect 298002 314440 298008 314452
rect 298060 314440 298066 314492
rect 311986 314440 311992 314492
rect 312044 314480 312050 314492
rect 318536 314480 318564 314520
rect 333606 314508 333612 314520
rect 333664 314508 333670 314560
rect 312044 314452 318564 314480
rect 312044 314440 312050 314452
rect 318610 314440 318616 314492
rect 318668 314480 318674 314492
rect 379146 314480 379152 314492
rect 318668 314452 379152 314480
rect 318668 314440 318674 314452
rect 379146 314440 379152 314452
rect 379204 314440 379210 314492
rect 296254 314372 296260 314424
rect 296312 314412 296318 314424
rect 356146 314412 356152 314424
rect 296312 314384 356152 314412
rect 296312 314372 296318 314384
rect 356146 314372 356152 314384
rect 356204 314372 356210 314424
rect 299474 314304 299480 314356
rect 299532 314344 299538 314356
rect 300854 314344 300860 314356
rect 299532 314316 300860 314344
rect 299532 314304 299538 314316
rect 300854 314304 300860 314316
rect 300912 314344 300918 314356
rect 360654 314344 360660 314356
rect 300912 314316 360660 314344
rect 300912 314304 300918 314316
rect 360654 314304 360660 314316
rect 360712 314304 360718 314356
rect 270218 314236 270224 314288
rect 270276 314276 270282 314288
rect 300302 314276 300308 314288
rect 270276 314248 300308 314276
rect 270276 314236 270282 314248
rect 300302 314236 300308 314248
rect 300360 314236 300366 314288
rect 318426 314236 318432 314288
rect 318484 314276 318490 314288
rect 376938 314276 376944 314288
rect 318484 314248 376944 314276
rect 318484 314236 318490 314248
rect 376938 314236 376944 314248
rect 376996 314236 377002 314288
rect 260466 314168 260472 314220
rect 260524 314208 260530 314220
rect 260650 314208 260656 314220
rect 260524 314180 260656 314208
rect 260524 314168 260530 314180
rect 260650 314168 260656 314180
rect 260708 314168 260714 314220
rect 297634 314168 297640 314220
rect 297692 314208 297698 314220
rect 341886 314208 341892 314220
rect 297692 314180 341892 314208
rect 297692 314168 297698 314180
rect 341886 314168 341892 314180
rect 341944 314168 341950 314220
rect 298002 314100 298008 314152
rect 298060 314140 298066 314152
rect 300578 314140 300584 314152
rect 298060 314112 300584 314140
rect 298060 314100 298066 314112
rect 300578 314100 300584 314112
rect 300636 314140 300642 314152
rect 332318 314140 332324 314152
rect 300636 314112 332324 314140
rect 300636 314100 300642 314112
rect 332318 314100 332324 314112
rect 332376 314100 332382 314152
rect 222194 314032 222200 314084
rect 222252 314072 222258 314084
rect 242434 314072 242440 314084
rect 222252 314044 242440 314072
rect 222252 314032 222258 314044
rect 242434 314032 242440 314044
rect 242492 314032 242498 314084
rect 248046 314032 248052 314084
rect 248104 314072 248110 314084
rect 308490 314072 308496 314084
rect 248104 314044 308496 314072
rect 248104 314032 248110 314044
rect 308490 314032 308496 314044
rect 308548 314032 308554 314084
rect 311250 314032 311256 314084
rect 311308 314072 311314 314084
rect 341426 314072 341432 314084
rect 311308 314044 341432 314072
rect 311308 314032 311314 314044
rect 341426 314032 341432 314044
rect 341484 314032 341490 314084
rect 210970 313964 210976 314016
rect 211028 314004 211034 314016
rect 271414 314004 271420 314016
rect 211028 313976 271420 314004
rect 211028 313964 211034 313976
rect 271414 313964 271420 313976
rect 271472 313964 271478 314016
rect 321094 314004 321100 314016
rect 311866 313976 321100 314004
rect 211890 313896 211896 313948
rect 211948 313936 211954 313948
rect 273714 313936 273720 313948
rect 211948 313908 273720 313936
rect 211948 313896 211954 313908
rect 273714 313896 273720 313908
rect 273772 313936 273778 313948
rect 274542 313936 274548 313948
rect 273772 313908 274548 313936
rect 273772 313896 273778 313908
rect 274542 313896 274548 313908
rect 274600 313896 274606 313948
rect 282454 313896 282460 313948
rect 282512 313936 282518 313948
rect 311866 313936 311894 313976
rect 321094 313964 321100 313976
rect 321152 314004 321158 314016
rect 321152 313976 321554 314004
rect 321152 313964 321158 313976
rect 282512 313908 311894 313936
rect 321526 313936 321554 313976
rect 330018 313964 330024 314016
rect 330076 314004 330082 314016
rect 390830 314004 390836 314016
rect 330076 313976 390836 314004
rect 330076 313964 330082 313976
rect 390830 313964 390836 313976
rect 390888 313964 390894 314016
rect 336274 313936 336280 313948
rect 321526 313908 336280 313936
rect 282512 313896 282518 313908
rect 336274 313896 336280 313908
rect 336332 313896 336338 313948
rect 379238 313896 379244 313948
rect 379296 313936 379302 313948
rect 466454 313936 466460 313948
rect 379296 313908 466460 313936
rect 379296 313896 379302 313908
rect 466454 313896 466460 313908
rect 466512 313896 466518 313948
rect 310514 313828 310520 313880
rect 310572 313868 310578 313880
rect 311342 313868 311348 313880
rect 310572 313840 311348 313868
rect 310572 313828 310578 313840
rect 311342 313828 311348 313840
rect 311400 313868 311406 313880
rect 329834 313868 329840 313880
rect 311400 313840 329840 313868
rect 311400 313828 311406 313840
rect 329834 313828 329840 313840
rect 329892 313828 329898 313880
rect 317874 313760 317880 313812
rect 317932 313800 317938 313812
rect 318702 313800 318708 313812
rect 317932 313772 318708 313800
rect 317932 313760 317938 313772
rect 318702 313760 318708 313772
rect 318760 313800 318766 313812
rect 379238 313800 379244 313812
rect 318760 313772 379244 313800
rect 318760 313760 318766 313772
rect 379238 313760 379244 313772
rect 379296 313760 379302 313812
rect 319438 313692 319444 313744
rect 319496 313732 319502 313744
rect 319806 313732 319812 313744
rect 319496 313704 319812 313732
rect 319496 313692 319502 313704
rect 319806 313692 319812 313704
rect 319864 313732 319870 313744
rect 379698 313732 379704 313744
rect 319864 313704 379704 313732
rect 319864 313692 319870 313704
rect 379698 313692 379704 313704
rect 379756 313692 379762 313744
rect 298738 313624 298744 313676
rect 298796 313664 298802 313676
rect 330662 313664 330668 313676
rect 298796 313636 330668 313664
rect 298796 313624 298802 313636
rect 330662 313624 330668 313636
rect 330720 313624 330726 313676
rect 279786 313556 279792 313608
rect 279844 313596 279850 313608
rect 284294 313596 284300 313608
rect 279844 313568 284300 313596
rect 279844 313556 279850 313568
rect 284294 313556 284300 313568
rect 284352 313556 284358 313608
rect 279418 313420 279424 313472
rect 279476 313460 279482 313472
rect 286042 313460 286048 313472
rect 279476 313432 286048 313460
rect 279476 313420 279482 313432
rect 286042 313420 286048 313432
rect 286100 313420 286106 313472
rect 292666 313420 292672 313472
rect 292724 313460 292730 313472
rect 293402 313460 293408 313472
rect 292724 313432 293408 313460
rect 292724 313420 292730 313432
rect 293402 313420 293408 313432
rect 293460 313420 293466 313472
rect 275738 313352 275744 313404
rect 275796 313392 275802 313404
rect 287698 313392 287704 313404
rect 275796 313364 287704 313392
rect 275796 313352 275802 313364
rect 287698 313352 287704 313364
rect 287756 313352 287762 313404
rect 270218 313284 270224 313336
rect 270276 313324 270282 313336
rect 270678 313324 270684 313336
rect 270276 313296 270684 313324
rect 270276 313284 270282 313296
rect 270678 313284 270684 313296
rect 270736 313284 270742 313336
rect 272610 313284 272616 313336
rect 272668 313324 272674 313336
rect 312446 313324 312452 313336
rect 272668 313296 312452 313324
rect 272668 313284 272674 313296
rect 312446 313284 312452 313296
rect 312504 313284 312510 313336
rect 260558 313216 260564 313268
rect 260616 313256 260622 313268
rect 260742 313256 260748 313268
rect 260616 313228 260748 313256
rect 260616 313216 260622 313228
rect 260742 313216 260748 313228
rect 260800 313256 260806 313268
rect 287054 313256 287060 313268
rect 260800 313228 287060 313256
rect 260800 313216 260806 313228
rect 287054 313216 287060 313228
rect 287112 313216 287118 313268
rect 309870 313216 309876 313268
rect 309928 313256 309934 313268
rect 310422 313256 310428 313268
rect 309928 313228 310428 313256
rect 309928 313216 309934 313228
rect 310422 313216 310428 313228
rect 310480 313216 310486 313268
rect 322106 313216 322112 313268
rect 322164 313256 322170 313268
rect 389266 313256 389272 313268
rect 322164 313228 389272 313256
rect 322164 313216 322170 313228
rect 389266 313216 389272 313228
rect 389324 313216 389330 313268
rect 523678 313216 523684 313268
rect 523736 313256 523742 313268
rect 579614 313256 579620 313268
rect 523736 313228 579620 313256
rect 523736 313216 523742 313228
rect 579614 313216 579620 313228
rect 579672 313216 579678 313268
rect 305638 313148 305644 313200
rect 305696 313188 305702 313200
rect 330570 313188 330576 313200
rect 305696 313160 330576 313188
rect 305696 313148 305702 313160
rect 330570 313148 330576 313160
rect 330628 313148 330634 313200
rect 313090 313080 313096 313132
rect 313148 313120 313154 313132
rect 372798 313120 372804 313132
rect 313148 313092 372804 313120
rect 313148 313080 313154 313092
rect 372798 313080 372804 313092
rect 372856 313080 372862 313132
rect 309686 313012 309692 313064
rect 309744 313052 309750 313064
rect 310054 313052 310060 313064
rect 309744 313024 310060 313052
rect 309744 313012 309750 313024
rect 310054 313012 310060 313024
rect 310112 313052 310118 313064
rect 329926 313052 329932 313064
rect 310112 313024 329932 313052
rect 310112 313012 310118 313024
rect 329926 313012 329932 313024
rect 329984 313012 329990 313064
rect 294874 312944 294880 312996
rect 294932 312984 294938 312996
rect 341794 312984 341800 312996
rect 294932 312956 341800 312984
rect 294932 312944 294938 312956
rect 341794 312944 341800 312956
rect 341852 312944 341858 312996
rect 295426 312876 295432 312928
rect 295484 312916 295490 312928
rect 331030 312916 331036 312928
rect 295484 312888 331036 312916
rect 295484 312876 295490 312888
rect 331030 312876 331036 312888
rect 331088 312876 331094 312928
rect 315206 312808 315212 312860
rect 315264 312848 315270 312860
rect 350166 312848 350172 312860
rect 315264 312820 350172 312848
rect 315264 312808 315270 312820
rect 350166 312808 350172 312820
rect 350224 312808 350230 312860
rect 202690 312740 202696 312792
rect 202748 312780 202754 312792
rect 260742 312780 260748 312792
rect 202748 312752 260748 312780
rect 202748 312740 202754 312752
rect 260742 312740 260748 312752
rect 260800 312740 260806 312792
rect 322842 312780 322848 312792
rect 316696 312752 322848 312780
rect 253658 312672 253664 312724
rect 253716 312712 253722 312724
rect 313090 312712 313096 312724
rect 253716 312684 313096 312712
rect 253716 312672 253722 312684
rect 313090 312672 313096 312684
rect 313148 312672 313154 312724
rect 252462 312604 252468 312656
rect 252520 312644 252526 312656
rect 312814 312644 312820 312656
rect 252520 312616 312820 312644
rect 252520 312604 252526 312616
rect 312814 312604 312820 312616
rect 312872 312604 312878 312656
rect 210602 312536 210608 312588
rect 210660 312576 210666 312588
rect 278406 312576 278412 312588
rect 210660 312548 278412 312576
rect 210660 312536 210666 312548
rect 278406 312536 278412 312548
rect 278464 312536 278470 312588
rect 278682 312536 278688 312588
rect 278740 312576 278746 312588
rect 316696 312576 316724 312752
rect 322842 312740 322848 312752
rect 322900 312740 322906 312792
rect 329834 312740 329840 312792
rect 329892 312780 329898 312792
rect 330938 312780 330944 312792
rect 329892 312752 330944 312780
rect 329892 312740 329898 312752
rect 330938 312740 330944 312752
rect 330996 312740 331002 312792
rect 343358 312780 343364 312792
rect 331186 312752 343364 312780
rect 317138 312672 317144 312724
rect 317196 312712 317202 312724
rect 331186 312712 331214 312752
rect 343358 312740 343364 312752
rect 343416 312740 343422 312792
rect 317196 312684 331214 312712
rect 317196 312672 317202 312684
rect 328362 312604 328368 312656
rect 328420 312644 328426 312656
rect 333146 312644 333152 312656
rect 328420 312616 333152 312644
rect 328420 312604 328426 312616
rect 333146 312604 333152 312616
rect 333204 312644 333210 312656
rect 387886 312644 387892 312656
rect 333204 312616 387892 312644
rect 333204 312604 333210 312616
rect 387886 312604 387892 312616
rect 387944 312604 387950 312656
rect 278740 312548 316724 312576
rect 278740 312536 278746 312548
rect 322842 312536 322848 312588
rect 322900 312576 322906 312588
rect 336182 312576 336188 312588
rect 322900 312548 336188 312576
rect 322900 312536 322906 312548
rect 336182 312536 336188 312548
rect 336240 312536 336246 312588
rect 502334 312576 502340 312588
rect 383626 312548 502340 312576
rect 301498 312468 301504 312520
rect 301556 312508 301562 312520
rect 301866 312508 301872 312520
rect 301556 312480 301872 312508
rect 301556 312468 301562 312480
rect 301866 312468 301872 312480
rect 301924 312508 301930 312520
rect 335078 312508 335084 312520
rect 301924 312480 335084 312508
rect 301924 312468 301930 312480
rect 335078 312468 335084 312480
rect 335136 312468 335142 312520
rect 304994 312400 305000 312452
rect 305052 312440 305058 312452
rect 305638 312440 305644 312452
rect 305052 312412 305644 312440
rect 305052 312400 305058 312412
rect 305638 312400 305644 312412
rect 305696 312400 305702 312452
rect 321002 312400 321008 312452
rect 321060 312440 321066 312452
rect 321278 312440 321284 312452
rect 321060 312412 321284 312440
rect 321060 312400 321066 312412
rect 321278 312400 321284 312412
rect 321336 312440 321342 312452
rect 381354 312440 381360 312452
rect 321336 312412 381360 312440
rect 321336 312400 321342 312412
rect 381354 312400 381360 312412
rect 381412 312440 381418 312452
rect 383626 312440 383654 312548
rect 502334 312536 502340 312548
rect 502392 312536 502398 312588
rect 381412 312412 383654 312440
rect 381412 312400 381418 312412
rect 277854 312332 277860 312384
rect 277912 312372 277918 312384
rect 322106 312372 322112 312384
rect 277912 312344 322112 312372
rect 277912 312332 277918 312344
rect 322106 312332 322112 312344
rect 322164 312332 322170 312384
rect 322750 312332 322756 312384
rect 322808 312372 322814 312384
rect 371878 312372 371884 312384
rect 322808 312344 371884 312372
rect 322808 312332 322814 312344
rect 371878 312332 371884 312344
rect 371936 312332 371942 312384
rect 336366 312304 336372 312316
rect 311866 312276 336372 312304
rect 310422 312196 310428 312248
rect 310480 312236 310486 312248
rect 311866 312236 311894 312276
rect 336366 312264 336372 312276
rect 336424 312264 336430 312316
rect 310480 312208 311894 312236
rect 310480 312196 310486 312208
rect 312814 312128 312820 312180
rect 312872 312168 312878 312180
rect 321554 312168 321560 312180
rect 312872 312140 321560 312168
rect 312872 312128 312878 312140
rect 321554 312128 321560 312140
rect 321612 312128 321618 312180
rect 262030 311788 262036 311840
rect 262088 311828 262094 311840
rect 287238 311828 287244 311840
rect 262088 311800 287244 311828
rect 262088 311788 262094 311800
rect 287238 311788 287244 311800
rect 287296 311788 287302 311840
rect 295334 311788 295340 311840
rect 295392 311828 295398 311840
rect 297910 311828 297916 311840
rect 295392 311800 297916 311828
rect 295392 311788 295398 311800
rect 297910 311788 297916 311800
rect 297968 311828 297974 311840
rect 333238 311828 333244 311840
rect 297968 311800 333244 311828
rect 297968 311788 297974 311800
rect 333238 311788 333244 311800
rect 333296 311788 333302 311840
rect 266354 311720 266360 311772
rect 266412 311760 266418 311772
rect 267550 311760 267556 311772
rect 266412 311732 267556 311760
rect 266412 311720 266418 311732
rect 267550 311720 267556 311732
rect 267608 311760 267614 311772
rect 287422 311760 287428 311772
rect 267608 311732 287428 311760
rect 267608 311720 267614 311732
rect 287422 311720 287428 311732
rect 287480 311720 287486 311772
rect 299106 311720 299112 311772
rect 299164 311760 299170 311772
rect 358078 311760 358084 311772
rect 299164 311732 358084 311760
rect 299164 311720 299170 311732
rect 358078 311720 358084 311732
rect 358136 311720 358142 311772
rect 293034 311652 293040 311704
rect 293092 311692 293098 311704
rect 293402 311692 293408 311704
rect 293092 311664 293408 311692
rect 293092 311652 293098 311664
rect 293402 311652 293408 311664
rect 293460 311692 293466 311704
rect 352374 311692 352380 311704
rect 293460 311664 352380 311692
rect 293460 311652 293466 311664
rect 352374 311652 352380 311664
rect 352432 311652 352438 311704
rect 309106 311596 313136 311624
rect 301590 311556 301596 311568
rect 296686 311528 301596 311556
rect 287790 311448 287796 311500
rect 287848 311488 287854 311500
rect 296686 311488 296714 311528
rect 301590 311516 301596 311528
rect 301648 311556 301654 311568
rect 309106 311556 309134 311596
rect 301648 311528 309134 311556
rect 313108 311556 313136 311596
rect 313734 311584 313740 311636
rect 313792 311624 313798 311636
rect 369762 311624 369768 311636
rect 313792 311596 369768 311624
rect 313792 311584 313798 311596
rect 369762 311584 369768 311596
rect 369820 311624 369826 311636
rect 374086 311624 374092 311636
rect 369820 311596 374092 311624
rect 369820 311584 369826 311596
rect 374086 311584 374092 311596
rect 374144 311584 374150 311636
rect 355594 311556 355600 311568
rect 313108 311528 355600 311556
rect 301648 311516 301654 311528
rect 355594 311516 355600 311528
rect 355652 311516 355658 311568
rect 287848 311460 296714 311488
rect 287848 311448 287854 311460
rect 304350 311448 304356 311500
rect 304408 311488 304414 311500
rect 306006 311488 306012 311500
rect 304408 311460 306012 311488
rect 304408 311448 304414 311460
rect 306006 311448 306012 311460
rect 306064 311448 306070 311500
rect 311526 311448 311532 311500
rect 311584 311488 311590 311500
rect 313734 311488 313740 311500
rect 311584 311460 313740 311488
rect 311584 311448 311590 311460
rect 313734 311448 313740 311460
rect 313792 311448 313798 311500
rect 321554 311448 321560 311500
rect 321612 311488 321618 311500
rect 371418 311488 371424 311500
rect 321612 311460 371424 311488
rect 321612 311448 321618 311460
rect 371418 311448 371424 311460
rect 371476 311448 371482 311500
rect 289170 311380 289176 311432
rect 289228 311420 289234 311432
rect 298002 311420 298008 311432
rect 289228 311392 298008 311420
rect 289228 311380 289234 311392
rect 298002 311380 298008 311392
rect 298060 311380 298066 311432
rect 300762 311380 300768 311432
rect 300820 311420 300826 311432
rect 346210 311420 346216 311432
rect 300820 311392 346216 311420
rect 300820 311380 300826 311392
rect 346210 311380 346216 311392
rect 346268 311380 346274 311432
rect 287974 311312 287980 311364
rect 288032 311352 288038 311364
rect 288032 311324 289216 311352
rect 288032 311312 288038 311324
rect 288894 311244 288900 311296
rect 288952 311284 288958 311296
rect 289078 311284 289084 311296
rect 288952 311256 289084 311284
rect 288952 311244 288958 311256
rect 289078 311244 289084 311256
rect 289136 311244 289142 311296
rect 289188 311284 289216 311324
rect 293218 311312 293224 311364
rect 293276 311352 293282 311364
rect 336090 311352 336096 311364
rect 293276 311324 336096 311352
rect 293276 311312 293282 311324
rect 336090 311312 336096 311324
rect 336148 311312 336154 311364
rect 299842 311284 299848 311296
rect 289188 311256 299848 311284
rect 299842 311244 299848 311256
rect 299900 311284 299906 311296
rect 300670 311284 300676 311296
rect 299900 311256 300676 311284
rect 299900 311244 299906 311256
rect 300670 311244 300676 311256
rect 300728 311244 300734 311296
rect 342898 311284 342904 311296
rect 300964 311256 342904 311284
rect 219158 311176 219164 311228
rect 219216 311216 219222 311228
rect 262030 311216 262036 311228
rect 219216 311188 262036 311216
rect 219216 311176 219222 311188
rect 262030 311176 262036 311188
rect 262088 311176 262094 311228
rect 282730 311176 282736 311228
rect 282788 311216 282794 311228
rect 298278 311216 298284 311228
rect 282788 311188 298284 311216
rect 282788 311176 282794 311188
rect 298278 311176 298284 311188
rect 298336 311216 298342 311228
rect 299106 311216 299112 311228
rect 298336 311188 299112 311216
rect 298336 311176 298342 311188
rect 299106 311176 299112 311188
rect 299164 311176 299170 311228
rect 299934 311176 299940 311228
rect 299992 311216 299998 311228
rect 300964 311216 300992 311256
rect 342898 311244 342904 311256
rect 342956 311244 342962 311296
rect 339126 311216 339132 311228
rect 299992 311188 300992 311216
rect 306346 311188 339132 311216
rect 299992 311176 299998 311188
rect 209406 311108 209412 311160
rect 209464 311148 209470 311160
rect 266354 311148 266360 311160
rect 209464 311120 266360 311148
rect 209464 311108 209470 311120
rect 266354 311108 266360 311120
rect 266412 311108 266418 311160
rect 285030 311108 285036 311160
rect 285088 311148 285094 311160
rect 300210 311148 300216 311160
rect 285088 311120 300216 311148
rect 285088 311108 285094 311120
rect 300210 311108 300216 311120
rect 300268 311148 300274 311160
rect 300762 311148 300768 311160
rect 300268 311120 300768 311148
rect 300268 311108 300274 311120
rect 300762 311108 300768 311120
rect 300820 311108 300826 311160
rect 300670 310972 300676 311024
rect 300728 311012 300734 311024
rect 306346 311012 306374 311188
rect 339126 311176 339132 311188
rect 339184 311176 339190 311228
rect 310882 311108 310888 311160
rect 310940 311148 310946 311160
rect 311250 311148 311256 311160
rect 310940 311120 311256 311148
rect 310940 311108 310946 311120
rect 311250 311108 311256 311120
rect 311308 311108 311314 311160
rect 315942 311108 315948 311160
rect 316000 311148 316006 311160
rect 351546 311148 351552 311160
rect 316000 311120 351552 311148
rect 316000 311108 316006 311120
rect 351546 311108 351552 311120
rect 351604 311108 351610 311160
rect 311066 311040 311072 311092
rect 311124 311080 311130 311092
rect 311802 311080 311808 311092
rect 311124 311052 311808 311080
rect 311124 311040 311130 311052
rect 311802 311040 311808 311052
rect 311860 311080 311866 311092
rect 347406 311080 347412 311092
rect 311860 311052 347412 311080
rect 311860 311040 311866 311052
rect 347406 311040 347412 311052
rect 347464 311040 347470 311092
rect 300728 310984 306374 311012
rect 300728 310972 300734 310984
rect 308306 310972 308312 311024
rect 308364 311012 308370 311024
rect 342346 311012 342352 311024
rect 308364 310984 342352 311012
rect 308364 310972 308370 310984
rect 342346 310972 342352 310984
rect 342404 310972 342410 311024
rect 311250 310904 311256 310956
rect 311308 310944 311314 310956
rect 371234 310944 371240 310956
rect 311308 310916 371240 310944
rect 311308 310904 311314 310916
rect 371234 310904 371240 310916
rect 371292 310904 371298 310956
rect 271690 310496 271696 310548
rect 271748 310536 271754 310548
rect 291102 310536 291108 310548
rect 271748 310508 291108 310536
rect 271748 310496 271754 310508
rect 291102 310496 291108 310508
rect 291160 310496 291166 310548
rect 315022 310496 315028 310548
rect 315080 310536 315086 310548
rect 315942 310536 315948 310548
rect 315080 310508 315948 310536
rect 315080 310496 315086 310508
rect 315942 310496 315948 310508
rect 316000 310496 316006 310548
rect 259362 310428 259368 310480
rect 259420 310468 259426 310480
rect 284478 310468 284484 310480
rect 259420 310440 284484 310468
rect 259420 310428 259426 310440
rect 284478 310428 284484 310440
rect 284536 310428 284542 310480
rect 299106 310428 299112 310480
rect 299164 310468 299170 310480
rect 305086 310468 305092 310480
rect 299164 310440 305092 310468
rect 299164 310428 299170 310440
rect 305086 310428 305092 310440
rect 305144 310468 305150 310480
rect 333514 310468 333520 310480
rect 305144 310440 333520 310468
rect 305144 310428 305150 310440
rect 333514 310428 333520 310440
rect 333572 310428 333578 310480
rect 283282 310360 283288 310412
rect 283340 310400 283346 310412
rect 283558 310400 283564 310412
rect 283340 310372 283564 310400
rect 283340 310360 283346 310372
rect 283558 310360 283564 310372
rect 283616 310360 283622 310412
rect 297358 310360 297364 310412
rect 297416 310400 297422 310412
rect 304994 310400 305000 310412
rect 297416 310372 305000 310400
rect 297416 310360 297422 310372
rect 304994 310360 305000 310372
rect 305052 310360 305058 310412
rect 317506 310360 317512 310412
rect 317564 310400 317570 310412
rect 317564 310372 325694 310400
rect 317564 310360 317570 310372
rect 325666 310332 325694 310372
rect 327718 310360 327724 310412
rect 327776 310400 327782 310412
rect 341702 310400 341708 310412
rect 327776 310372 341708 310400
rect 327776 310360 327782 310372
rect 341702 310360 341708 310372
rect 341760 310360 341766 310412
rect 381170 310332 381176 310344
rect 325666 310304 381176 310332
rect 381170 310292 381176 310304
rect 381228 310292 381234 310344
rect 313550 310224 313556 310276
rect 313608 310264 313614 310276
rect 374914 310264 374920 310276
rect 313608 310236 374920 310264
rect 313608 310224 313614 310236
rect 374914 310224 374920 310236
rect 374972 310224 374978 310276
rect 330386 310156 330392 310208
rect 330444 310196 330450 310208
rect 383746 310196 383752 310208
rect 330444 310168 383752 310196
rect 330444 310156 330450 310168
rect 383746 310156 383752 310168
rect 383804 310156 383810 310208
rect 297818 310088 297824 310140
rect 297876 310128 297882 310140
rect 298922 310128 298928 310140
rect 297876 310100 298928 310128
rect 297876 310088 297882 310100
rect 298922 310088 298928 310100
rect 298980 310128 298986 310140
rect 356790 310128 356796 310140
rect 298980 310100 356796 310128
rect 298980 310088 298986 310100
rect 356790 310088 356796 310100
rect 356848 310088 356854 310140
rect 286502 310020 286508 310072
rect 286560 310060 286566 310072
rect 295426 310060 295432 310072
rect 286560 310032 295432 310060
rect 286560 310020 286566 310032
rect 295426 310020 295432 310032
rect 295484 310020 295490 310072
rect 313918 310020 313924 310072
rect 313976 310060 313982 310072
rect 373258 310060 373264 310072
rect 313976 310032 373264 310060
rect 313976 310020 313982 310032
rect 373258 310020 373264 310032
rect 373316 310020 373322 310072
rect 286870 309952 286876 310004
rect 286928 309992 286934 310004
rect 297174 309992 297180 310004
rect 286928 309964 297180 309992
rect 286928 309952 286934 309964
rect 297174 309952 297180 309964
rect 297232 309992 297238 310004
rect 355318 309992 355324 310004
rect 297232 309964 355324 309992
rect 297232 309952 297238 309964
rect 355318 309952 355324 309964
rect 355376 309952 355382 310004
rect 226058 309884 226064 309936
rect 226116 309924 226122 309936
rect 259362 309924 259368 309936
rect 226116 309896 259368 309924
rect 226116 309884 226122 309896
rect 259362 309884 259368 309896
rect 259420 309884 259426 309936
rect 340506 309924 340512 309936
rect 296686 309896 340512 309924
rect 219066 309816 219072 309868
rect 219124 309856 219130 309868
rect 295702 309856 295708 309868
rect 219124 309828 295708 309856
rect 219124 309816 219130 309828
rect 295702 309816 295708 309828
rect 295760 309856 295766 309868
rect 296686 309856 296714 309896
rect 340506 309884 340512 309896
rect 340564 309884 340570 309936
rect 342346 309884 342352 309936
rect 342404 309924 342410 309936
rect 342898 309924 342904 309936
rect 342404 309896 342904 309924
rect 342404 309884 342410 309896
rect 342898 309884 342904 309896
rect 342956 309924 342962 309936
rect 369210 309924 369216 309936
rect 342956 309896 369216 309924
rect 342956 309884 342962 309896
rect 369210 309884 369216 309896
rect 369268 309884 369274 309936
rect 295760 309828 296714 309856
rect 295760 309816 295766 309828
rect 302878 309816 302884 309868
rect 302936 309856 302942 309868
rect 344830 309856 344836 309868
rect 302936 309828 344836 309856
rect 302936 309816 302942 309828
rect 344830 309816 344836 309828
rect 344888 309816 344894 309868
rect 217778 309748 217784 309800
rect 217836 309788 217842 309800
rect 294506 309788 294512 309800
rect 217836 309760 294512 309788
rect 217836 309748 217842 309760
rect 294506 309748 294512 309760
rect 294564 309788 294570 309800
rect 338942 309788 338948 309800
rect 294564 309760 338948 309788
rect 294564 309748 294570 309760
rect 338942 309748 338948 309760
rect 339000 309748 339006 309800
rect 316954 309680 316960 309732
rect 317012 309720 317018 309732
rect 354122 309720 354128 309732
rect 317012 309692 354128 309720
rect 317012 309680 317018 309692
rect 354122 309680 354128 309692
rect 354180 309680 354186 309732
rect 316218 309612 316224 309664
rect 316276 309652 316282 309664
rect 390738 309652 390744 309664
rect 316276 309624 390744 309652
rect 316276 309612 316282 309624
rect 390738 309612 390744 309624
rect 390796 309612 390802 309664
rect 310974 309544 310980 309596
rect 311032 309584 311038 309596
rect 311526 309584 311532 309596
rect 311032 309556 311532 309584
rect 311032 309544 311038 309556
rect 311526 309544 311532 309556
rect 311584 309544 311590 309596
rect 319990 309544 319996 309596
rect 320048 309584 320054 309596
rect 387794 309584 387800 309596
rect 320048 309556 387800 309584
rect 320048 309544 320054 309556
rect 387794 309544 387800 309556
rect 387852 309544 387858 309596
rect 283558 309476 283564 309528
rect 283616 309516 283622 309528
rect 327994 309516 328000 309528
rect 283616 309488 328000 309516
rect 283616 309476 283622 309488
rect 327994 309476 328000 309488
rect 328052 309476 328058 309528
rect 323670 309408 323676 309460
rect 323728 309448 323734 309460
rect 330386 309448 330392 309460
rect 323728 309420 330392 309448
rect 323728 309408 323734 309420
rect 330386 309408 330392 309420
rect 330444 309408 330450 309460
rect 275922 309204 275928 309256
rect 275980 309244 275986 309256
rect 285674 309244 285680 309256
rect 275980 309216 285680 309244
rect 275980 309204 275986 309216
rect 285674 309204 285680 309216
rect 285732 309204 285738 309256
rect 316310 309204 316316 309256
rect 316368 309244 316374 309256
rect 316954 309244 316960 309256
rect 316368 309216 316960 309244
rect 316368 309204 316374 309216
rect 316954 309204 316960 309216
rect 317012 309204 317018 309256
rect 327166 309204 327172 309256
rect 327224 309244 327230 309256
rect 327534 309244 327540 309256
rect 327224 309216 327540 309244
rect 327224 309204 327230 309216
rect 327534 309204 327540 309216
rect 327592 309204 327598 309256
rect 274542 309136 274548 309188
rect 274600 309176 274606 309188
rect 288250 309176 288256 309188
rect 274600 309148 288256 309176
rect 274600 309136 274606 309148
rect 288250 309136 288256 309148
rect 288308 309136 288314 309188
rect 302712 309148 303108 309176
rect 260466 309068 260472 309120
rect 260524 309108 260530 309120
rect 260742 309108 260748 309120
rect 260524 309080 260748 309108
rect 260524 309068 260530 309080
rect 260742 309068 260748 309080
rect 260800 309108 260806 309120
rect 285950 309108 285956 309120
rect 260800 309080 285956 309108
rect 260800 309068 260806 309080
rect 285950 309068 285956 309080
rect 286008 309068 286014 309120
rect 300302 309068 300308 309120
rect 300360 309108 300366 309120
rect 302142 309108 302148 309120
rect 300360 309080 302148 309108
rect 300360 309068 300366 309080
rect 302142 309068 302148 309080
rect 302200 309108 302206 309120
rect 302712 309108 302740 309148
rect 302200 309080 302740 309108
rect 302200 309068 302206 309080
rect 302786 309068 302792 309120
rect 302844 309108 302850 309120
rect 302970 309108 302976 309120
rect 302844 309080 302976 309108
rect 302844 309068 302850 309080
rect 302970 309068 302976 309080
rect 303028 309068 303034 309120
rect 303080 309108 303108 309148
rect 316218 309136 316224 309188
rect 316276 309176 316282 309188
rect 316678 309176 316684 309188
rect 316276 309148 316684 309176
rect 316276 309136 316282 309148
rect 316678 309136 316684 309148
rect 316736 309136 316742 309188
rect 317506 309136 317512 309188
rect 317564 309176 317570 309188
rect 318518 309176 318524 309188
rect 317564 309148 318524 309176
rect 317564 309136 317570 309148
rect 318518 309136 318524 309148
rect 318576 309136 318582 309188
rect 364610 309108 364616 309120
rect 303080 309080 364616 309108
rect 364610 309068 364616 309080
rect 364668 309068 364674 309120
rect 270402 309000 270408 309052
rect 270460 309040 270466 309052
rect 288066 309040 288072 309052
rect 270460 309012 288072 309040
rect 270460 309000 270466 309012
rect 288066 309000 288072 309012
rect 288124 309000 288130 309052
rect 302602 309000 302608 309052
rect 302660 309040 302666 309052
rect 303154 309040 303160 309052
rect 302660 309012 303160 309040
rect 302660 309000 302666 309012
rect 303154 309000 303160 309012
rect 303212 309000 303218 309052
rect 310790 309000 310796 309052
rect 310848 309040 310854 309052
rect 311342 309040 311348 309052
rect 310848 309012 311348 309040
rect 310848 309000 310854 309012
rect 311342 309000 311348 309012
rect 311400 309040 311406 309052
rect 371326 309040 371332 309052
rect 311400 309012 371332 309040
rect 311400 309000 311406 309012
rect 371326 309000 371332 309012
rect 371384 309000 371390 309052
rect 301682 308932 301688 308984
rect 301740 308972 301746 308984
rect 304166 308972 304172 308984
rect 301740 308944 304172 308972
rect 301740 308932 301746 308944
rect 304166 308932 304172 308944
rect 304224 308972 304230 308984
rect 364518 308972 364524 308984
rect 304224 308944 364524 308972
rect 304224 308932 304230 308944
rect 364518 308932 364524 308944
rect 364576 308932 364582 308984
rect 302970 308864 302976 308916
rect 303028 308904 303034 308916
rect 360930 308904 360936 308916
rect 303028 308876 360936 308904
rect 303028 308864 303034 308876
rect 360930 308864 360936 308876
rect 360988 308864 360994 308916
rect 303154 308796 303160 308848
rect 303212 308836 303218 308848
rect 359642 308836 359648 308848
rect 303212 308808 359648 308836
rect 303212 308796 303218 308808
rect 359642 308796 359648 308808
rect 359700 308796 359706 308848
rect 293954 308728 293960 308780
rect 294012 308768 294018 308780
rect 294414 308768 294420 308780
rect 294012 308740 294420 308768
rect 294012 308728 294018 308740
rect 294414 308728 294420 308740
rect 294472 308768 294478 308780
rect 350074 308768 350080 308780
rect 294472 308740 350080 308768
rect 294472 308728 294478 308740
rect 350074 308728 350080 308740
rect 350132 308728 350138 308780
rect 294046 308660 294052 308712
rect 294104 308700 294110 308712
rect 294322 308700 294328 308712
rect 294104 308672 294328 308700
rect 294104 308660 294110 308672
rect 294322 308660 294328 308672
rect 294380 308700 294386 308712
rect 348878 308700 348884 308712
rect 294380 308672 348884 308700
rect 294380 308660 294386 308672
rect 348878 308660 348884 308672
rect 348936 308660 348942 308712
rect 207934 308592 207940 308644
rect 207992 308632 207998 308644
rect 270402 308632 270408 308644
rect 207992 308604 270408 308632
rect 207992 308592 207998 308604
rect 270402 308592 270408 308604
rect 270460 308592 270466 308644
rect 304074 308592 304080 308644
rect 304132 308632 304138 308644
rect 304442 308632 304448 308644
rect 304132 308604 304448 308632
rect 304132 308592 304138 308604
rect 304442 308592 304448 308604
rect 304500 308632 304506 308644
rect 355502 308632 355508 308644
rect 304500 308604 355508 308632
rect 304500 308592 304506 308604
rect 355502 308592 355508 308604
rect 355560 308592 355566 308644
rect 219802 308524 219808 308576
rect 219860 308564 219866 308576
rect 260742 308564 260748 308576
rect 219860 308536 260748 308564
rect 219860 308524 219866 308536
rect 260742 308524 260748 308536
rect 260800 308524 260806 308576
rect 264882 308524 264888 308576
rect 264940 308564 264946 308576
rect 332962 308564 332968 308576
rect 264940 308536 332968 308564
rect 264940 308524 264946 308536
rect 332962 308524 332968 308536
rect 333020 308524 333026 308576
rect 259638 308456 259644 308508
rect 259696 308496 259702 308508
rect 332594 308496 332600 308508
rect 259696 308468 332600 308496
rect 259696 308456 259702 308468
rect 332594 308456 332600 308468
rect 332652 308456 332658 308508
rect 217410 308388 217416 308440
rect 217468 308428 217474 308440
rect 293954 308428 293960 308440
rect 217468 308400 293960 308428
rect 217468 308388 217474 308400
rect 293954 308388 293960 308400
rect 294012 308388 294018 308440
rect 300210 308388 300216 308440
rect 300268 308428 300274 308440
rect 302694 308428 302700 308440
rect 300268 308400 302700 308428
rect 300268 308388 300274 308400
rect 302694 308388 302700 308400
rect 302752 308428 302758 308440
rect 340598 308428 340604 308440
rect 302752 308400 340604 308428
rect 302752 308388 302758 308400
rect 340598 308388 340604 308400
rect 340656 308388 340662 308440
rect 371326 308388 371332 308440
rect 371384 308428 371390 308440
rect 372154 308428 372160 308440
rect 371384 308400 372160 308428
rect 371384 308388 371390 308400
rect 372154 308388 372160 308400
rect 372212 308428 372218 308440
rect 378134 308428 378140 308440
rect 372212 308400 378140 308428
rect 372212 308388 372218 308400
rect 378134 308388 378140 308400
rect 378192 308388 378198 308440
rect 305270 308320 305276 308372
rect 305328 308360 305334 308372
rect 305822 308360 305828 308372
rect 305328 308332 305828 308360
rect 305328 308320 305334 308332
rect 305822 308320 305828 308332
rect 305880 308360 305886 308372
rect 340414 308360 340420 308372
rect 305880 308332 340420 308360
rect 305880 308320 305886 308332
rect 340414 308320 340420 308332
rect 340472 308320 340478 308372
rect 292942 308252 292948 308304
rect 293000 308292 293006 308304
rect 298278 308292 298284 308304
rect 293000 308264 298284 308292
rect 293000 308252 293006 308264
rect 298278 308252 298284 308264
rect 298336 308292 298342 308304
rect 331950 308292 331956 308304
rect 298336 308264 331956 308292
rect 298336 308252 298342 308264
rect 331950 308252 331956 308264
rect 332008 308252 332014 308304
rect 319622 308184 319628 308236
rect 319680 308224 319686 308236
rect 339218 308224 339224 308236
rect 319680 308196 339224 308224
rect 319680 308184 319686 308196
rect 339218 308184 339224 308196
rect 339276 308184 339282 308236
rect 216122 307844 216128 307896
rect 216180 307884 216186 307896
rect 292942 307884 292948 307896
rect 216180 307856 292948 307884
rect 216180 307844 216186 307856
rect 292942 307844 292948 307856
rect 293000 307844 293006 307896
rect 216214 307776 216220 307828
rect 216272 307816 216278 307828
rect 293954 307816 293960 307828
rect 216272 307788 293960 307816
rect 216272 307776 216278 307788
rect 293954 307776 293960 307788
rect 294012 307776 294018 307828
rect 263134 307708 263140 307760
rect 263192 307748 263198 307760
rect 263410 307748 263416 307760
rect 263192 307720 263416 307748
rect 263192 307708 263198 307720
rect 263410 307708 263416 307720
rect 263468 307748 263474 307760
rect 283190 307748 283196 307760
rect 263468 307720 283196 307748
rect 263468 307708 263474 307720
rect 283190 307708 283196 307720
rect 283248 307708 283254 307760
rect 338666 307748 338672 307760
rect 306346 307720 338672 307748
rect 287698 307640 287704 307692
rect 287756 307680 287762 307692
rect 303982 307680 303988 307692
rect 287756 307652 303988 307680
rect 287756 307640 287762 307652
rect 303982 307640 303988 307652
rect 304040 307680 304046 307692
rect 306346 307680 306374 307720
rect 338666 307708 338672 307720
rect 338724 307708 338730 307760
rect 304040 307652 306374 307680
rect 304040 307640 304046 307652
rect 310698 307640 310704 307692
rect 310756 307680 310762 307692
rect 311434 307680 311440 307692
rect 310756 307652 311440 307680
rect 310756 307640 310762 307652
rect 311434 307640 311440 307652
rect 311492 307640 311498 307692
rect 323762 307640 323768 307692
rect 323820 307680 323826 307692
rect 334066 307680 334072 307692
rect 323820 307652 334072 307680
rect 323820 307640 323826 307652
rect 334066 307640 334072 307652
rect 334124 307680 334130 307692
rect 335262 307680 335268 307692
rect 334124 307652 335268 307680
rect 334124 307640 334130 307652
rect 335262 307640 335268 307652
rect 335320 307640 335326 307692
rect 292942 307572 292948 307624
rect 293000 307612 293006 307624
rect 293310 307612 293316 307624
rect 293000 307584 293316 307612
rect 293000 307572 293006 307584
rect 293310 307572 293316 307584
rect 293368 307612 293374 307624
rect 351362 307612 351368 307624
rect 293368 307584 351368 307612
rect 293368 307572 293374 307584
rect 351362 307572 351368 307584
rect 351420 307572 351426 307624
rect 291102 307504 291108 307556
rect 291160 307544 291166 307556
rect 348418 307544 348424 307556
rect 291160 307516 348424 307544
rect 291160 307504 291166 307516
rect 348418 307504 348424 307516
rect 348476 307504 348482 307556
rect 281902 307436 281908 307488
rect 281960 307476 281966 307488
rect 299474 307476 299480 307488
rect 281960 307448 299480 307476
rect 281960 307436 281966 307448
rect 299474 307436 299480 307448
rect 299532 307476 299538 307488
rect 356698 307476 356704 307488
rect 299532 307448 356704 307476
rect 299532 307436 299538 307448
rect 356698 307436 356704 307448
rect 356756 307436 356762 307488
rect 280706 307368 280712 307420
rect 280764 307408 280770 307420
rect 290826 307408 290832 307420
rect 280764 307380 290832 307408
rect 280764 307368 280770 307380
rect 290826 307368 290832 307380
rect 290884 307408 290890 307420
rect 291102 307408 291108 307420
rect 290884 307380 291108 307408
rect 290884 307368 290890 307380
rect 291102 307368 291108 307380
rect 291160 307368 291166 307420
rect 294230 307368 294236 307420
rect 294288 307408 294294 307420
rect 347130 307408 347136 307420
rect 294288 307380 347136 307408
rect 294288 307368 294294 307380
rect 347130 307368 347136 307380
rect 347188 307368 347194 307420
rect 285214 307300 285220 307352
rect 285272 307340 285278 307352
rect 298094 307340 298100 307352
rect 285272 307312 298100 307340
rect 285272 307300 285278 307312
rect 298094 307300 298100 307312
rect 298152 307340 298158 307352
rect 344554 307340 344560 307352
rect 298152 307312 344560 307340
rect 298152 307300 298158 307312
rect 344554 307300 344560 307312
rect 344612 307300 344618 307352
rect 285490 307232 285496 307284
rect 285548 307272 285554 307284
rect 331858 307272 331864 307284
rect 285548 307244 331864 307272
rect 285548 307232 285554 307244
rect 331858 307232 331864 307244
rect 331916 307232 331922 307284
rect 213362 307164 213368 307216
rect 213420 307204 213426 307216
rect 263134 307204 263140 307216
rect 213420 307176 263140 307204
rect 213420 307164 213426 307176
rect 263134 307164 263140 307176
rect 263192 307164 263198 307216
rect 283834 307164 283840 307216
rect 283892 307204 283898 307216
rect 283892 307176 293908 307204
rect 283892 307164 283898 307176
rect 217502 307096 217508 307148
rect 217560 307136 217566 307148
rect 293218 307136 293224 307148
rect 217560 307108 293224 307136
rect 217560 307096 217566 307108
rect 293218 307096 293224 307108
rect 293276 307096 293282 307148
rect 293880 307136 293908 307176
rect 293954 307164 293960 307216
rect 294012 307204 294018 307216
rect 294966 307204 294972 307216
rect 294012 307176 294972 307204
rect 294012 307164 294018 307176
rect 294966 307164 294972 307176
rect 295024 307204 295030 307216
rect 337654 307204 337660 307216
rect 295024 307176 337660 307204
rect 295024 307164 295030 307176
rect 337654 307164 337660 307176
rect 337712 307164 337718 307216
rect 294046 307136 294052 307148
rect 293880 307108 294052 307136
rect 294046 307096 294052 307108
rect 294104 307096 294110 307148
rect 314470 307096 314476 307148
rect 314528 307136 314534 307148
rect 355410 307136 355416 307148
rect 314528 307108 355416 307136
rect 314528 307096 314534 307108
rect 355410 307096 355416 307108
rect 355468 307096 355474 307148
rect 217594 307028 217600 307080
rect 217652 307068 217658 307080
rect 299934 307068 299940 307080
rect 217652 307040 299940 307068
rect 217652 307028 217658 307040
rect 299934 307028 299940 307040
rect 299992 307028 299998 307080
rect 314930 307028 314936 307080
rect 314988 307068 314994 307080
rect 315574 307068 315580 307080
rect 314988 307040 315580 307068
rect 314988 307028 314994 307040
rect 315574 307028 315580 307040
rect 315632 307068 315638 307080
rect 376294 307068 376300 307080
rect 315632 307040 376300 307068
rect 315632 307028 315638 307040
rect 376294 307028 376300 307040
rect 376352 307068 376358 307080
rect 431954 307068 431960 307080
rect 376352 307040 431960 307068
rect 376352 307028 376358 307040
rect 431954 307028 431960 307040
rect 432012 307028 432018 307080
rect 311434 306960 311440 307012
rect 311492 307000 311498 307012
rect 370498 307000 370504 307012
rect 311492 306972 370504 307000
rect 311492 306960 311498 306972
rect 370498 306960 370504 306972
rect 370556 306960 370562 307012
rect 313550 306892 313556 306944
rect 313608 306932 313614 306944
rect 314470 306932 314476 306944
rect 313608 306904 314476 306932
rect 313608 306892 313614 306904
rect 314470 306892 314476 306904
rect 314528 306892 314534 306944
rect 209222 306348 209228 306400
rect 209280 306388 209286 306400
rect 266998 306388 267004 306400
rect 209280 306360 267004 306388
rect 209280 306348 209286 306360
rect 266998 306348 267004 306360
rect 267056 306348 267062 306400
rect 266354 306280 266360 306332
rect 266412 306320 266418 306332
rect 267642 306320 267648 306332
rect 266412 306292 267648 306320
rect 266412 306280 266418 306292
rect 267642 306280 267648 306292
rect 267700 306320 267706 306332
rect 286410 306320 286416 306332
rect 267700 306292 286416 306320
rect 267700 306280 267706 306292
rect 286410 306280 286416 306292
rect 286468 306280 286474 306332
rect 305178 306280 305184 306332
rect 305236 306320 305242 306332
rect 365806 306320 365812 306332
rect 305236 306292 365812 306320
rect 305236 306280 305242 306292
rect 365806 306280 365812 306292
rect 365864 306280 365870 306332
rect 308214 306212 308220 306264
rect 308272 306252 308278 306264
rect 367922 306252 367928 306264
rect 308272 306224 367928 306252
rect 308272 306212 308278 306224
rect 367922 306212 367928 306224
rect 367980 306212 367986 306264
rect 308122 306144 308128 306196
rect 308180 306184 308186 306196
rect 367830 306184 367836 306196
rect 308180 306156 367836 306184
rect 308180 306144 308186 306156
rect 367830 306144 367836 306156
rect 367888 306144 367894 306196
rect 293218 306076 293224 306128
rect 293276 306116 293282 306128
rect 309778 306116 309784 306128
rect 293276 306088 309784 306116
rect 293276 306076 293282 306088
rect 309778 306076 309784 306088
rect 309836 306116 309842 306128
rect 365070 306116 365076 306128
rect 309836 306088 365076 306116
rect 309836 306076 309842 306088
rect 365070 306076 365076 306088
rect 365128 306076 365134 306128
rect 285858 306008 285864 306060
rect 285916 306048 285922 306060
rect 339034 306048 339040 306060
rect 285916 306020 339040 306048
rect 285916 306008 285922 306020
rect 339034 306008 339040 306020
rect 339092 306008 339098 306060
rect 296070 305940 296076 305992
rect 296128 305980 296134 305992
rect 308122 305980 308128 305992
rect 296128 305952 308128 305980
rect 296128 305940 296134 305952
rect 308122 305940 308128 305952
rect 308180 305940 308186 305992
rect 309594 305940 309600 305992
rect 309652 305980 309658 305992
rect 362218 305980 362224 305992
rect 309652 305952 362224 305980
rect 309652 305940 309658 305952
rect 362218 305940 362224 305952
rect 362276 305940 362282 305992
rect 292850 305872 292856 305924
rect 292908 305912 292914 305924
rect 344278 305912 344284 305924
rect 292908 305884 344284 305912
rect 292908 305872 292914 305884
rect 344278 305872 344284 305884
rect 344336 305872 344342 305924
rect 286318 305804 286324 305856
rect 286376 305844 286382 305856
rect 302510 305844 302516 305856
rect 286376 305816 302516 305844
rect 286376 305804 286382 305816
rect 302510 305804 302516 305816
rect 302568 305844 302574 305856
rect 348694 305844 348700 305856
rect 302568 305816 348700 305844
rect 302568 305804 302574 305816
rect 348694 305804 348700 305816
rect 348752 305804 348758 305856
rect 291470 305736 291476 305788
rect 291528 305776 291534 305788
rect 335998 305776 336004 305788
rect 291528 305748 336004 305776
rect 291528 305736 291534 305748
rect 335998 305736 336004 305748
rect 336056 305736 336062 305788
rect 210694 305668 210700 305720
rect 210752 305708 210758 305720
rect 266354 305708 266360 305720
rect 210752 305680 266360 305708
rect 210752 305668 210758 305680
rect 266354 305668 266360 305680
rect 266412 305668 266418 305720
rect 330478 305708 330484 305720
rect 296686 305680 330484 305708
rect 214834 305600 214840 305652
rect 214892 305640 214898 305652
rect 292850 305640 292856 305652
rect 214892 305612 292856 305640
rect 214892 305600 214898 305612
rect 292850 305600 292856 305612
rect 292908 305600 292914 305652
rect 290090 305532 290096 305584
rect 290148 305572 290154 305584
rect 291010 305572 291016 305584
rect 290148 305544 291016 305572
rect 290148 305532 290154 305544
rect 291010 305532 291016 305544
rect 291068 305572 291074 305584
rect 296686 305572 296714 305680
rect 330478 305668 330484 305680
rect 330536 305668 330542 305720
rect 307386 305600 307392 305652
rect 307444 305640 307450 305652
rect 343082 305640 343088 305652
rect 307444 305612 343088 305640
rect 307444 305600 307450 305612
rect 343082 305600 343088 305612
rect 343140 305600 343146 305652
rect 334894 305572 334900 305584
rect 291068 305544 296714 305572
rect 306346 305544 334900 305572
rect 291068 305532 291074 305544
rect 299750 305396 299756 305448
rect 299808 305436 299814 305448
rect 300578 305436 300584 305448
rect 299808 305408 300584 305436
rect 299808 305396 299814 305408
rect 300578 305396 300584 305408
rect 300636 305436 300642 305448
rect 306346 305436 306374 305544
rect 334894 305532 334900 305544
rect 334952 305532 334958 305584
rect 322750 305464 322756 305516
rect 322808 305504 322814 305516
rect 349890 305504 349896 305516
rect 322808 305476 349896 305504
rect 322808 305464 322814 305476
rect 349890 305464 349896 305476
rect 349948 305464 349954 305516
rect 300636 305408 306374 305436
rect 300636 305396 300642 305408
rect 306742 305396 306748 305448
rect 306800 305436 306806 305448
rect 307386 305436 307392 305448
rect 306800 305408 307392 305436
rect 306800 305396 306806 305408
rect 307386 305396 307392 305408
rect 307444 305396 307450 305448
rect 314102 305396 314108 305448
rect 314160 305436 314166 305448
rect 339586 305436 339592 305448
rect 314160 305408 339592 305436
rect 314160 305396 314166 305408
rect 339586 305396 339592 305408
rect 339644 305396 339650 305448
rect 321646 305124 321652 305176
rect 321704 305164 321710 305176
rect 322750 305164 322756 305176
rect 321704 305136 322756 305164
rect 321704 305124 321710 305136
rect 322750 305124 322756 305136
rect 322808 305124 322814 305176
rect 216030 305056 216036 305108
rect 216088 305096 216094 305108
rect 259638 305096 259644 305108
rect 216088 305068 259644 305096
rect 216088 305056 216094 305068
rect 259638 305056 259644 305068
rect 259696 305056 259702 305108
rect 206278 304988 206284 305040
rect 206336 305028 206342 305040
rect 265894 305028 265900 305040
rect 206336 305000 265900 305028
rect 206336 304988 206342 305000
rect 265894 304988 265900 305000
rect 265952 304988 265958 305040
rect 288158 304988 288164 305040
rect 288216 305028 288222 305040
rect 291470 305028 291476 305040
rect 288216 305000 291476 305028
rect 288216 304988 288222 305000
rect 291470 304988 291476 305000
rect 291528 304988 291534 305040
rect 305178 304988 305184 305040
rect 305236 305028 305242 305040
rect 305638 305028 305644 305040
rect 305236 305000 305644 305028
rect 305236 304988 305242 305000
rect 305638 304988 305644 305000
rect 305696 304988 305702 305040
rect 308214 304988 308220 305040
rect 308272 305028 308278 305040
rect 308582 305028 308588 305040
rect 308272 305000 308588 305028
rect 308272 304988 308278 305000
rect 308582 304988 308588 305000
rect 308640 304988 308646 305040
rect 339586 304988 339592 305040
rect 339644 305028 339650 305040
rect 340782 305028 340788 305040
rect 339644 305000 340788 305028
rect 339644 304988 339650 305000
rect 340782 304988 340788 305000
rect 340840 304988 340846 305040
rect 282638 304920 282644 304972
rect 282696 304960 282702 304972
rect 359550 304960 359556 304972
rect 282696 304932 359556 304960
rect 282696 304920 282702 304932
rect 359550 304920 359556 304932
rect 359608 304920 359614 304972
rect 264974 304852 264980 304904
rect 265032 304892 265038 304904
rect 266170 304892 266176 304904
rect 265032 304864 266176 304892
rect 265032 304852 265038 304864
rect 266170 304852 266176 304864
rect 266228 304892 266234 304904
rect 288986 304892 288992 304904
rect 266228 304864 288992 304892
rect 266228 304852 266234 304864
rect 288986 304852 288992 304864
rect 289044 304852 289050 304904
rect 295334 304852 295340 304904
rect 295392 304892 295398 304904
rect 295610 304892 295616 304904
rect 295392 304864 295616 304892
rect 295392 304852 295398 304864
rect 295610 304852 295616 304864
rect 295668 304892 295674 304904
rect 357066 304892 357072 304904
rect 295668 304864 357072 304892
rect 295668 304852 295674 304864
rect 357066 304852 357072 304864
rect 357124 304852 357130 304904
rect 271782 304784 271788 304836
rect 271840 304824 271846 304836
rect 291378 304824 291384 304836
rect 271840 304796 291384 304824
rect 271840 304784 271846 304796
rect 291378 304784 291384 304796
rect 291436 304784 291442 304836
rect 302418 304784 302424 304836
rect 302476 304824 302482 304836
rect 360838 304824 360844 304836
rect 302476 304796 360844 304824
rect 302476 304784 302482 304796
rect 360838 304784 360844 304796
rect 360896 304784 360902 304836
rect 266998 304716 267004 304768
rect 267056 304756 267062 304768
rect 283098 304756 283104 304768
rect 267056 304728 283104 304756
rect 267056 304716 267062 304728
rect 283098 304716 283104 304728
rect 283156 304716 283162 304768
rect 300946 304716 300952 304768
rect 301004 304756 301010 304768
rect 351270 304756 351276 304768
rect 301004 304728 351276 304756
rect 301004 304716 301010 304728
rect 351270 304716 351276 304728
rect 351328 304716 351334 304768
rect 299658 304648 299664 304700
rect 299716 304688 299722 304700
rect 349798 304688 349804 304700
rect 299716 304660 349804 304688
rect 299716 304648 299722 304660
rect 349798 304648 349804 304660
rect 349856 304648 349862 304700
rect 261294 304580 261300 304632
rect 261352 304620 261358 304632
rect 261754 304620 261760 304632
rect 261352 304592 261760 304620
rect 261352 304580 261358 304592
rect 261754 304580 261760 304592
rect 261812 304580 261818 304632
rect 298646 304580 298652 304632
rect 298704 304620 298710 304632
rect 347314 304620 347320 304632
rect 298704 304592 347320 304620
rect 298704 304580 298710 304592
rect 347314 304580 347320 304592
rect 347372 304580 347378 304632
rect 220630 304512 220636 304564
rect 220688 304552 220694 304564
rect 271782 304552 271788 304564
rect 220688 304524 271788 304552
rect 220688 304512 220694 304524
rect 271782 304512 271788 304524
rect 271840 304512 271846 304564
rect 286686 304512 286692 304564
rect 286744 304552 286750 304564
rect 301222 304552 301228 304564
rect 286744 304524 301228 304552
rect 286744 304512 286750 304524
rect 301222 304512 301228 304524
rect 301280 304552 301286 304564
rect 348510 304552 348516 304564
rect 301280 304524 348516 304552
rect 301280 304512 301286 304524
rect 348510 304512 348516 304524
rect 348568 304512 348574 304564
rect 208118 304444 208124 304496
rect 208176 304484 208182 304496
rect 264974 304484 264980 304496
rect 208176 304456 264980 304484
rect 208176 304444 208182 304456
rect 264974 304444 264980 304456
rect 265032 304444 265038 304496
rect 293310 304444 293316 304496
rect 293368 304484 293374 304496
rect 300946 304484 300952 304496
rect 293368 304456 300952 304484
rect 293368 304444 293374 304456
rect 300946 304444 300952 304456
rect 301004 304444 301010 304496
rect 301130 304444 301136 304496
rect 301188 304484 301194 304496
rect 345934 304484 345940 304496
rect 301188 304456 345940 304484
rect 301188 304444 301194 304456
rect 345934 304444 345940 304456
rect 345992 304444 345998 304496
rect 218882 304376 218888 304428
rect 218940 304416 218946 304428
rect 218940 304388 296714 304416
rect 218940 304376 218946 304388
rect 208026 304308 208032 304360
rect 208084 304348 208090 304360
rect 285858 304348 285864 304360
rect 208084 304320 285864 304348
rect 208084 304308 208090 304320
rect 285858 304308 285864 304320
rect 285916 304308 285922 304360
rect 296686 304348 296714 304388
rect 301038 304376 301044 304428
rect 301096 304416 301102 304428
rect 344462 304416 344468 304428
rect 301096 304388 344468 304416
rect 301096 304376 301102 304388
rect 344462 304376 344468 304388
rect 344520 304376 344526 304428
rect 296898 304348 296904 304360
rect 296686 304320 296904 304348
rect 296898 304308 296904 304320
rect 296956 304348 296962 304360
rect 340322 304348 340328 304360
rect 296956 304320 340328 304348
rect 296956 304308 296962 304320
rect 340322 304308 340328 304320
rect 340380 304308 340386 304360
rect 213270 304240 213276 304292
rect 213328 304280 213334 304292
rect 295334 304280 295340 304292
rect 213328 304252 295340 304280
rect 213328 304240 213334 304252
rect 295334 304240 295340 304252
rect 295392 304240 295398 304292
rect 299566 304240 299572 304292
rect 299624 304280 299630 304292
rect 348602 304280 348608 304292
rect 299624 304252 348608 304280
rect 299624 304240 299630 304252
rect 348602 304240 348608 304252
rect 348660 304240 348666 304292
rect 300486 304172 300492 304224
rect 300544 304212 300550 304224
rect 341610 304212 341616 304224
rect 300544 304184 341616 304212
rect 300544 304172 300550 304184
rect 341610 304172 341616 304184
rect 341668 304172 341674 304224
rect 299106 304104 299112 304156
rect 299164 304144 299170 304156
rect 334710 304144 334716 304156
rect 299164 304116 334716 304144
rect 299164 304104 299170 304116
rect 334710 304104 334716 304116
rect 334768 304104 334774 304156
rect 284110 304036 284116 304088
rect 284168 304076 284174 304088
rect 302418 304076 302424 304088
rect 284168 304048 302424 304076
rect 284168 304036 284174 304048
rect 302418 304036 302424 304048
rect 302476 304036 302482 304088
rect 307018 304036 307024 304088
rect 307076 304076 307082 304088
rect 313182 304076 313188 304088
rect 307076 304048 313188 304076
rect 307076 304036 307082 304048
rect 313182 304036 313188 304048
rect 313240 304076 313246 304088
rect 334802 304076 334808 304088
rect 313240 304048 334808 304076
rect 313240 304036 313246 304048
rect 334802 304036 334808 304048
rect 334860 304036 334866 304088
rect 298554 303968 298560 304020
rect 298612 304008 298618 304020
rect 299566 304008 299572 304020
rect 298612 303980 299572 304008
rect 298612 303968 298618 303980
rect 299566 303968 299572 303980
rect 299624 303968 299630 304020
rect 264054 303804 264060 303816
rect 258046 303776 264060 303804
rect 204530 303696 204536 303748
rect 204588 303736 204594 303748
rect 258046 303736 258074 303776
rect 264054 303764 264060 303776
rect 264112 303804 264118 303816
rect 264514 303804 264520 303816
rect 264112 303776 264520 303804
rect 264112 303764 264118 303776
rect 264514 303764 264520 303776
rect 264572 303764 264578 303816
rect 204588 303708 258074 303736
rect 204588 303696 204594 303708
rect 297450 303696 297456 303748
rect 297508 303736 297514 303748
rect 301130 303736 301136 303748
rect 297508 303708 301136 303736
rect 297508 303696 297514 303708
rect 301130 303696 301136 303708
rect 301188 303696 301194 303748
rect 201402 303628 201408 303680
rect 201460 303668 201466 303680
rect 261294 303668 261300 303680
rect 201460 303640 261300 303668
rect 201460 303628 201466 303640
rect 261294 303628 261300 303640
rect 261352 303628 261358 303680
rect 298646 303628 298652 303680
rect 298704 303668 298710 303680
rect 299014 303668 299020 303680
rect 298704 303640 299020 303668
rect 298704 303628 298710 303640
rect 299014 303628 299020 303640
rect 299072 303628 299078 303680
rect 299658 303628 299664 303680
rect 299716 303668 299722 303680
rect 300118 303668 300124 303680
rect 299716 303640 300124 303668
rect 299716 303628 299722 303640
rect 300118 303628 300124 303640
rect 300176 303628 300182 303680
rect 301038 303628 301044 303680
rect 301096 303668 301102 303680
rect 301590 303668 301596 303680
rect 301096 303640 301596 303668
rect 301096 303628 301102 303640
rect 301590 303628 301596 303640
rect 301648 303628 301654 303680
rect 317506 303560 317512 303612
rect 317564 303600 317570 303612
rect 390554 303600 390560 303612
rect 317564 303572 390560 303600
rect 317564 303560 317570 303572
rect 390554 303560 390560 303572
rect 390612 303560 390618 303612
rect 320726 303492 320732 303544
rect 320784 303532 320790 303544
rect 320910 303532 320916 303544
rect 320784 303504 320916 303532
rect 320784 303492 320790 303504
rect 320910 303492 320916 303504
rect 320968 303532 320974 303544
rect 390646 303532 390652 303544
rect 320968 303504 390652 303532
rect 320968 303492 320974 303504
rect 390646 303492 390652 303504
rect 390704 303492 390710 303544
rect 301774 303424 301780 303476
rect 301832 303464 301838 303476
rect 362126 303464 362132 303476
rect 301832 303436 362132 303464
rect 301832 303424 301838 303436
rect 362126 303424 362132 303436
rect 362184 303424 362190 303476
rect 320910 303356 320916 303408
rect 320968 303396 320974 303408
rect 321094 303396 321100 303408
rect 320968 303368 321100 303396
rect 320968 303356 320974 303368
rect 321094 303356 321100 303368
rect 321152 303356 321158 303408
rect 321186 303356 321192 303408
rect 321244 303396 321250 303408
rect 380158 303396 380164 303408
rect 321244 303368 380164 303396
rect 321244 303356 321250 303368
rect 380158 303356 380164 303368
rect 380216 303356 380222 303408
rect 320174 303288 320180 303340
rect 320232 303328 320238 303340
rect 320232 303300 321416 303328
rect 320232 303288 320238 303300
rect 321388 303272 321416 303300
rect 321462 303288 321468 303340
rect 321520 303328 321526 303340
rect 380066 303328 380072 303340
rect 321520 303300 380072 303328
rect 321520 303288 321526 303300
rect 380066 303288 380072 303300
rect 380124 303288 380130 303340
rect 321094 303220 321100 303272
rect 321152 303260 321158 303272
rect 321278 303260 321284 303272
rect 321152 303232 321284 303260
rect 321152 303220 321158 303232
rect 321278 303220 321284 303232
rect 321336 303220 321342 303272
rect 321370 303220 321376 303272
rect 321428 303260 321434 303272
rect 380342 303260 380348 303272
rect 321428 303232 380348 303260
rect 321428 303220 321434 303232
rect 380342 303220 380348 303232
rect 380400 303220 380406 303272
rect 295334 303152 295340 303204
rect 295392 303192 295398 303204
rect 296438 303192 296444 303204
rect 295392 303164 296444 303192
rect 295392 303152 295398 303164
rect 296438 303152 296444 303164
rect 296496 303192 296502 303204
rect 354030 303192 354036 303204
rect 296496 303164 354036 303192
rect 296496 303152 296502 303164
rect 354030 303152 354036 303164
rect 354088 303152 354094 303204
rect 292022 303084 292028 303136
rect 292080 303124 292086 303136
rect 294138 303124 294144 303136
rect 292080 303096 294144 303124
rect 292080 303084 292086 303096
rect 294138 303084 294144 303096
rect 294196 303124 294202 303136
rect 351178 303124 351184 303136
rect 294196 303096 351184 303124
rect 294196 303084 294202 303096
rect 351178 303084 351184 303096
rect 351236 303084 351242 303136
rect 288250 303016 288256 303068
rect 288308 303056 288314 303068
rect 295518 303056 295524 303068
rect 288308 303028 295524 303056
rect 288308 303016 288314 303028
rect 295518 303016 295524 303028
rect 295576 303056 295582 303068
rect 352558 303056 352564 303068
rect 295576 303028 352564 303056
rect 295576 303016 295582 303028
rect 352558 303016 352564 303028
rect 352616 303016 352622 303068
rect 213822 302948 213828 303000
rect 213880 302988 213886 303000
rect 291746 302988 291752 303000
rect 213880 302960 291752 302988
rect 213880 302948 213886 302960
rect 291746 302948 291752 302960
rect 291804 302988 291810 303000
rect 340230 302988 340236 303000
rect 291804 302960 340236 302988
rect 291804 302948 291810 302960
rect 340230 302948 340236 302960
rect 340288 302948 340294 303000
rect 215938 302880 215944 302932
rect 215996 302920 216002 302932
rect 295334 302920 295340 302932
rect 215996 302892 295340 302920
rect 215996 302880 216002 302892
rect 295334 302880 295340 302892
rect 295392 302880 295398 302932
rect 298002 302880 298008 302932
rect 298060 302920 298066 302932
rect 337470 302920 337476 302932
rect 298060 302892 337476 302920
rect 298060 302880 298066 302892
rect 337470 302880 337476 302892
rect 337528 302880 337534 302932
rect 305362 302812 305368 302864
rect 305420 302852 305426 302864
rect 329190 302852 329196 302864
rect 305420 302824 329196 302852
rect 305420 302812 305426 302824
rect 329190 302812 329196 302824
rect 329248 302812 329254 302864
rect 301958 302744 301964 302796
rect 302016 302784 302022 302796
rect 303890 302784 303896 302796
rect 302016 302756 303896 302784
rect 302016 302744 302022 302756
rect 303890 302744 303896 302756
rect 303948 302784 303954 302796
rect 343174 302784 343180 302796
rect 303948 302756 343180 302784
rect 303948 302744 303954 302756
rect 343174 302744 343180 302756
rect 343232 302744 343238 302796
rect 300026 302676 300032 302728
rect 300084 302716 300090 302728
rect 343266 302716 343272 302728
rect 300084 302688 343272 302716
rect 300084 302676 300090 302688
rect 343266 302676 343272 302688
rect 343324 302676 343330 302728
rect 204346 302268 204352 302320
rect 204404 302308 204410 302320
rect 204404 302280 264560 302308
rect 204404 302268 204410 302280
rect 264532 302252 264560 302280
rect 200114 302200 200120 302252
rect 200172 302240 200178 302252
rect 260926 302240 260932 302252
rect 200172 302212 260932 302240
rect 200172 302200 200178 302212
rect 260926 302200 260932 302212
rect 260984 302240 260990 302252
rect 260984 302212 262168 302240
rect 260984 302200 260990 302212
rect 262140 302172 262168 302212
rect 264514 302200 264520 302252
rect 264572 302240 264578 302252
rect 264882 302240 264888 302252
rect 264572 302212 264888 302240
rect 264572 302200 264578 302212
rect 264882 302200 264888 302212
rect 264940 302200 264946 302252
rect 296806 302200 296812 302252
rect 296864 302240 296870 302252
rect 298002 302240 298008 302252
rect 296864 302212 298008 302240
rect 296864 302200 296870 302212
rect 298002 302200 298008 302212
rect 298060 302200 298066 302252
rect 269942 302172 269948 302184
rect 262140 302144 269948 302172
rect 269942 302132 269948 302144
rect 270000 302132 270006 302184
rect 297542 302132 297548 302184
rect 297600 302172 297606 302184
rect 360562 302172 360568 302184
rect 297600 302144 360568 302172
rect 297600 302132 297606 302144
rect 360562 302132 360568 302144
rect 360620 302132 360626 302184
rect 289354 302064 289360 302116
rect 289412 302104 289418 302116
rect 296346 302104 296352 302116
rect 289412 302076 296352 302104
rect 289412 302064 289418 302076
rect 296346 302064 296352 302076
rect 296404 302104 296410 302116
rect 357802 302104 357808 302116
rect 296404 302076 357808 302104
rect 296404 302064 296410 302076
rect 357802 302064 357808 302076
rect 357860 302064 357866 302116
rect 312906 301996 312912 302048
rect 312964 302036 312970 302048
rect 374454 302036 374460 302048
rect 312964 302008 374460 302036
rect 312964 301996 312970 302008
rect 374454 301996 374460 302008
rect 374512 301996 374518 302048
rect 309778 301928 309784 301980
rect 309836 301968 309842 301980
rect 371694 301968 371700 301980
rect 309836 301940 371700 301968
rect 309836 301928 309842 301940
rect 371694 301928 371700 301940
rect 371752 301928 371758 301980
rect 307202 301860 307208 301912
rect 307260 301900 307266 301912
rect 307662 301900 307668 301912
rect 307260 301872 307668 301900
rect 307260 301860 307266 301872
rect 307662 301860 307668 301872
rect 307720 301900 307726 301912
rect 368842 301900 368848 301912
rect 307720 301872 368848 301900
rect 307720 301860 307726 301872
rect 368842 301860 368848 301872
rect 368900 301860 368906 301912
rect 300762 301792 300768 301844
rect 300820 301832 300826 301844
rect 361942 301832 361948 301844
rect 300820 301804 361948 301832
rect 300820 301792 300826 301804
rect 361942 301792 361948 301804
rect 362000 301792 362006 301844
rect 297542 301724 297548 301776
rect 297600 301764 297606 301776
rect 297910 301764 297916 301776
rect 297600 301736 297916 301764
rect 297600 301724 297606 301736
rect 297910 301724 297916 301736
rect 297968 301724 297974 301776
rect 309226 301724 309232 301776
rect 309284 301764 309290 301776
rect 310146 301764 310152 301776
rect 309284 301736 310152 301764
rect 309284 301724 309290 301736
rect 310146 301724 310152 301736
rect 310204 301724 310210 301776
rect 370314 301764 370320 301776
rect 310256 301736 370320 301764
rect 309318 301656 309324 301708
rect 309376 301696 309382 301708
rect 309778 301696 309784 301708
rect 309376 301668 309784 301696
rect 309376 301656 309382 301668
rect 309778 301656 309784 301668
rect 309836 301656 309842 301708
rect 310256 301640 310284 301736
rect 370314 301724 370320 301736
rect 370372 301724 370378 301776
rect 312078 301656 312084 301708
rect 312136 301696 312142 301708
rect 312354 301696 312360 301708
rect 312136 301668 312360 301696
rect 312136 301656 312142 301668
rect 312354 301656 312360 301668
rect 312412 301696 312418 301708
rect 372246 301696 372252 301708
rect 312412 301668 372252 301696
rect 312412 301656 312418 301668
rect 372246 301656 372252 301668
rect 372304 301656 372310 301708
rect 309410 301588 309416 301640
rect 309468 301628 309474 301640
rect 310238 301628 310244 301640
rect 309468 301600 310244 301628
rect 309468 301588 309474 301600
rect 310238 301588 310244 301600
rect 310296 301588 310302 301640
rect 310330 301588 310336 301640
rect 310388 301628 310394 301640
rect 369026 301628 369032 301640
rect 310388 301600 369032 301628
rect 310388 301588 310394 301600
rect 369026 301588 369032 301600
rect 369084 301588 369090 301640
rect 287514 301520 287520 301572
rect 287572 301560 287578 301572
rect 287882 301560 287888 301572
rect 287572 301532 287888 301560
rect 287572 301520 287578 301532
rect 287882 301520 287888 301532
rect 287940 301560 287946 301572
rect 345658 301560 345664 301572
rect 287940 301532 345664 301560
rect 287940 301520 287946 301532
rect 345658 301520 345664 301532
rect 345716 301520 345722 301572
rect 224310 301452 224316 301504
rect 224368 301492 224374 301504
rect 293402 301492 293408 301504
rect 224368 301464 293408 301492
rect 224368 301452 224374 301464
rect 293402 301452 293408 301464
rect 293460 301452 293466 301504
rect 298370 301452 298376 301504
rect 298428 301492 298434 301504
rect 351454 301492 351460 301504
rect 298428 301464 351460 301492
rect 298428 301452 298434 301464
rect 351454 301452 351460 301464
rect 351512 301452 351518 301504
rect 305914 301384 305920 301436
rect 305972 301424 305978 301436
rect 344370 301424 344376 301436
rect 305972 301396 344376 301424
rect 305972 301384 305978 301396
rect 344370 301384 344376 301396
rect 344428 301384 344434 301436
rect 256694 301316 256700 301368
rect 256752 301356 256758 301368
rect 257246 301356 257252 301368
rect 256752 301328 257252 301356
rect 256752 301316 256758 301328
rect 257246 301316 257252 301328
rect 257304 301316 257310 301368
rect 262306 301316 262312 301368
rect 262364 301356 262370 301368
rect 262950 301356 262956 301368
rect 262364 301328 262956 301356
rect 262364 301316 262370 301328
rect 262950 301316 262956 301328
rect 263008 301316 263014 301368
rect 320726 301316 320732 301368
rect 320784 301356 320790 301368
rect 321278 301356 321284 301368
rect 320784 301328 321284 301356
rect 320784 301316 320790 301328
rect 321278 301316 321284 301328
rect 321336 301316 321342 301368
rect 197354 300908 197360 300960
rect 197412 300948 197418 300960
rect 256694 300948 256700 300960
rect 197412 300920 256700 300948
rect 197412 300908 197418 300920
rect 256694 300908 256700 300920
rect 256752 300908 256758 300960
rect 202782 300840 202788 300892
rect 202840 300880 202846 300892
rect 262306 300880 262312 300892
rect 202840 300852 262312 300880
rect 202840 300840 202846 300852
rect 262306 300840 262312 300852
rect 262364 300840 262370 300892
rect 255314 300772 255320 300824
rect 255372 300812 255378 300824
rect 256142 300812 256148 300824
rect 255372 300784 256148 300812
rect 255372 300772 255378 300784
rect 256142 300772 256148 300784
rect 256200 300772 256206 300824
rect 262398 300772 262404 300824
rect 262456 300812 262462 300824
rect 262858 300812 262864 300824
rect 262456 300784 262864 300812
rect 262456 300772 262462 300784
rect 262858 300772 262864 300784
rect 262916 300772 262922 300824
rect 308030 300772 308036 300824
rect 308088 300812 308094 300824
rect 308674 300812 308680 300824
rect 308088 300784 308680 300812
rect 308088 300772 308094 300784
rect 308674 300772 308680 300784
rect 308732 300772 308738 300824
rect 369854 300812 369860 300824
rect 310716 300784 369860 300812
rect 307478 300704 307484 300756
rect 307536 300744 307542 300756
rect 310716 300744 310744 300784
rect 369854 300772 369860 300784
rect 369912 300772 369918 300824
rect 307536 300716 310744 300744
rect 307536 300704 307542 300716
rect 312630 300704 312636 300756
rect 312688 300744 312694 300756
rect 312998 300744 313004 300756
rect 312688 300716 313004 300744
rect 312688 300704 312694 300716
rect 312998 300704 313004 300716
rect 313056 300744 313062 300756
rect 374362 300744 374368 300756
rect 313056 300716 374368 300744
rect 313056 300704 313062 300716
rect 374362 300704 374368 300716
rect 374420 300704 374426 300756
rect 300394 300636 300400 300688
rect 300452 300676 300458 300688
rect 306006 300676 306012 300688
rect 300452 300648 306012 300676
rect 300452 300636 300458 300648
rect 306006 300636 306012 300648
rect 306064 300676 306070 300688
rect 367646 300676 367652 300688
rect 306064 300648 367652 300676
rect 306064 300636 306070 300648
rect 367646 300636 367652 300648
rect 367704 300636 367710 300688
rect 304626 300568 304632 300620
rect 304684 300608 304690 300620
rect 364886 300608 364892 300620
rect 304684 300580 364892 300608
rect 304684 300568 304690 300580
rect 364886 300568 364892 300580
rect 364944 300568 364950 300620
rect 302326 300500 302332 300552
rect 302384 300540 302390 300552
rect 302970 300540 302976 300552
rect 302384 300512 302976 300540
rect 302384 300500 302390 300512
rect 302970 300500 302976 300512
rect 303028 300540 303034 300552
rect 363874 300540 363880 300552
rect 303028 300512 363880 300540
rect 303028 300500 303034 300512
rect 363874 300500 363880 300512
rect 363932 300500 363938 300552
rect 307662 300432 307668 300484
rect 307720 300472 307726 300484
rect 366542 300472 366548 300484
rect 307720 300444 366548 300472
rect 307720 300432 307726 300444
rect 366542 300432 366548 300444
rect 366600 300432 366606 300484
rect 318702 300364 318708 300416
rect 318760 300404 318766 300416
rect 377950 300404 377956 300416
rect 318760 300376 377956 300404
rect 318760 300364 318766 300376
rect 377950 300364 377956 300376
rect 378008 300364 378014 300416
rect 306926 300296 306932 300348
rect 306984 300336 306990 300348
rect 363598 300336 363604 300348
rect 306984 300308 363604 300336
rect 306984 300296 306990 300308
rect 363598 300296 363604 300308
rect 363656 300296 363662 300348
rect 303798 300268 303804 300280
rect 296686 300240 303804 300268
rect 289078 300092 289084 300144
rect 289136 300132 289142 300144
rect 296686 300132 296714 300240
rect 303798 300228 303804 300240
rect 303856 300268 303862 300280
rect 359458 300268 359464 300280
rect 303856 300240 359464 300268
rect 303856 300228 303862 300240
rect 359458 300228 359464 300240
rect 359516 300228 359522 300280
rect 305730 300160 305736 300212
rect 305788 300200 305794 300212
rect 306558 300200 306564 300212
rect 305788 300172 306564 300200
rect 305788 300160 305794 300172
rect 306558 300160 306564 300172
rect 306616 300200 306622 300212
rect 307662 300200 307668 300212
rect 306616 300172 307668 300200
rect 306616 300160 306622 300172
rect 307662 300160 307668 300172
rect 307720 300160 307726 300212
rect 307754 300160 307760 300212
rect 307812 300200 307818 300212
rect 349982 300200 349988 300212
rect 307812 300172 349988 300200
rect 307812 300160 307818 300172
rect 349982 300160 349988 300172
rect 350040 300160 350046 300212
rect 289136 300104 296714 300132
rect 289136 300092 289142 300104
rect 304350 300092 304356 300144
rect 304408 300132 304414 300144
rect 345842 300132 345848 300144
rect 304408 300104 345848 300132
rect 304408 300092 304414 300104
rect 345842 300092 345848 300104
rect 345900 300092 345906 300144
rect 230750 300024 230756 300076
rect 230808 300064 230814 300076
rect 231762 300064 231768 300076
rect 230808 300036 231768 300064
rect 230808 300024 230814 300036
rect 231762 300024 231768 300036
rect 231820 300024 231826 300076
rect 307202 300024 307208 300076
rect 307260 300064 307266 300076
rect 307662 300064 307668 300076
rect 307260 300036 307668 300064
rect 307260 300024 307266 300036
rect 307662 300024 307668 300036
rect 307720 300024 307726 300076
rect 308674 300024 308680 300076
rect 308732 300064 308738 300076
rect 340138 300064 340144 300076
rect 308732 300036 340144 300064
rect 308732 300024 308738 300036
rect 340138 300024 340144 300036
rect 340196 300024 340202 300076
rect 209038 299684 209044 299736
rect 209096 299724 209102 299736
rect 253198 299724 253204 299736
rect 209096 299696 253204 299724
rect 209096 299684 209102 299696
rect 253198 299684 253204 299696
rect 253256 299684 253262 299736
rect 195974 299616 195980 299668
rect 196032 299656 196038 299668
rect 256142 299656 256148 299668
rect 196032 299628 256148 299656
rect 196032 299616 196038 299628
rect 256142 299616 256148 299628
rect 256200 299616 256206 299668
rect 201678 299548 201684 299600
rect 201736 299588 201742 299600
rect 262398 299588 262404 299600
rect 201736 299560 262404 299588
rect 201736 299548 201742 299560
rect 262398 299548 262404 299560
rect 262456 299548 262462 299600
rect 231762 299480 231768 299532
rect 231820 299520 231826 299532
rect 577498 299520 577504 299532
rect 231820 299492 577504 299520
rect 231820 299480 231826 299492
rect 577498 299480 577504 299492
rect 577556 299480 577562 299532
rect 310330 299412 310336 299464
rect 310388 299452 310394 299464
rect 371602 299452 371608 299464
rect 310388 299424 371608 299452
rect 310388 299412 310394 299424
rect 371602 299412 371608 299424
rect 371660 299412 371666 299464
rect 316126 299344 316132 299396
rect 316184 299384 316190 299396
rect 316770 299384 316776 299396
rect 316184 299356 316776 299384
rect 316184 299344 316190 299356
rect 316770 299344 316776 299356
rect 316828 299344 316834 299396
rect 317414 299344 317420 299396
rect 317472 299384 317478 299396
rect 318058 299384 318064 299396
rect 317472 299356 318064 299384
rect 317472 299344 317478 299356
rect 318058 299344 318064 299356
rect 318116 299344 318122 299396
rect 318702 299344 318708 299396
rect 318760 299384 318766 299396
rect 378686 299384 378692 299396
rect 318760 299356 378692 299384
rect 318760 299344 318766 299356
rect 378686 299344 378692 299356
rect 378744 299344 378750 299396
rect 295058 299276 295064 299328
rect 295116 299316 295122 299328
rect 353938 299316 353944 299328
rect 295116 299288 353944 299316
rect 295116 299276 295122 299288
rect 353938 299276 353944 299288
rect 353996 299276 354002 299328
rect 310146 299208 310152 299260
rect 310204 299248 310210 299260
rect 310330 299248 310336 299260
rect 310204 299220 310336 299248
rect 310204 299208 310210 299220
rect 310330 299208 310336 299220
rect 310388 299208 310394 299260
rect 372706 299248 372712 299260
rect 316006 299220 372712 299248
rect 310054 299140 310060 299192
rect 310112 299180 310118 299192
rect 314286 299180 314292 299192
rect 310112 299152 314292 299180
rect 310112 299140 310118 299152
rect 314286 299140 314292 299152
rect 314344 299180 314350 299192
rect 316006 299180 316034 299220
rect 372706 299208 372712 299220
rect 372764 299208 372770 299260
rect 314344 299152 316034 299180
rect 314344 299140 314350 299152
rect 318058 299140 318064 299192
rect 318116 299180 318122 299192
rect 377674 299180 377680 299192
rect 318116 299152 377680 299180
rect 318116 299140 318122 299152
rect 377674 299140 377680 299152
rect 377732 299140 377738 299192
rect 316770 299072 316776 299124
rect 316828 299112 316834 299124
rect 376202 299112 376208 299124
rect 316828 299084 376208 299112
rect 316828 299072 316834 299084
rect 376202 299072 376208 299084
rect 376260 299072 376266 299124
rect 311710 299004 311716 299056
rect 311768 299044 311774 299056
rect 364978 299044 364984 299056
rect 311768 299016 364984 299044
rect 311768 299004 311774 299016
rect 364978 299004 364984 299016
rect 365036 299004 365042 299056
rect 285582 298936 285588 298988
rect 285640 298976 285646 298988
rect 337562 298976 337568 298988
rect 285640 298948 337568 298976
rect 285640 298936 285646 298948
rect 337562 298936 337568 298948
rect 337620 298936 337626 298988
rect 4154 298800 4160 298852
rect 4212 298840 4218 298852
rect 221918 298840 221924 298852
rect 4212 298812 221924 298840
rect 4212 298800 4218 298812
rect 221918 298800 221924 298812
rect 221976 298800 221982 298852
rect 233142 298732 233148 298784
rect 233200 298772 233206 298784
rect 580166 298772 580172 298784
rect 233200 298744 580172 298772
rect 233200 298732 233206 298744
rect 580166 298732 580172 298744
rect 580224 298732 580230 298784
rect 207842 298256 207848 298308
rect 207900 298296 207906 298308
rect 265618 298296 265624 298308
rect 207900 298268 265624 298296
rect 207900 298256 207906 298268
rect 265618 298256 265624 298268
rect 265676 298296 265682 298308
rect 265676 298268 265848 298296
rect 265676 298256 265682 298268
rect 202874 298188 202880 298240
rect 202932 298228 202938 298240
rect 263042 298228 263048 298240
rect 202932 298200 263048 298228
rect 202932 298188 202938 298200
rect 263042 298188 263048 298200
rect 263100 298188 263106 298240
rect 194594 298120 194600 298172
rect 194652 298160 194658 298172
rect 254762 298160 254768 298172
rect 194652 298132 254768 298160
rect 194652 298120 194658 298132
rect 254762 298120 254768 298132
rect 254820 298120 254826 298172
rect 233694 298052 233700 298104
rect 233752 298092 233758 298104
rect 233970 298092 233976 298104
rect 233752 298064 233976 298092
rect 233752 298052 233758 298064
rect 233970 298052 233976 298064
rect 234028 298052 234034 298104
rect 255958 298052 255964 298104
rect 256016 298092 256022 298104
rect 256326 298092 256332 298104
rect 256016 298064 256332 298092
rect 256016 298052 256022 298064
rect 256326 298052 256332 298064
rect 256384 298052 256390 298104
rect 259270 298052 259276 298104
rect 259328 298092 259334 298104
rect 265710 298092 265716 298104
rect 259328 298064 265716 298092
rect 259328 298052 259334 298064
rect 265710 298052 265716 298064
rect 265768 298052 265774 298104
rect 265820 298024 265848 298268
rect 282822 298052 282828 298104
rect 282880 298092 282886 298104
rect 349062 298092 349068 298104
rect 282880 298064 349068 298092
rect 282880 298052 282886 298064
rect 349062 298052 349068 298064
rect 349120 298052 349126 298104
rect 287146 298024 287152 298036
rect 265820 297996 287152 298024
rect 287146 297984 287152 297996
rect 287204 297984 287210 298036
rect 303246 297984 303252 298036
rect 303304 298024 303310 298036
rect 366174 298024 366180 298036
rect 303304 297996 366180 298024
rect 303304 297984 303310 297996
rect 366174 297984 366180 297996
rect 366232 297984 366238 298036
rect 307938 297916 307944 297968
rect 307996 297956 308002 297968
rect 308490 297956 308496 297968
rect 307996 297928 308496 297956
rect 307996 297916 308002 297928
rect 308490 297916 308496 297928
rect 308548 297916 308554 297968
rect 309042 297916 309048 297968
rect 309100 297956 309106 297968
rect 370222 297956 370228 297968
rect 309100 297928 370228 297956
rect 309100 297916 309106 297928
rect 370222 297916 370228 297928
rect 370280 297916 370286 297968
rect 304718 297848 304724 297900
rect 304776 297888 304782 297900
rect 363414 297888 363420 297900
rect 304776 297860 363420 297888
rect 304776 297848 304782 297860
rect 363414 297848 363420 297860
rect 363472 297848 363478 297900
rect 305454 297780 305460 297832
rect 305512 297820 305518 297832
rect 306098 297820 306104 297832
rect 305512 297792 306104 297820
rect 305512 297780 305518 297792
rect 306098 297780 306104 297792
rect 306156 297820 306162 297832
rect 364794 297820 364800 297832
rect 306156 297792 364800 297820
rect 306156 297780 306162 297792
rect 364794 297780 364800 297792
rect 364852 297780 364858 297832
rect 308490 297712 308496 297764
rect 308548 297752 308554 297764
rect 368198 297752 368204 297764
rect 308548 297724 368204 297752
rect 308548 297712 308554 297724
rect 368198 297712 368204 297724
rect 368256 297712 368262 297764
rect 309042 297644 309048 297696
rect 309100 297684 309106 297696
rect 347222 297684 347228 297696
rect 309100 297656 347228 297684
rect 309100 297644 309106 297656
rect 347222 297644 347228 297656
rect 347280 297644 347286 297696
rect 308950 297576 308956 297628
rect 309008 297616 309014 297628
rect 345750 297616 345756 297628
rect 309008 297588 345756 297616
rect 309008 297576 309014 297588
rect 345750 297576 345756 297588
rect 345808 297576 345814 297628
rect 264054 297440 264060 297492
rect 264112 297480 264118 297492
rect 264238 297480 264244 297492
rect 264112 297452 264244 297480
rect 264112 297440 264118 297452
rect 264238 297440 264244 297452
rect 264296 297440 264302 297492
rect 209130 297372 209136 297424
rect 209188 297412 209194 297424
rect 236638 297412 236644 297424
rect 209188 297384 236644 297412
rect 209188 297372 209194 297384
rect 236638 297372 236644 297384
rect 236696 297372 236702 297424
rect 218790 297304 218796 297356
rect 218848 297344 218854 297356
rect 258718 297344 258724 297356
rect 218848 297316 258724 297344
rect 218848 297304 218854 297316
rect 258718 297304 258724 297316
rect 258776 297304 258782 297356
rect 211798 297236 211804 297288
rect 211856 297276 211862 297288
rect 256326 297276 256332 297288
rect 211856 297248 256332 297276
rect 211856 297236 211862 297248
rect 256326 297236 256332 297248
rect 256384 297236 256390 297288
rect 179414 297168 179420 297220
rect 179472 297208 179478 297220
rect 238110 297208 238116 297220
rect 179472 297180 238116 297208
rect 179472 297168 179478 297180
rect 238110 297168 238116 297180
rect 238168 297168 238174 297220
rect 248598 297168 248604 297220
rect 248656 297208 248662 297220
rect 249058 297208 249064 297220
rect 248656 297180 249064 297208
rect 248656 297168 248662 297180
rect 249058 297168 249064 297180
rect 249116 297168 249122 297220
rect 282086 297168 282092 297220
rect 282144 297208 282150 297220
rect 282822 297208 282828 297220
rect 282144 297180 282828 297208
rect 282144 297168 282150 297180
rect 282822 297168 282828 297180
rect 282880 297168 282886 297220
rect 204438 297100 204444 297152
rect 204496 297140 204502 297152
rect 264330 297140 264336 297152
rect 204496 297112 264336 297140
rect 204496 297100 204502 297112
rect 264330 297100 264336 297112
rect 264388 297100 264394 297152
rect 173894 297032 173900 297084
rect 173952 297072 173958 297084
rect 233694 297072 233700 297084
rect 173952 297044 233700 297072
rect 173952 297032 173958 297044
rect 233694 297032 233700 297044
rect 233752 297032 233758 297084
rect 186314 296964 186320 297016
rect 186372 297004 186378 297016
rect 246390 297004 246396 297016
rect 186372 296976 246396 297004
rect 186372 296964 186378 296976
rect 246390 296964 246396 296976
rect 246448 296964 246454 297016
rect 175274 296896 175280 296948
rect 175332 296936 175338 296948
rect 235350 296936 235356 296948
rect 175332 296908 235356 296936
rect 175332 296896 175338 296908
rect 235350 296896 235356 296908
rect 235408 296896 235414 296948
rect 187694 296828 187700 296880
rect 187752 296868 187758 296880
rect 248598 296868 248604 296880
rect 187752 296840 248604 296868
rect 187752 296828 187758 296840
rect 248598 296828 248604 296840
rect 248656 296828 248662 296880
rect 183554 296760 183560 296812
rect 183612 296800 183618 296812
rect 244550 296800 244556 296812
rect 183612 296772 244556 296800
rect 183612 296760 183618 296772
rect 244550 296760 244556 296772
rect 244608 296800 244614 296812
rect 245010 296800 245016 296812
rect 244608 296772 245016 296800
rect 244608 296760 244614 296772
rect 245010 296760 245016 296772
rect 245068 296760 245074 296812
rect 206646 296692 206652 296744
rect 206704 296732 206710 296744
rect 284570 296732 284576 296744
rect 206704 296704 284576 296732
rect 206704 296692 206710 296704
rect 284570 296692 284576 296704
rect 284628 296692 284634 296744
rect 288710 296624 288716 296676
rect 288768 296664 288774 296676
rect 348970 296664 348976 296676
rect 288768 296636 348976 296664
rect 288768 296624 288774 296636
rect 348970 296624 348976 296636
rect 349028 296624 349034 296676
rect 288342 296556 288348 296608
rect 288400 296596 288406 296608
rect 342990 296596 342996 296608
rect 288400 296568 342996 296596
rect 288400 296556 288406 296568
rect 342990 296556 342996 296568
rect 343048 296556 343054 296608
rect 230566 296148 230572 296200
rect 230624 296188 230630 296200
rect 231210 296188 231216 296200
rect 230624 296160 231216 296188
rect 230624 296148 230630 296160
rect 231210 296148 231216 296160
rect 231268 296148 231274 296200
rect 240042 296080 240048 296132
rect 240100 296120 240106 296132
rect 265986 296120 265992 296132
rect 240100 296092 265992 296120
rect 240100 296080 240106 296092
rect 265986 296080 265992 296092
rect 266044 296080 266050 296132
rect 242802 296012 242808 296064
rect 242860 296052 242866 296064
rect 273162 296052 273168 296064
rect 242860 296024 273168 296052
rect 242860 296012 242866 296024
rect 273162 296012 273168 296024
rect 273220 296012 273226 296064
rect 222286 295944 222292 295996
rect 222344 295984 222350 295996
rect 283558 295984 283564 295996
rect 222344 295956 283564 295984
rect 222344 295944 222350 295956
rect 283558 295944 283564 295956
rect 283616 295944 283622 295996
rect 169754 295876 169760 295928
rect 169812 295916 169818 295928
rect 230566 295916 230572 295928
rect 169812 295888 230572 295916
rect 169812 295876 169818 295888
rect 230566 295876 230572 295888
rect 230624 295876 230630 295928
rect 214742 295808 214748 295860
rect 214800 295848 214806 295860
rect 243354 295848 243360 295860
rect 214800 295820 243360 295848
rect 214800 295808 214806 295820
rect 243354 295808 243360 295820
rect 243412 295808 243418 295860
rect 186958 295740 186964 295792
rect 187016 295780 187022 295792
rect 234890 295780 234896 295792
rect 187016 295752 234896 295780
rect 187016 295740 187022 295752
rect 234890 295740 234896 295752
rect 234948 295740 234954 295792
rect 202138 295672 202144 295724
rect 202196 295712 202202 295724
rect 261662 295712 261668 295724
rect 202196 295684 261668 295712
rect 202196 295672 202202 295684
rect 261662 295672 261668 295684
rect 261720 295672 261726 295724
rect 182174 295604 182180 295656
rect 182232 295644 182238 295656
rect 242158 295644 242164 295656
rect 182232 295616 242164 295644
rect 182232 295604 182238 295616
rect 242158 295604 242164 295616
rect 242216 295604 242222 295656
rect 178034 295536 178040 295588
rect 178092 295576 178098 295588
rect 239030 295576 239036 295588
rect 178092 295548 239036 295576
rect 178092 295536 178098 295548
rect 239030 295536 239036 295548
rect 239088 295576 239094 295588
rect 240042 295576 240048 295588
rect 239088 295548 240048 295576
rect 239088 295536 239094 295548
rect 240042 295536 240048 295548
rect 240100 295536 240106 295588
rect 172514 295468 172520 295520
rect 172572 295508 172578 295520
rect 233510 295508 233516 295520
rect 172572 295480 233516 295508
rect 172572 295468 172578 295480
rect 233510 295468 233516 295480
rect 233568 295508 233574 295520
rect 233878 295508 233884 295520
rect 233568 295480 233884 295508
rect 233568 295468 233574 295480
rect 233878 295468 233884 295480
rect 233936 295468 233942 295520
rect 234982 295468 234988 295520
rect 235040 295508 235046 295520
rect 239398 295508 239404 295520
rect 235040 295480 239404 295508
rect 235040 295468 235046 295480
rect 239398 295468 239404 295480
rect 239456 295468 239462 295520
rect 214650 295400 214656 295452
rect 214708 295440 214714 295452
rect 241974 295440 241980 295452
rect 214708 295412 241980 295440
rect 214708 295400 214714 295412
rect 241974 295400 241980 295412
rect 242032 295440 242038 295452
rect 242802 295440 242808 295452
rect 242032 295412 242808 295440
rect 242032 295400 242038 295412
rect 242802 295400 242808 295412
rect 242860 295400 242866 295452
rect 189074 295332 189080 295384
rect 189132 295372 189138 295384
rect 250530 295372 250536 295384
rect 189132 295344 250536 295372
rect 189132 295332 189138 295344
rect 250530 295332 250536 295344
rect 250588 295332 250594 295384
rect 243078 295264 243084 295316
rect 243136 295304 243142 295316
rect 243354 295304 243360 295316
rect 243136 295276 243360 295304
rect 243136 295264 243142 295276
rect 243354 295264 243360 295276
rect 243412 295304 243418 295316
rect 273070 295304 273076 295316
rect 243412 295276 273076 295304
rect 243412 295264 243418 295276
rect 273070 295264 273076 295276
rect 273128 295264 273134 295316
rect 284018 295264 284024 295316
rect 284076 295304 284082 295316
rect 341518 295304 341524 295316
rect 284076 295276 341524 295304
rect 284076 295264 284082 295276
rect 341518 295264 341524 295276
rect 341576 295264 341582 295316
rect 288618 295196 288624 295248
rect 288676 295236 288682 295248
rect 347038 295236 347044 295248
rect 288676 295208 347044 295236
rect 288676 295196 288682 295208
rect 347038 295196 347044 295208
rect 347096 295196 347102 295248
rect 284570 295128 284576 295180
rect 284628 295168 284634 295180
rect 338850 295168 338856 295180
rect 284628 295140 338856 295168
rect 284628 295128 284634 295140
rect 338850 295128 338856 295140
rect 338908 295128 338914 295180
rect 193214 294788 193220 294840
rect 193272 294828 193278 294840
rect 254486 294828 254492 294840
rect 193272 294800 254492 294828
rect 193272 294788 193278 294800
rect 254486 294788 254492 294800
rect 254544 294788 254550 294840
rect 234246 294720 234252 294772
rect 234304 294760 234310 294772
rect 264606 294760 264612 294772
rect 234304 294732 264612 294760
rect 234304 294720 234310 294732
rect 264606 294720 264612 294732
rect 264664 294720 264670 294772
rect 166994 294652 167000 294704
rect 167052 294692 167058 294704
rect 227990 294692 227996 294704
rect 167052 294664 227996 294692
rect 167052 294652 167058 294664
rect 227990 294652 227996 294664
rect 228048 294692 228054 294704
rect 228450 294692 228456 294704
rect 228048 294664 228456 294692
rect 228048 294652 228054 294664
rect 228450 294652 228456 294664
rect 228508 294652 228514 294704
rect 240042 294652 240048 294704
rect 240100 294692 240106 294704
rect 275186 294692 275192 294704
rect 240100 294664 275192 294692
rect 240100 294652 240106 294664
rect 275186 294652 275192 294664
rect 275244 294652 275250 294704
rect 164510 294584 164516 294636
rect 164568 294624 164574 294636
rect 222010 294624 222016 294636
rect 164568 294596 222016 294624
rect 164568 294584 164574 294596
rect 222010 294584 222016 294596
rect 222068 294584 222074 294636
rect 238386 294584 238392 294636
rect 238444 294624 238450 294636
rect 277946 294624 277952 294636
rect 238444 294596 277952 294624
rect 238444 294584 238450 294596
rect 277946 294584 277952 294596
rect 278004 294584 278010 294636
rect 165890 294516 165896 294568
rect 165948 294556 165954 294568
rect 227070 294556 227076 294568
rect 165948 294528 227076 294556
rect 165948 294516 165954 294528
rect 227070 294516 227076 294528
rect 227128 294516 227134 294568
rect 170398 294448 170404 294500
rect 170456 294488 170462 294500
rect 225690 294488 225696 294500
rect 170456 294460 225696 294488
rect 170456 294448 170462 294460
rect 225690 294448 225696 294460
rect 225748 294448 225754 294500
rect 169846 294380 169852 294432
rect 169904 294420 169910 294432
rect 229830 294420 229836 294432
rect 169904 294392 229836 294420
rect 169904 294380 169910 294392
rect 229830 294380 229836 294392
rect 229888 294420 229894 294432
rect 230198 294420 230204 294432
rect 229888 294392 230204 294420
rect 229888 294380 229894 294392
rect 230198 294380 230204 294392
rect 230256 294380 230262 294432
rect 180794 294312 180800 294364
rect 180852 294352 180858 294364
rect 241606 294352 241612 294364
rect 180852 294324 241612 294352
rect 180852 294312 180858 294324
rect 241606 294312 241612 294324
rect 241664 294312 241670 294364
rect 171134 294244 171140 294296
rect 171192 294284 171198 294296
rect 232406 294284 232412 294296
rect 171192 294256 232412 294284
rect 171192 294244 171198 294256
rect 232406 294244 232412 294256
rect 232464 294244 232470 294296
rect 168374 294176 168380 294228
rect 168432 294216 168438 294228
rect 229094 294216 229100 294228
rect 168432 294188 229100 294216
rect 168432 294176 168438 294188
rect 229094 294176 229100 294188
rect 229152 294216 229158 294228
rect 229370 294216 229376 294228
rect 229152 294188 229376 294216
rect 229152 294176 229158 294188
rect 229370 294176 229376 294188
rect 229428 294176 229434 294228
rect 212074 294108 212080 294160
rect 212132 294148 212138 294160
rect 234246 294148 234252 294160
rect 212132 294120 234252 294148
rect 212132 294108 212138 294120
rect 234246 294108 234252 294120
rect 234304 294108 234310 294160
rect 215018 294040 215024 294092
rect 215076 294080 215082 294092
rect 247034 294080 247040 294092
rect 215076 294052 247040 294080
rect 215076 294040 215082 294052
rect 247034 294040 247040 294052
rect 247092 294040 247098 294092
rect 222010 293972 222016 294024
rect 222068 294012 222074 294024
rect 225046 294012 225052 294024
rect 222068 293984 225052 294012
rect 222068 293972 222074 293984
rect 225046 293972 225052 293984
rect 225104 293972 225110 294024
rect 225690 293972 225696 294024
rect 225748 294012 225754 294024
rect 225966 294012 225972 294024
rect 225748 293984 225972 294012
rect 225748 293972 225754 293984
rect 225966 293972 225972 293984
rect 226024 293972 226030 294024
rect 178126 293632 178132 293684
rect 178184 293672 178190 293684
rect 237374 293672 237380 293684
rect 178184 293644 237380 293672
rect 178184 293632 178190 293644
rect 237374 293632 237380 293644
rect 237432 293632 237438 293684
rect 178218 293564 178224 293616
rect 178276 293604 178282 293616
rect 238386 293604 238392 293616
rect 178276 293576 238392 293604
rect 178276 293564 178282 293576
rect 238386 293564 238392 293576
rect 238444 293564 238450 293616
rect 199654 293496 199660 293548
rect 199712 293536 199718 293548
rect 256970 293536 256976 293548
rect 199712 293508 256976 293536
rect 199712 293496 199718 293508
rect 256970 293496 256976 293508
rect 257028 293536 257034 293548
rect 257338 293536 257344 293548
rect 257028 293508 257344 293536
rect 257028 293496 257034 293508
rect 257338 293496 257344 293508
rect 257396 293496 257402 293548
rect 237466 293360 237472 293412
rect 237524 293400 237530 293412
rect 275830 293400 275836 293412
rect 237524 293372 275836 293400
rect 237524 293360 237530 293372
rect 275830 293360 275836 293372
rect 275888 293360 275894 293412
rect 231946 293292 231952 293344
rect 232004 293332 232010 293344
rect 236454 293332 236460 293344
rect 232004 293304 236460 293332
rect 232004 293292 232010 293304
rect 236454 293292 236460 293304
rect 236512 293332 236518 293344
rect 278590 293332 278596 293344
rect 236512 293304 278596 293332
rect 236512 293292 236518 293304
rect 278590 293292 278596 293304
rect 278648 293292 278654 293344
rect 162670 293224 162676 293276
rect 162728 293264 162734 293276
rect 220354 293264 220360 293276
rect 162728 293236 220360 293264
rect 162728 293224 162734 293236
rect 220354 293224 220360 293236
rect 220412 293264 220418 293276
rect 226518 293264 226524 293276
rect 220412 293236 226524 293264
rect 220412 293224 220418 293236
rect 226518 293224 226524 293236
rect 226576 293224 226582 293276
rect 235350 293224 235356 293276
rect 235408 293264 235414 293276
rect 278130 293264 278136 293276
rect 235408 293236 278136 293264
rect 235408 293224 235414 293236
rect 278130 293224 278136 293236
rect 278188 293224 278194 293276
rect 212258 293156 212264 293208
rect 212316 293196 212322 293208
rect 232038 293196 232044 293208
rect 212316 293168 232044 293196
rect 212316 293156 212322 293168
rect 232038 293156 232044 293168
rect 232096 293156 232102 293208
rect 217226 293088 217232 293140
rect 217284 293128 217290 293140
rect 241882 293128 241888 293140
rect 217284 293100 241888 293128
rect 217284 293088 217290 293100
rect 241882 293088 241888 293100
rect 241940 293088 241946 293140
rect 200758 293020 200764 293072
rect 200816 293060 200822 293072
rect 231946 293060 231952 293072
rect 200816 293032 231952 293060
rect 200816 293020 200822 293032
rect 231946 293020 231952 293032
rect 232004 293020 232010 293072
rect 232038 293020 232044 293072
rect 232096 293060 232102 293072
rect 233142 293060 233148 293072
rect 232096 293032 233148 293060
rect 232096 293020 232102 293032
rect 233142 293020 233148 293032
rect 233200 293020 233206 293072
rect 259638 293020 259644 293072
rect 259696 293060 259702 293072
rect 260190 293060 260196 293072
rect 259696 293032 260196 293060
rect 259696 293020 259702 293032
rect 260190 293020 260196 293032
rect 260248 293020 260254 293072
rect 262306 293020 262312 293072
rect 262364 293060 262370 293072
rect 263134 293060 263140 293072
rect 262364 293032 263140 293060
rect 262364 293020 262370 293032
rect 263134 293020 263140 293032
rect 263192 293020 263198 293072
rect 189718 292952 189724 293004
rect 189776 292992 189782 293004
rect 240042 292992 240048 293004
rect 189776 292964 240048 292992
rect 189776 292952 189782 292964
rect 240042 292952 240048 292964
rect 240100 292952 240106 293004
rect 178678 292884 178684 292936
rect 178736 292924 178742 292936
rect 237466 292924 237472 292936
rect 178736 292896 237472 292924
rect 178736 292884 178742 292896
rect 237466 292884 237472 292896
rect 237524 292884 237530 292936
rect 172606 292816 172612 292868
rect 172664 292856 172670 292868
rect 232774 292856 232780 292868
rect 172664 292828 232780 292856
rect 172664 292816 172670 292828
rect 232774 292816 232780 292828
rect 232832 292856 232838 292868
rect 238018 292856 238024 292868
rect 232832 292828 238024 292856
rect 232832 292816 232838 292828
rect 238018 292816 238024 292828
rect 238076 292816 238082 292868
rect 171226 292748 171232 292800
rect 171284 292788 171290 292800
rect 231118 292788 231124 292800
rect 171284 292760 231124 292788
rect 171284 292748 171290 292760
rect 231118 292748 231124 292760
rect 231176 292788 231182 292800
rect 231302 292788 231308 292800
rect 231176 292760 231308 292788
rect 231176 292748 231182 292760
rect 231302 292748 231308 292760
rect 231360 292748 231366 292800
rect 218514 292680 218520 292732
rect 218572 292720 218578 292732
rect 226978 292720 226984 292732
rect 218572 292692 226984 292720
rect 218572 292680 218578 292692
rect 226978 292680 226984 292692
rect 227036 292680 227042 292732
rect 219250 292612 219256 292664
rect 219308 292652 219314 292664
rect 227714 292652 227720 292664
rect 219308 292624 227720 292652
rect 219308 292612 219314 292624
rect 227714 292612 227720 292624
rect 227772 292612 227778 292664
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 198734 292584 198740 292596
rect 3476 292556 198740 292584
rect 3476 292544 3482 292556
rect 198734 292544 198740 292556
rect 198792 292584 198798 292596
rect 199654 292584 199660 292596
rect 198792 292556 199660 292584
rect 198792 292544 198798 292556
rect 199654 292544 199660 292556
rect 199712 292544 199718 292596
rect 217686 292544 217692 292596
rect 217744 292584 217750 292596
rect 235350 292584 235356 292596
rect 217744 292556 235356 292584
rect 217744 292544 217750 292556
rect 235350 292544 235356 292556
rect 235408 292544 235414 292596
rect 226978 292476 226984 292528
rect 227036 292516 227042 292528
rect 228726 292516 228732 292528
rect 227036 292488 228732 292516
rect 227036 292476 227042 292488
rect 228726 292476 228732 292488
rect 228784 292476 228790 292528
rect 241882 292476 241888 292528
rect 241940 292516 241946 292528
rect 275646 292516 275652 292528
rect 241940 292488 275652 292516
rect 241940 292476 241946 292488
rect 275646 292476 275652 292488
rect 275704 292476 275710 292528
rect 307202 292476 307208 292528
rect 307260 292516 307266 292528
rect 314102 292516 314108 292528
rect 307260 292488 314108 292516
rect 307260 292476 307266 292488
rect 314102 292476 314108 292488
rect 314160 292516 314166 292528
rect 372614 292516 372620 292528
rect 314160 292488 372620 292516
rect 314160 292476 314166 292488
rect 372614 292476 372620 292488
rect 372672 292516 372678 292528
rect 373166 292516 373172 292528
rect 372672 292488 373172 292516
rect 372672 292476 372678 292488
rect 373166 292476 373172 292488
rect 373224 292476 373230 292528
rect 227714 292408 227720 292460
rect 227772 292448 227778 292460
rect 228358 292448 228364 292460
rect 227772 292420 228364 292448
rect 227772 292408 227778 292420
rect 228358 292408 228364 292420
rect 228416 292448 228422 292460
rect 229830 292448 229836 292460
rect 228416 292420 229836 292448
rect 228416 292408 228422 292420
rect 229830 292408 229836 292420
rect 229888 292408 229894 292460
rect 247034 292408 247040 292460
rect 247092 292448 247098 292460
rect 247494 292448 247500 292460
rect 247092 292420 247500 292448
rect 247092 292408 247098 292420
rect 247494 292408 247500 292420
rect 247552 292448 247558 292460
rect 281166 292448 281172 292460
rect 247552 292420 281172 292448
rect 247552 292408 247558 292420
rect 281166 292408 281172 292420
rect 281224 292408 281230 292460
rect 241606 292340 241612 292392
rect 241664 292380 241670 292392
rect 271322 292380 271328 292392
rect 241664 292352 271328 292380
rect 241664 292340 241670 292352
rect 271322 292340 271328 292352
rect 271380 292340 271386 292392
rect 219986 292272 219992 292324
rect 220044 292312 220050 292324
rect 220044 292284 246528 292312
rect 220044 292272 220050 292284
rect 237374 292204 237380 292256
rect 237432 292244 237438 292256
rect 238294 292244 238300 292256
rect 237432 292216 238300 292244
rect 237432 292204 237438 292216
rect 238294 292204 238300 292216
rect 238352 292244 238358 292256
rect 238352 292216 246436 292244
rect 238352 292204 238358 292216
rect 189902 292136 189908 292188
rect 189960 292176 189966 292188
rect 246298 292176 246304 292188
rect 189960 292148 246304 292176
rect 189960 292136 189966 292148
rect 246298 292136 246304 292148
rect 246356 292136 246362 292188
rect 227714 292068 227720 292120
rect 227772 292108 227778 292120
rect 233142 292108 233148 292120
rect 227772 292080 233148 292108
rect 227772 292068 227778 292080
rect 233142 292068 233148 292080
rect 233200 292068 233206 292120
rect 246408 292108 246436 292216
rect 246500 292176 246528 292284
rect 256970 292272 256976 292324
rect 257028 292312 257034 292324
rect 257028 292284 258672 292312
rect 257028 292272 257034 292284
rect 249334 292204 249340 292256
rect 249392 292244 249398 292256
rect 258534 292244 258540 292256
rect 249392 292216 258540 292244
rect 249392 292204 249398 292216
rect 258534 292204 258540 292216
rect 258592 292204 258598 292256
rect 258644 292244 258672 292284
rect 258718 292272 258724 292324
rect 258776 292312 258782 292324
rect 260006 292312 260012 292324
rect 258776 292284 260012 292312
rect 258776 292272 258782 292284
rect 260006 292272 260012 292284
rect 260064 292272 260070 292324
rect 263042 292272 263048 292324
rect 263100 292312 263106 292324
rect 264054 292312 264060 292324
rect 263100 292284 264060 292312
rect 263100 292272 263106 292284
rect 264054 292272 264060 292284
rect 264112 292272 264118 292324
rect 264514 292272 264520 292324
rect 264572 292312 264578 292324
rect 265526 292312 265532 292324
rect 264572 292284 265532 292312
rect 264572 292272 264578 292284
rect 265526 292272 265532 292284
rect 265584 292272 265590 292324
rect 258902 292244 258908 292256
rect 258644 292216 258908 292244
rect 258902 292204 258908 292216
rect 258960 292204 258966 292256
rect 264330 292204 264336 292256
rect 264388 292244 264394 292256
rect 265158 292244 265164 292256
rect 264388 292216 265164 292244
rect 264388 292204 264394 292216
rect 265158 292204 265164 292216
rect 265216 292204 265222 292256
rect 257062 292176 257068 292188
rect 246500 292148 257068 292176
rect 257062 292136 257068 292148
rect 257120 292176 257126 292188
rect 257430 292176 257436 292188
rect 257120 292148 257436 292176
rect 257120 292136 257126 292148
rect 257430 292136 257436 292148
rect 257488 292136 257494 292188
rect 258166 292136 258172 292188
rect 258224 292176 258230 292188
rect 268470 292176 268476 292188
rect 258224 292148 268476 292176
rect 258224 292136 258230 292148
rect 268470 292136 268476 292148
rect 268528 292176 268534 292188
rect 271966 292176 271972 292188
rect 268528 292148 271972 292176
rect 268528 292136 268534 292148
rect 271966 292136 271972 292148
rect 272024 292136 272030 292188
rect 249334 292108 249340 292120
rect 246408 292080 249340 292108
rect 249334 292068 249340 292080
rect 249392 292068 249398 292120
rect 252830 292068 252836 292120
rect 252888 292108 252894 292120
rect 263962 292108 263968 292120
rect 252888 292080 263968 292108
rect 252888 292068 252894 292080
rect 263962 292068 263968 292080
rect 264020 292068 264026 292120
rect 245286 292000 245292 292052
rect 245344 292040 245350 292052
rect 267274 292040 267280 292052
rect 245344 292012 267280 292040
rect 245344 292000 245350 292012
rect 267274 292000 267280 292012
rect 267332 292000 267338 292052
rect 218606 291932 218612 291984
rect 218664 291972 218670 291984
rect 222102 291972 222108 291984
rect 218664 291944 222108 291972
rect 218664 291932 218670 291944
rect 222102 291932 222108 291944
rect 222160 291972 222166 291984
rect 227254 291972 227260 291984
rect 222160 291944 227260 291972
rect 222160 291932 222166 291944
rect 227254 291932 227260 291944
rect 227312 291932 227318 291984
rect 242710 291932 242716 291984
rect 242768 291972 242774 291984
rect 250438 291972 250444 291984
rect 242768 291944 250444 291972
rect 242768 291932 242774 291944
rect 250438 291932 250444 291944
rect 250496 291932 250502 291984
rect 252554 291932 252560 291984
rect 252612 291972 252618 291984
rect 282270 291972 282276 291984
rect 252612 291944 282276 291972
rect 252612 291932 252618 291944
rect 282270 291932 282276 291944
rect 282328 291932 282334 291984
rect 308858 291932 308864 291984
rect 308916 291972 308922 291984
rect 336366 291972 336372 291984
rect 308916 291944 336372 291972
rect 308916 291932 308922 291944
rect 336366 291932 336372 291944
rect 336424 291932 336430 291984
rect 214558 291864 214564 291916
rect 214616 291904 214622 291916
rect 234982 291904 234988 291916
rect 214616 291876 234988 291904
rect 214616 291864 214622 291876
rect 234982 291864 234988 291876
rect 235040 291864 235046 291916
rect 247862 291864 247868 291916
rect 247920 291904 247926 291916
rect 279326 291904 279332 291916
rect 247920 291876 279332 291904
rect 247920 291864 247926 291876
rect 279326 291864 279332 291876
rect 279384 291864 279390 291916
rect 309134 291864 309140 291916
rect 309192 291904 309198 291916
rect 310514 291904 310520 291916
rect 309192 291876 310520 291904
rect 309192 291864 309198 291876
rect 310514 291864 310520 291876
rect 310572 291904 310578 291916
rect 355962 291904 355968 291916
rect 310572 291876 355968 291904
rect 310572 291864 310578 291876
rect 355962 291864 355968 291876
rect 356020 291904 356026 291916
rect 357434 291904 357440 291916
rect 356020 291876 357440 291904
rect 356020 291864 356026 291876
rect 357434 291864 357440 291876
rect 357492 291864 357498 291916
rect 166902 291796 166908 291848
rect 166960 291836 166966 291848
rect 220446 291836 220452 291848
rect 166960 291808 220452 291836
rect 166960 291796 166966 291808
rect 220446 291796 220452 291808
rect 220504 291836 220510 291848
rect 220722 291836 220728 291848
rect 220504 291808 220728 291836
rect 220504 291796 220510 291808
rect 220722 291796 220728 291808
rect 220780 291796 220786 291848
rect 220814 291796 220820 291848
rect 220872 291836 220878 291848
rect 231670 291836 231676 291848
rect 220872 291808 231676 291836
rect 220872 291796 220878 291808
rect 215846 291728 215852 291780
rect 215904 291768 215910 291780
rect 220924 291768 220952 291808
rect 231670 291796 231676 291808
rect 231728 291796 231734 291848
rect 236822 291796 236828 291848
rect 236880 291836 236886 291848
rect 264422 291836 264428 291848
rect 236880 291808 264428 291836
rect 236880 291796 236886 291808
rect 264422 291796 264428 291808
rect 264480 291796 264486 291848
rect 272426 291796 272432 291848
rect 272484 291836 272490 291848
rect 331674 291836 331680 291848
rect 272484 291808 331680 291836
rect 272484 291796 272490 291808
rect 331674 291796 331680 291808
rect 331732 291796 331738 291848
rect 372614 291796 372620 291848
rect 372672 291836 372678 291848
rect 402974 291836 402980 291848
rect 372672 291808 402980 291836
rect 372672 291796 372678 291808
rect 402974 291796 402980 291808
rect 403032 291796 403038 291848
rect 215904 291740 220952 291768
rect 215904 291728 215910 291740
rect 220998 291728 221004 291780
rect 221056 291768 221062 291780
rect 243630 291768 243636 291780
rect 221056 291740 243636 291768
rect 221056 291728 221062 291740
rect 243630 291728 243636 291740
rect 243688 291728 243694 291780
rect 256142 291728 256148 291780
rect 256200 291768 256206 291780
rect 256694 291768 256700 291780
rect 256200 291740 256700 291768
rect 256200 291728 256206 291740
rect 256694 291728 256700 291740
rect 256752 291728 256758 291780
rect 256786 291728 256792 291780
rect 256844 291768 256850 291780
rect 259730 291768 259736 291780
rect 256844 291740 259736 291768
rect 256844 291728 256850 291740
rect 259730 291728 259736 291740
rect 259788 291728 259794 291780
rect 222010 291660 222016 291712
rect 222068 291700 222074 291712
rect 244182 291700 244188 291712
rect 222068 291672 244188 291700
rect 222068 291660 222074 291672
rect 244182 291660 244188 291672
rect 244240 291660 244246 291712
rect 254486 291660 254492 291712
rect 254544 291700 254550 291712
rect 254544 291672 258074 291700
rect 254544 291660 254550 291672
rect 220354 291592 220360 291644
rect 220412 291632 220418 291644
rect 247770 291632 247776 291644
rect 220412 291604 247776 291632
rect 220412 291592 220418 291604
rect 247770 291592 247776 291604
rect 247828 291592 247834 291644
rect 254762 291592 254768 291644
rect 254820 291632 254826 291644
rect 255590 291632 255596 291644
rect 254820 291604 255596 291632
rect 254820 291592 254826 291604
rect 255590 291592 255596 291604
rect 255648 291592 255654 291644
rect 258046 291632 258074 291672
rect 271874 291660 271880 291712
rect 271932 291700 271938 291712
rect 272518 291700 272524 291712
rect 271932 291672 272524 291700
rect 271932 291660 271938 291672
rect 272518 291660 272524 291672
rect 272576 291660 272582 291712
rect 281442 291632 281448 291644
rect 258046 291604 281448 291632
rect 281442 291592 281448 291604
rect 281500 291592 281506 291644
rect 220078 291524 220084 291576
rect 220136 291564 220142 291576
rect 247402 291564 247408 291576
rect 220136 291536 247408 291564
rect 220136 291524 220142 291536
rect 247402 291524 247408 291536
rect 247460 291524 247466 291576
rect 220814 291456 220820 291508
rect 220872 291496 220878 291508
rect 253290 291496 253296 291508
rect 220872 291468 253296 291496
rect 220872 291456 220878 291468
rect 253290 291456 253296 291468
rect 253348 291496 253354 291508
rect 253750 291496 253756 291508
rect 253348 291468 253756 291496
rect 253348 291456 253354 291468
rect 253750 291456 253756 291468
rect 253808 291456 253814 291508
rect 220906 291388 220912 291440
rect 220964 291428 220970 291440
rect 254578 291428 254584 291440
rect 220964 291400 254584 291428
rect 220964 291388 220970 291400
rect 254578 291388 254584 291400
rect 254636 291388 254642 291440
rect 221274 291320 221280 291372
rect 221332 291360 221338 291372
rect 255958 291360 255964 291372
rect 221332 291332 255964 291360
rect 221332 291320 221338 291332
rect 255958 291320 255964 291332
rect 256016 291320 256022 291372
rect 264790 291320 264796 291372
rect 264848 291360 264854 291372
rect 268378 291360 268384 291372
rect 264848 291332 268384 291360
rect 264848 291320 264854 291332
rect 268378 291320 268384 291332
rect 268436 291360 268442 291372
rect 269022 291360 269028 291372
rect 268436 291332 269028 291360
rect 268436 291320 268442 291332
rect 269022 291320 269028 291332
rect 269080 291320 269086 291372
rect 217318 291252 217324 291304
rect 217376 291292 217382 291304
rect 228542 291292 228548 291304
rect 217376 291264 228548 291292
rect 217376 291252 217382 291264
rect 228542 291252 228548 291264
rect 228600 291252 228606 291304
rect 234586 291264 240824 291292
rect 221366 291184 221372 291236
rect 221424 291224 221430 291236
rect 234586 291224 234614 291264
rect 221424 291196 234614 291224
rect 221424 291184 221430 291196
rect 235442 291184 235448 291236
rect 235500 291224 235506 291236
rect 236086 291224 236092 291236
rect 235500 291196 236092 291224
rect 235500 291184 235506 291196
rect 236086 291184 236092 291196
rect 236144 291184 236150 291236
rect 238110 291184 238116 291236
rect 238168 291224 238174 291236
rect 239398 291224 239404 291236
rect 238168 291196 239404 291224
rect 238168 291184 238174 291196
rect 239398 291184 239404 291196
rect 239456 291184 239462 291236
rect 240796 291224 240824 291264
rect 240870 291252 240876 291304
rect 240928 291292 240934 291304
rect 241882 291292 241888 291304
rect 240928 291264 241888 291292
rect 240928 291252 240934 291264
rect 241882 291252 241888 291264
rect 241940 291252 241946 291304
rect 263686 291252 263692 291304
rect 263744 291292 263750 291304
rect 272426 291292 272432 291304
rect 263744 291264 272432 291292
rect 263744 291252 263750 291264
rect 272426 291252 272432 291264
rect 272484 291252 272490 291304
rect 242710 291224 242716 291236
rect 240796 291196 242716 291224
rect 242710 291184 242716 291196
rect 242768 291184 242774 291236
rect 244274 291184 244280 291236
rect 244332 291224 244338 291236
rect 244918 291224 244924 291236
rect 244332 291196 244924 291224
rect 244332 291184 244338 291196
rect 244918 291184 244924 291196
rect 244976 291184 244982 291236
rect 247770 291184 247776 291236
rect 247828 291224 247834 291236
rect 248230 291224 248236 291236
rect 247828 291196 248236 291224
rect 247828 291184 247834 291196
rect 248230 291184 248236 291196
rect 248288 291184 248294 291236
rect 248322 291184 248328 291236
rect 248380 291224 248386 291236
rect 250806 291224 250812 291236
rect 248380 291196 250812 291224
rect 248380 291184 248386 291196
rect 250806 291184 250812 291196
rect 250864 291184 250870 291236
rect 262582 291184 262588 291236
rect 262640 291224 262646 291236
rect 271874 291224 271880 291236
rect 262640 291196 271880 291224
rect 262640 291184 262646 291196
rect 271874 291184 271880 291196
rect 271932 291184 271938 291236
rect 269022 291116 269028 291168
rect 269080 291156 269086 291168
rect 272242 291156 272248 291168
rect 269080 291128 272248 291156
rect 269080 291116 269086 291128
rect 272242 291116 272248 291128
rect 272300 291116 272306 291168
rect 335998 291116 336004 291168
rect 336056 291156 336062 291168
rect 336366 291156 336372 291168
rect 336056 291128 336372 291156
rect 336056 291116 336062 291128
rect 336366 291116 336372 291128
rect 336424 291156 336430 291168
rect 367738 291156 367744 291168
rect 336424 291128 367744 291156
rect 336424 291116 336430 291128
rect 367738 291116 367744 291128
rect 367796 291116 367802 291168
rect 262214 290776 262220 290828
rect 262272 290816 262278 290828
rect 262950 290816 262956 290828
rect 262272 290788 262956 290816
rect 262272 290776 262278 290788
rect 262950 290776 262956 290788
rect 263008 290776 263014 290828
rect 172698 290708 172704 290760
rect 172756 290748 172762 290760
rect 219894 290748 219900 290760
rect 172756 290720 219900 290748
rect 172756 290708 172762 290720
rect 219894 290708 219900 290720
rect 219952 290748 219958 290760
rect 227714 290748 227720 290760
rect 219952 290720 227720 290748
rect 219952 290708 219958 290720
rect 227714 290708 227720 290720
rect 227772 290708 227778 290760
rect 240134 290708 240140 290760
rect 240192 290748 240198 290760
rect 261570 290748 261576 290760
rect 240192 290720 261576 290748
rect 240192 290708 240198 290720
rect 261570 290708 261576 290720
rect 261628 290708 261634 290760
rect 197538 290640 197544 290692
rect 197596 290680 197602 290692
rect 256510 290680 256516 290692
rect 197596 290652 256516 290680
rect 197596 290640 197602 290652
rect 256510 290640 256516 290652
rect 256568 290680 256574 290692
rect 256786 290680 256792 290692
rect 256568 290652 256792 290680
rect 256568 290640 256574 290652
rect 256786 290640 256792 290652
rect 256844 290640 256850 290692
rect 194686 290572 194692 290624
rect 194744 290612 194750 290624
rect 254670 290612 254676 290624
rect 194744 290584 254676 290612
rect 194744 290572 194750 290584
rect 254670 290572 254676 290584
rect 254728 290572 254734 290624
rect 193306 290504 193312 290556
rect 193364 290544 193370 290556
rect 253842 290544 253848 290556
rect 193364 290516 253848 290544
rect 193364 290504 193370 290516
rect 253842 290504 253848 290516
rect 253900 290504 253906 290556
rect 179506 290436 179512 290488
rect 179564 290476 179570 290488
rect 240134 290476 240140 290488
rect 179564 290448 240140 290476
rect 179564 290436 179570 290448
rect 240134 290436 240140 290448
rect 240192 290436 240198 290488
rect 244182 290436 244188 290488
rect 244240 290476 244246 290488
rect 272794 290476 272800 290488
rect 244240 290448 272800 290476
rect 244240 290436 244246 290448
rect 272794 290436 272800 290448
rect 272852 290436 272858 290488
rect 221734 290368 221740 290420
rect 221792 290408 221798 290420
rect 240502 290408 240508 290420
rect 221792 290380 240508 290408
rect 221792 290368 221798 290380
rect 240502 290368 240508 290380
rect 240560 290368 240566 290420
rect 168282 290300 168288 290352
rect 168340 290340 168346 290352
rect 220722 290340 220728 290352
rect 168340 290312 220728 290340
rect 168340 290300 168346 290312
rect 220722 290300 220728 290312
rect 220780 290300 220786 290352
rect 221918 290300 221924 290352
rect 221976 290340 221982 290352
rect 259270 290340 259276 290352
rect 221976 290312 259276 290340
rect 221976 290300 221982 290312
rect 259270 290300 259276 290312
rect 259328 290300 259334 290352
rect 219894 290232 219900 290284
rect 219952 290272 219958 290284
rect 260558 290272 260564 290284
rect 219952 290244 260564 290272
rect 219952 290232 219958 290244
rect 260558 290232 260564 290244
rect 260616 290232 260622 290284
rect 202966 290164 202972 290216
rect 203024 290204 203030 290216
rect 262214 290204 262220 290216
rect 203024 290176 262220 290204
rect 203024 290164 203030 290176
rect 262214 290164 262220 290176
rect 262272 290164 262278 290216
rect 176654 290096 176660 290148
rect 176712 290136 176718 290148
rect 236822 290136 236828 290148
rect 176712 290108 236828 290136
rect 176712 290096 176718 290108
rect 236822 290096 236828 290108
rect 236880 290096 236886 290148
rect 199378 290028 199384 290080
rect 199436 290068 199442 290080
rect 259546 290068 259552 290080
rect 199436 290040 259552 290068
rect 199436 290028 199442 290040
rect 259546 290028 259552 290040
rect 259604 290028 259610 290080
rect 169938 289960 169944 290012
rect 169996 290000 170002 290012
rect 230750 290000 230756 290012
rect 169996 289972 230756 290000
rect 169996 289960 170002 289972
rect 230750 289960 230756 289972
rect 230808 289960 230814 290012
rect 256510 289960 256516 290012
rect 256568 290000 256574 290012
rect 257246 290000 257252 290012
rect 256568 289972 257252 290000
rect 256568 289960 256574 289972
rect 257246 289960 257252 289972
rect 257304 289960 257310 290012
rect 197446 289892 197452 289944
rect 197504 289932 197510 289944
rect 258350 289932 258356 289944
rect 197504 289904 258356 289932
rect 197504 289892 197510 289904
rect 258350 289892 258356 289904
rect 258408 289892 258414 289944
rect 182266 289824 182272 289876
rect 182324 289864 182330 289876
rect 243262 289864 243268 289876
rect 182324 289836 243268 289864
rect 182324 289824 182330 289836
rect 243262 289824 243268 289836
rect 243320 289824 243326 289876
rect 220538 289756 220544 289808
rect 220596 289796 220602 289808
rect 223574 289796 223580 289808
rect 220596 289768 223580 289796
rect 220596 289756 220602 289768
rect 223574 289756 223580 289768
rect 223632 289756 223638 289808
rect 241486 289564 244274 289592
rect 241486 289524 241514 289564
rect 236472 289496 241514 289524
rect 234522 289388 234528 289400
rect 219406 289360 234528 289388
rect 180058 289212 180064 289264
rect 180116 289252 180122 289264
rect 219406 289252 219434 289360
rect 234522 289348 234528 289360
rect 234580 289388 234586 289400
rect 235534 289388 235540 289400
rect 234580 289360 235540 289388
rect 234580 289348 234586 289360
rect 235534 289348 235540 289360
rect 235592 289348 235598 289400
rect 180116 289224 219434 289252
rect 180116 289212 180122 289224
rect 184934 289144 184940 289196
rect 184992 289184 184998 289196
rect 236472 289184 236500 289496
rect 244246 289456 244274 289564
rect 245194 289456 245200 289468
rect 243832 289428 244136 289456
rect 244246 289428 245200 289456
rect 243832 289320 243860 289428
rect 243998 289348 244004 289400
rect 244056 289348 244062 289400
rect 244108 289388 244136 289428
rect 245194 289416 245200 289428
rect 245252 289416 245258 289468
rect 245470 289388 245476 289400
rect 244108 289360 245476 289388
rect 245470 289348 245476 289360
rect 245528 289348 245534 289400
rect 236840 289292 240134 289320
rect 236840 289184 236868 289292
rect 240106 289252 240134 289292
rect 240244 289292 243860 289320
rect 240244 289252 240272 289292
rect 240106 289224 240272 289252
rect 184992 289156 236500 289184
rect 236656 289156 236868 289184
rect 184992 289144 184998 289156
rect 185026 289076 185032 289128
rect 185084 289116 185090 289128
rect 236656 289116 236684 289156
rect 185084 289088 236684 289116
rect 185084 289076 185090 289088
rect 183646 288396 183652 288448
rect 183704 288436 183710 288448
rect 244016 288436 244044 289348
rect 323486 289076 323492 289128
rect 323544 289116 323550 289128
rect 328822 289116 328828 289128
rect 323544 289088 328828 289116
rect 323544 289076 323550 289088
rect 328822 289076 328828 289088
rect 328880 289116 328886 289128
rect 389174 289116 389180 289128
rect 328880 289088 389180 289116
rect 328880 289076 328886 289088
rect 389174 289076 389180 289088
rect 389232 289116 389238 289128
rect 538214 289116 538220 289128
rect 389232 289088 538220 289116
rect 389232 289076 389238 289088
rect 538214 289076 538220 289088
rect 538272 289076 538278 289128
rect 183704 288408 244044 288436
rect 183704 288396 183710 288408
rect 306006 288396 306012 288448
rect 306064 288436 306070 288448
rect 307478 288436 307484 288448
rect 306064 288408 307484 288436
rect 306064 288396 306070 288408
rect 307478 288396 307484 288408
rect 307536 288396 307542 288448
rect 268378 287648 268384 287700
rect 268436 287688 268442 287700
rect 325418 287688 325424 287700
rect 268436 287660 325424 287688
rect 268436 287648 268442 287660
rect 325418 287648 325424 287660
rect 325476 287648 325482 287700
rect 194778 286356 194784 286408
rect 194836 286396 194842 286408
rect 220906 286396 220912 286408
rect 194836 286368 220912 286396
rect 194836 286356 194842 286368
rect 220906 286356 220912 286368
rect 220964 286356 220970 286408
rect 183738 286288 183744 286340
rect 183796 286328 183802 286340
rect 183796 286300 200114 286328
rect 183796 286288 183802 286300
rect 200086 286260 200114 286300
rect 268930 286288 268936 286340
rect 268988 286328 268994 286340
rect 321186 286328 321192 286340
rect 268988 286300 321192 286328
rect 268988 286288 268994 286300
rect 321186 286288 321192 286300
rect 321244 286288 321250 286340
rect 220906 286260 220912 286272
rect 200086 286232 220912 286260
rect 220906 286220 220912 286232
rect 220964 286220 220970 286272
rect 219342 285132 219348 285184
rect 219400 285172 219406 285184
rect 220906 285172 220912 285184
rect 219400 285144 220912 285172
rect 219400 285132 219406 285144
rect 220906 285132 220912 285144
rect 220964 285132 220970 285184
rect 220814 285104 220820 285116
rect 200086 285076 220820 285104
rect 193398 284928 193404 284980
rect 193456 284968 193462 284980
rect 200086 284968 200114 285076
rect 220814 285064 220820 285076
rect 220872 285064 220878 285116
rect 193456 284940 200114 284968
rect 193456 284928 193462 284940
rect 269022 284928 269028 284980
rect 269080 284968 269086 284980
rect 325234 284968 325240 284980
rect 269080 284940 325240 284968
rect 269080 284928 269086 284940
rect 325234 284928 325240 284940
rect 325292 284928 325298 284980
rect 196066 283568 196072 283620
rect 196124 283608 196130 283620
rect 220906 283608 220912 283620
rect 196124 283580 220912 283608
rect 196124 283568 196130 283580
rect 220906 283568 220912 283580
rect 220964 283568 220970 283620
rect 271322 283568 271328 283620
rect 271380 283608 271386 283620
rect 290918 283608 290924 283620
rect 271380 283580 290924 283608
rect 271380 283568 271386 283580
rect 290918 283568 290924 283580
rect 290976 283568 290982 283620
rect 271414 282140 271420 282192
rect 271472 282180 271478 282192
rect 292482 282180 292488 282192
rect 271472 282152 292488 282180
rect 271472 282140 271478 282152
rect 292482 282140 292488 282152
rect 292540 282140 292546 282192
rect 196158 280780 196164 280832
rect 196216 280820 196222 280832
rect 219986 280820 219992 280832
rect 196216 280792 219992 280820
rect 196216 280780 196222 280792
rect 219986 280780 219992 280792
rect 220044 280780 220050 280832
rect 271506 280780 271512 280832
rect 271564 280820 271570 280832
rect 292390 280820 292396 280832
rect 271564 280792 292396 280820
rect 271564 280780 271570 280792
rect 292390 280780 292396 280792
rect 292448 280780 292454 280832
rect 182358 279420 182364 279472
rect 182416 279460 182422 279472
rect 220906 279460 220912 279472
rect 182416 279432 220912 279460
rect 182416 279420 182422 279432
rect 220906 279420 220912 279432
rect 220964 279420 220970 279472
rect 271598 279420 271604 279472
rect 271656 279460 271662 279472
rect 292298 279460 292304 279472
rect 271656 279432 292304 279460
rect 271656 279420 271662 279432
rect 292298 279420 292304 279432
rect 292356 279420 292362 279472
rect 323946 277380 323952 277432
rect 324004 277420 324010 277432
rect 327258 277420 327264 277432
rect 324004 277392 327264 277420
rect 324004 277380 324010 277392
rect 327258 277380 327264 277392
rect 327316 277420 327322 277432
rect 531314 277420 531320 277432
rect 327316 277392 531320 277420
rect 327316 277380 327322 277392
rect 531314 277380 531320 277392
rect 531372 277380 531378 277432
rect 185118 276632 185124 276684
rect 185176 276672 185182 276684
rect 220906 276672 220912 276684
rect 185176 276644 220912 276672
rect 185176 276632 185182 276644
rect 220906 276632 220912 276644
rect 220964 276632 220970 276684
rect 322658 276020 322664 276072
rect 322716 276060 322722 276072
rect 322934 276060 322940 276072
rect 322716 276032 322940 276060
rect 322716 276020 322722 276032
rect 322934 276020 322940 276032
rect 322992 276060 322998 276072
rect 516134 276060 516140 276072
rect 322992 276032 516140 276060
rect 322992 276020 322998 276032
rect 516134 276020 516140 276032
rect 516192 276020 516198 276072
rect 187878 273912 187884 273964
rect 187936 273952 187942 273964
rect 220354 273952 220360 273964
rect 187936 273924 220360 273952
rect 187936 273912 187942 273924
rect 220354 273912 220360 273924
rect 220412 273912 220418 273964
rect 321278 273232 321284 273284
rect 321336 273272 321342 273284
rect 321646 273272 321652 273284
rect 321336 273244 321652 273272
rect 321336 273232 321342 273244
rect 321646 273232 321652 273244
rect 321704 273272 321710 273284
rect 495434 273272 495440 273284
rect 321704 273244 495440 273272
rect 321704 273232 321710 273244
rect 495434 273232 495440 273244
rect 495492 273232 495498 273284
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 14458 266404 14464 266416
rect 3108 266376 14464 266404
rect 3108 266364 3114 266376
rect 14458 266364 14464 266376
rect 14516 266364 14522 266416
rect 325142 266364 325148 266416
rect 325200 266404 325206 266416
rect 325602 266404 325608 266416
rect 325200 266376 325608 266404
rect 325200 266364 325206 266376
rect 325602 266364 325608 266376
rect 325660 266404 325666 266416
rect 542998 266404 543004 266416
rect 325660 266376 543004 266404
rect 325660 266364 325666 266376
rect 542998 266364 543004 266376
rect 543056 266364 543062 266416
rect 317046 264596 317052 264648
rect 317104 264636 317110 264648
rect 317414 264636 317420 264648
rect 317104 264608 317420 264636
rect 317104 264596 317110 264608
rect 317414 264596 317420 264608
rect 317472 264596 317478 264648
rect 314102 263644 314108 263696
rect 314160 263684 314166 263696
rect 314378 263684 314384 263696
rect 314160 263656 314384 263684
rect 314160 263644 314166 263656
rect 314378 263644 314384 263656
rect 314436 263684 314442 263696
rect 414014 263684 414020 263696
rect 314436 263656 414020 263684
rect 314436 263644 314442 263656
rect 414014 263644 414020 263656
rect 414072 263644 414078 263696
rect 317414 263576 317420 263628
rect 317472 263616 317478 263628
rect 445754 263616 445760 263628
rect 317472 263588 445760 263616
rect 317472 263576 317478 263588
rect 445754 263576 445760 263588
rect 445812 263576 445818 263628
rect 312446 262828 312452 262880
rect 312504 262868 312510 262880
rect 347498 262868 347504 262880
rect 312504 262840 347504 262868
rect 312504 262828 312510 262840
rect 347498 262828 347504 262840
rect 347556 262868 347562 262880
rect 389174 262868 389180 262880
rect 347556 262840 389180 262868
rect 347556 262828 347562 262840
rect 389174 262828 389180 262840
rect 389232 262828 389238 262880
rect 318242 262692 318248 262744
rect 318300 262732 318306 262744
rect 318518 262732 318524 262744
rect 318300 262704 318524 262732
rect 318300 262692 318306 262704
rect 318518 262692 318524 262704
rect 318576 262692 318582 262744
rect 318242 262216 318248 262268
rect 318300 262256 318306 262268
rect 452654 262256 452660 262268
rect 318300 262228 452660 262256
rect 318300 262216 318306 262228
rect 452654 262216 452660 262228
rect 452712 262216 452718 262268
rect 295058 260108 295064 260160
rect 295116 260148 295122 260160
rect 322290 260148 322296 260160
rect 295116 260120 322296 260148
rect 295116 260108 295122 260120
rect 322290 260108 322296 260120
rect 322348 260108 322354 260160
rect 310238 259428 310244 259480
rect 310296 259468 310302 259480
rect 360194 259468 360200 259480
rect 310296 259440 360200 259468
rect 310296 259428 310302 259440
rect 360194 259428 360200 259440
rect 360252 259428 360258 259480
rect 316954 258068 316960 258120
rect 317012 258108 317018 258120
rect 441614 258108 441620 258120
rect 317012 258080 441620 258108
rect 317012 258068 317018 258080
rect 441614 258068 441620 258080
rect 441672 258068 441678 258120
rect 269942 257320 269948 257372
rect 270000 257360 270006 257372
rect 313090 257360 313096 257372
rect 270000 257332 313096 257360
rect 270000 257320 270006 257332
rect 313090 257320 313096 257332
rect 313148 257360 313154 257372
rect 391934 257360 391940 257372
rect 313148 257332 391940 257360
rect 313148 257320 313154 257332
rect 391934 257320 391940 257332
rect 391992 257320 391998 257372
rect 319714 256708 319720 256760
rect 319772 256748 319778 256760
rect 470594 256748 470600 256760
rect 319772 256720 470600 256748
rect 319772 256708 319778 256720
rect 470594 256708 470600 256720
rect 470652 256708 470658 256760
rect 315574 255280 315580 255332
rect 315632 255320 315638 255332
rect 315850 255320 315856 255332
rect 315632 255292 315856 255320
rect 315632 255280 315638 255292
rect 315850 255280 315856 255292
rect 315908 255320 315914 255332
rect 427814 255320 427820 255332
rect 315908 255292 427820 255320
rect 315908 255280 315914 255292
rect 427814 255280 427820 255292
rect 427872 255280 427878 255332
rect 268930 254532 268936 254584
rect 268988 254572 268994 254584
rect 290366 254572 290372 254584
rect 268988 254544 290372 254572
rect 268988 254532 268994 254544
rect 290366 254532 290372 254544
rect 290424 254532 290430 254584
rect 311526 253988 311532 254040
rect 311584 254028 311590 254040
rect 364334 254028 364340 254040
rect 311584 254000 364340 254028
rect 311584 253988 311590 254000
rect 364334 253988 364340 254000
rect 364392 253988 364398 254040
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 3476 253932 200114 253960
rect 3476 253920 3482 253932
rect 200086 253892 200114 253932
rect 323762 253920 323768 253972
rect 323820 253960 323826 253972
rect 527174 253960 527180 253972
rect 323820 253932 527180 253960
rect 323820 253920 323826 253932
rect 527174 253920 527180 253932
rect 527232 253920 527238 253972
rect 200206 253892 200212 253904
rect 200086 253864 200212 253892
rect 200206 253852 200212 253864
rect 200264 253892 200270 253904
rect 216030 253892 216036 253904
rect 200264 253864 216036 253892
rect 200264 253852 200270 253864
rect 216030 253852 216036 253864
rect 216088 253852 216094 253904
rect 275646 253172 275652 253224
rect 275704 253212 275710 253224
rect 321094 253212 321100 253224
rect 275704 253184 321100 253212
rect 275704 253172 275710 253184
rect 321094 253172 321100 253184
rect 321152 253172 321158 253224
rect 316770 253036 316776 253088
rect 316828 253076 316834 253088
rect 317230 253076 317236 253088
rect 316828 253048 317236 253076
rect 316828 253036 316834 253048
rect 317230 253036 317236 253048
rect 317288 253036 317294 253088
rect 310330 252696 310336 252748
rect 310388 252736 310394 252748
rect 349246 252736 349252 252748
rect 310388 252708 349252 252736
rect 310388 252696 310394 252708
rect 349246 252696 349252 252708
rect 349304 252696 349310 252748
rect 317230 252628 317236 252680
rect 317288 252668 317294 252680
rect 448606 252668 448612 252680
rect 317288 252640 448612 252668
rect 317288 252628 317294 252640
rect 448606 252628 448612 252640
rect 448664 252628 448670 252680
rect 323854 252560 323860 252612
rect 323912 252600 323918 252612
rect 324130 252600 324136 252612
rect 323912 252572 324136 252600
rect 323912 252560 323918 252572
rect 324130 252560 324136 252572
rect 324188 252600 324194 252612
rect 523126 252600 523132 252612
rect 324188 252572 523132 252600
rect 324188 252560 324194 252572
rect 523126 252560 523132 252572
rect 523184 252560 523190 252612
rect 268930 251812 268936 251864
rect 268988 251852 268994 251864
rect 290642 251852 290648 251864
rect 268988 251824 290648 251852
rect 268988 251812 268994 251824
rect 290642 251812 290648 251824
rect 290700 251812 290706 251864
rect 214926 251608 214932 251660
rect 214984 251648 214990 251660
rect 215662 251648 215668 251660
rect 214984 251620 215668 251648
rect 214984 251608 214990 251620
rect 215662 251608 215668 251620
rect 215720 251608 215726 251660
rect 315666 251268 315672 251320
rect 315724 251308 315730 251320
rect 315942 251308 315948 251320
rect 315724 251280 315948 251308
rect 315724 251268 315730 251280
rect 315942 251268 315948 251280
rect 316000 251308 316006 251320
rect 423766 251308 423772 251320
rect 316000 251280 423772 251308
rect 316000 251268 316006 251280
rect 423766 251268 423772 251280
rect 423824 251268 423830 251320
rect 321370 251200 321376 251252
rect 321428 251240 321434 251252
rect 491294 251240 491300 251252
rect 321428 251212 491300 251240
rect 321428 251200 321434 251212
rect 491294 251200 491300 251212
rect 491352 251200 491358 251252
rect 271782 250452 271788 250504
rect 271840 250492 271846 250504
rect 317138 250492 317144 250504
rect 271840 250464 317144 250492
rect 271840 250452 271846 250464
rect 317138 250452 317144 250464
rect 317196 250492 317202 250504
rect 438854 250492 438860 250504
rect 317196 250464 438860 250492
rect 317196 250452 317202 250464
rect 438854 250452 438860 250464
rect 438912 250452 438918 250504
rect 323026 249772 323032 249824
rect 323084 249812 323090 249824
rect 324222 249812 324228 249824
rect 323084 249784 324228 249812
rect 323084 249772 323090 249784
rect 324222 249772 324228 249784
rect 324280 249812 324286 249824
rect 534074 249812 534080 249824
rect 324280 249784 534080 249812
rect 324280 249772 324286 249784
rect 534074 249772 534080 249784
rect 534132 249772 534138 249824
rect 307478 249704 307484 249756
rect 307536 249744 307542 249756
rect 308674 249744 308680 249756
rect 307536 249716 308680 249744
rect 307536 249704 307542 249716
rect 308674 249704 308680 249716
rect 308732 249704 308738 249756
rect 314194 249704 314200 249756
rect 314252 249744 314258 249756
rect 314562 249744 314568 249756
rect 314252 249716 314568 249744
rect 314252 249704 314258 249716
rect 314562 249704 314568 249716
rect 314620 249704 314626 249756
rect 292298 249092 292304 249144
rect 292356 249132 292362 249144
rect 316678 249132 316684 249144
rect 292356 249104 316684 249132
rect 292356 249092 292362 249104
rect 316678 249092 316684 249104
rect 316736 249092 316742 249144
rect 171318 249024 171324 249076
rect 171376 249064 171382 249076
rect 215846 249064 215852 249076
rect 171376 249036 215852 249064
rect 171376 249024 171382 249036
rect 215846 249024 215852 249036
rect 215904 249024 215910 249076
rect 273070 249024 273076 249076
rect 273128 249064 273134 249076
rect 323026 249064 323032 249076
rect 273128 249036 323032 249064
rect 273128 249024 273134 249036
rect 323026 249024 323032 249036
rect 323084 249024 323090 249076
rect 312906 248480 312912 248532
rect 312964 248520 312970 248532
rect 382274 248520 382280 248532
rect 312964 248492 382280 248520
rect 312964 248480 312970 248492
rect 382274 248480 382280 248492
rect 382332 248480 382338 248532
rect 314194 248412 314200 248464
rect 314252 248452 314258 248464
rect 407114 248452 407120 248464
rect 314252 248424 407120 248452
rect 314252 248412 314258 248424
rect 407114 248412 407120 248424
rect 407172 248412 407178 248464
rect 168466 247664 168472 247716
rect 168524 247704 168530 247716
rect 217134 247704 217140 247716
rect 168524 247676 217140 247704
rect 168524 247664 168530 247676
rect 217134 247664 217140 247676
rect 217192 247664 217198 247716
rect 281994 247664 282000 247716
rect 282052 247704 282058 247716
rect 307386 247704 307392 247716
rect 282052 247676 307392 247704
rect 282052 247664 282058 247676
rect 307386 247664 307392 247676
rect 307444 247664 307450 247716
rect 314286 247120 314292 247172
rect 314344 247160 314350 247172
rect 409874 247160 409880 247172
rect 314344 247132 409880 247160
rect 314344 247120 314350 247132
rect 409874 247120 409880 247132
rect 409932 247120 409938 247172
rect 318150 247052 318156 247104
rect 318208 247092 318214 247104
rect 318610 247092 318616 247104
rect 318208 247064 318616 247092
rect 318208 247052 318214 247064
rect 318610 247052 318616 247064
rect 318668 247092 318674 247104
rect 459554 247092 459560 247104
rect 318668 247064 459560 247092
rect 318668 247052 318674 247064
rect 459554 247052 459560 247064
rect 459612 247052 459618 247104
rect 168558 246304 168564 246356
rect 168616 246344 168622 246356
rect 217318 246344 217324 246356
rect 168616 246316 217324 246344
rect 168616 246304 168622 246316
rect 217318 246304 217324 246316
rect 217376 246304 217382 246356
rect 269298 246304 269304 246356
rect 269356 246344 269362 246356
rect 292114 246344 292120 246356
rect 269356 246316 292120 246344
rect 269356 246304 269362 246316
rect 292114 246304 292120 246316
rect 292172 246304 292178 246356
rect 310422 245828 310428 245880
rect 310480 245868 310486 245880
rect 310480 245840 316034 245868
rect 310480 245828 310486 245840
rect 316006 245732 316034 245840
rect 353294 245732 353300 245744
rect 316006 245704 353300 245732
rect 353294 245692 353300 245704
rect 353352 245692 353358 245744
rect 310054 245624 310060 245676
rect 310112 245664 310118 245676
rect 310422 245664 310428 245676
rect 310112 245636 310428 245664
rect 310112 245624 310118 245636
rect 310422 245624 310428 245636
rect 310480 245624 310486 245676
rect 316678 245624 316684 245676
rect 316736 245664 316742 245676
rect 317322 245664 317328 245676
rect 316736 245636 317328 245664
rect 316736 245624 316742 245636
rect 317322 245624 317328 245636
rect 317380 245664 317386 245676
rect 434714 245664 434720 245676
rect 317380 245636 434720 245664
rect 317380 245624 317386 245636
rect 434714 245624 434720 245636
rect 434772 245624 434778 245676
rect 577498 245556 577504 245608
rect 577556 245596 577562 245608
rect 579614 245596 579620 245608
rect 577556 245568 579620 245596
rect 577556 245556 577562 245568
rect 579614 245556 579620 245568
rect 579672 245556 579678 245608
rect 287606 244944 287612 244996
rect 287664 244984 287670 244996
rect 312722 244984 312728 244996
rect 287664 244956 312728 244984
rect 287664 244944 287670 244956
rect 312722 244944 312728 244956
rect 312780 244944 312786 244996
rect 167086 244876 167092 244928
rect 167144 244916 167150 244928
rect 218606 244916 218612 244928
rect 167144 244888 218612 244916
rect 167144 244876 167150 244888
rect 218606 244876 218612 244888
rect 218664 244876 218670 244928
rect 285858 244876 285864 244928
rect 285916 244916 285922 244928
rect 314010 244916 314016 244928
rect 285916 244888 314016 244916
rect 285916 244876 285922 244888
rect 314010 244876 314016 244888
rect 314068 244876 314074 244928
rect 312354 244400 312360 244452
rect 312412 244440 312418 244452
rect 312906 244440 312912 244452
rect 312412 244412 312912 244440
rect 312412 244400 312418 244412
rect 312906 244400 312912 244412
rect 312964 244440 312970 244452
rect 385034 244440 385040 244452
rect 312964 244412 385040 244440
rect 312964 244400 312970 244412
rect 385034 244400 385040 244412
rect 385092 244400 385098 244452
rect 318334 244332 318340 244384
rect 318392 244372 318398 244384
rect 456794 244372 456800 244384
rect 318392 244344 456800 244372
rect 318392 244332 318398 244344
rect 456794 244332 456800 244344
rect 456852 244332 456858 244384
rect 321554 244264 321560 244316
rect 321612 244304 321618 244316
rect 322750 244304 322756 244316
rect 321612 244276 322756 244304
rect 321612 244264 321618 244276
rect 322750 244264 322756 244276
rect 322808 244304 322814 244316
rect 507118 244304 507124 244316
rect 322808 244276 507124 244304
rect 322808 244264 322814 244276
rect 507118 244264 507124 244276
rect 507176 244264 507182 244316
rect 288526 243720 288532 243772
rect 288584 243760 288590 243772
rect 288584 243732 296714 243760
rect 288584 243720 288590 243732
rect 270586 243652 270592 243704
rect 270644 243692 270650 243704
rect 288894 243692 288900 243704
rect 270644 243664 288900 243692
rect 270644 243652 270650 243664
rect 288894 243652 288900 243664
rect 288952 243652 288958 243704
rect 296686 243692 296714 243732
rect 313918 243692 313924 243704
rect 296686 243664 313924 243692
rect 313918 243652 313924 243664
rect 313976 243652 313982 243704
rect 273346 243584 273352 243636
rect 273404 243624 273410 243636
rect 315482 243624 315488 243636
rect 273404 243596 315488 243624
rect 273404 243584 273410 243596
rect 315482 243584 315488 243596
rect 315540 243584 315546 243636
rect 191926 243516 191932 243568
rect 191984 243556 191990 243568
rect 218698 243556 218704 243568
rect 191984 243528 218704 243556
rect 191984 243516 191990 243528
rect 218698 243516 218704 243528
rect 218756 243516 218762 243568
rect 274910 243516 274916 243568
rect 274968 243556 274974 243568
rect 321554 243556 321560 243568
rect 274968 243528 321560 243556
rect 274968 243516 274974 243528
rect 321554 243516 321560 243528
rect 321612 243516 321618 243568
rect 210510 243448 210516 243500
rect 210568 243488 210574 243500
rect 213822 243488 213828 243500
rect 210568 243460 213828 243488
rect 210568 243448 210574 243460
rect 213822 243448 213828 243460
rect 213880 243448 213886 243500
rect 320082 242972 320088 243024
rect 320140 243012 320146 243024
rect 471238 243012 471244 243024
rect 320140 242984 471244 243012
rect 320140 242972 320146 242984
rect 471238 242972 471244 242984
rect 471296 242972 471302 243024
rect 321554 242904 321560 242956
rect 321612 242944 321618 242956
rect 322842 242944 322848 242956
rect 321612 242916 322848 242944
rect 321612 242904 321618 242916
rect 322842 242904 322848 242916
rect 322900 242944 322906 242956
rect 520274 242944 520280 242956
rect 322900 242916 520280 242944
rect 322900 242904 322906 242916
rect 520274 242904 520280 242916
rect 520332 242904 520338 242956
rect 313918 242496 313924 242548
rect 313976 242536 313982 242548
rect 315390 242536 315396 242548
rect 313976 242508 315396 242536
rect 313976 242496 313982 242508
rect 315390 242496 315396 242508
rect 315448 242496 315454 242548
rect 268930 242360 268936 242412
rect 268988 242400 268994 242412
rect 271230 242400 271236 242412
rect 268988 242372 271236 242400
rect 268988 242360 268994 242372
rect 271230 242360 271236 242372
rect 271288 242360 271294 242412
rect 284846 242292 284852 242344
rect 284904 242332 284910 242344
rect 309870 242332 309876 242344
rect 284904 242304 309876 242332
rect 284904 242292 284910 242304
rect 309870 242292 309876 242304
rect 309928 242292 309934 242344
rect 271230 242224 271236 242276
rect 271288 242264 271294 242276
rect 277486 242264 277492 242276
rect 271288 242236 277492 242264
rect 271288 242224 271294 242236
rect 277486 242224 277492 242236
rect 277544 242264 277550 242276
rect 321554 242264 321560 242276
rect 277544 242236 321560 242264
rect 277544 242224 277550 242236
rect 321554 242224 321560 242236
rect 321612 242224 321618 242276
rect 173986 242156 173992 242208
rect 174044 242196 174050 242208
rect 214558 242196 214564 242208
rect 174044 242168 214564 242196
rect 174044 242156 174050 242168
rect 214558 242156 214564 242168
rect 214616 242156 214622 242208
rect 269206 242156 269212 242208
rect 269264 242196 269270 242208
rect 276106 242196 276112 242208
rect 269264 242168 276112 242196
rect 269264 242156 269270 242168
rect 276106 242156 276112 242168
rect 276164 242196 276170 242208
rect 324958 242196 324964 242208
rect 276164 242168 324964 242196
rect 276164 242156 276170 242168
rect 324958 242156 324964 242168
rect 325016 242156 325022 242208
rect 268286 242020 268292 242072
rect 268344 242060 268350 242072
rect 271598 242060 271604 242072
rect 268344 242032 271604 242060
rect 268344 242020 268350 242032
rect 271598 242020 271604 242032
rect 271656 242020 271662 242072
rect 274542 241884 274548 241936
rect 274600 241924 274606 241936
rect 275922 241924 275928 241936
rect 274600 241896 275928 241924
rect 274600 241884 274606 241896
rect 275922 241884 275928 241896
rect 275980 241884 275986 241936
rect 160002 241612 160008 241664
rect 160060 241652 160066 241664
rect 204898 241652 204904 241664
rect 160060 241624 204904 241652
rect 160060 241612 160066 241624
rect 204898 241612 204904 241624
rect 204956 241652 204962 241664
rect 221182 241652 221188 241664
rect 204956 241624 221188 241652
rect 204956 241612 204962 241624
rect 221182 241612 221188 241624
rect 221240 241612 221246 241664
rect 269390 241612 269396 241664
rect 269448 241652 269454 241664
rect 271322 241652 271328 241664
rect 269448 241624 271328 241652
rect 269448 241612 269454 241624
rect 271322 241612 271328 241624
rect 271380 241612 271386 241664
rect 157242 241544 157248 241596
rect 157300 241584 157306 241596
rect 206370 241584 206376 241596
rect 157300 241556 206376 241584
rect 157300 241544 157306 241556
rect 206370 241544 206376 241556
rect 206428 241544 206434 241596
rect 207658 241544 207664 241596
rect 207716 241584 207722 241596
rect 222286 241584 222292 241596
rect 207716 241556 222292 241584
rect 207716 241544 207722 241556
rect 222286 241544 222292 241556
rect 222344 241544 222350 241596
rect 269482 241544 269488 241596
rect 269540 241584 269546 241596
rect 271506 241584 271512 241596
rect 269540 241556 271512 241584
rect 269540 241544 269546 241556
rect 271506 241544 271512 241556
rect 271564 241544 271570 241596
rect 274634 241544 274640 241596
rect 274692 241584 274698 241596
rect 275646 241584 275652 241596
rect 274692 241556 275652 241584
rect 274692 241544 274698 241556
rect 275646 241544 275652 241556
rect 275704 241544 275710 241596
rect 320082 241544 320088 241596
rect 320140 241584 320146 241596
rect 481634 241584 481640 241596
rect 320140 241556 481640 241584
rect 320140 241544 320146 241556
rect 481634 241544 481640 241556
rect 481692 241544 481698 241596
rect 154298 241476 154304 241528
rect 154356 241516 154362 241528
rect 209222 241516 209228 241528
rect 154356 241488 209228 241516
rect 154356 241476 154362 241488
rect 209222 241476 209228 241488
rect 209280 241476 209286 241528
rect 215662 241476 215668 241528
rect 215720 241516 215726 241528
rect 215720 241488 234246 241516
rect 215720 241476 215726 241488
rect 14458 241408 14464 241460
rect 14516 241448 14522 241460
rect 198826 241448 198832 241460
rect 14516 241420 198832 241448
rect 14516 241408 14522 241420
rect 198826 241408 198832 241420
rect 198884 241448 198890 241460
rect 199378 241448 199384 241460
rect 198884 241420 199384 241448
rect 198884 241408 198890 241420
rect 199378 241408 199384 241420
rect 199436 241408 199442 241460
rect 219986 241408 219992 241460
rect 220044 241448 220050 241460
rect 220170 241448 220176 241460
rect 220044 241420 220176 241448
rect 220044 241408 220050 241420
rect 220170 241408 220176 241420
rect 220228 241408 220234 241460
rect 221366 241408 221372 241460
rect 221424 241448 221430 241460
rect 221424 241420 233786 241448
rect 221424 241408 221430 241420
rect 216122 241272 216128 241324
rect 216180 241312 216186 241324
rect 221366 241312 221372 241324
rect 216180 241284 221372 241312
rect 216180 241272 216186 241284
rect 221366 241272 221372 241284
rect 221424 241272 221430 241324
rect 214834 241136 214840 241188
rect 214892 241176 214898 241188
rect 214892 241148 230612 241176
rect 214892 241136 214898 241148
rect 219066 241068 219072 241120
rect 219124 241108 219130 241120
rect 220814 241108 220820 241120
rect 219124 241080 220820 241108
rect 219124 241068 219130 241080
rect 220814 241068 220820 241080
rect 220872 241068 220878 241120
rect 213914 241000 213920 241052
rect 213972 241040 213978 241052
rect 213972 241012 230152 241040
rect 213972 241000 213978 241012
rect 220262 240864 220268 240916
rect 220320 240904 220326 240916
rect 220320 240876 229968 240904
rect 220320 240864 220326 240876
rect 218882 240796 218888 240848
rect 218940 240836 218946 240848
rect 218940 240808 229830 240836
rect 218940 240796 218946 240808
rect 189166 240728 189172 240780
rect 189224 240768 189230 240780
rect 220170 240768 220176 240780
rect 189224 240740 220176 240768
rect 189224 240728 189230 240740
rect 220170 240728 220176 240740
rect 220228 240728 220234 240780
rect 220354 240728 220360 240780
rect 220412 240768 220418 240780
rect 220412 240740 228864 240768
rect 220412 240728 220418 240740
rect 206646 240660 206652 240712
rect 206704 240700 206710 240712
rect 222010 240700 222016 240712
rect 206704 240672 222016 240700
rect 206704 240660 206710 240672
rect 222010 240660 222016 240672
rect 222068 240660 222074 240712
rect 219526 240592 219532 240644
rect 219584 240632 219590 240644
rect 219584 240604 224724 240632
rect 219584 240592 219590 240604
rect 215846 240524 215852 240576
rect 215904 240564 215910 240576
rect 216398 240564 216404 240576
rect 215904 240536 216404 240564
rect 215904 240524 215910 240536
rect 216398 240524 216404 240536
rect 216456 240524 216462 240576
rect 224696 240564 224724 240604
rect 224696 240536 225138 240564
rect 213730 240456 213736 240508
rect 213788 240496 213794 240508
rect 225110 240496 225138 240536
rect 228836 240496 228864 240740
rect 213788 240468 225046 240496
rect 225110 240468 225414 240496
rect 228836 240468 229462 240496
rect 213788 240456 213794 240468
rect 225018 240428 225046 240468
rect 225018 240400 225138 240428
rect 214466 240320 214472 240372
rect 214524 240360 214530 240372
rect 216122 240360 216128 240372
rect 214524 240332 216128 240360
rect 214524 240320 214530 240332
rect 216122 240320 216128 240332
rect 216180 240320 216186 240372
rect 206370 240252 206376 240304
rect 206428 240292 206434 240304
rect 206428 240264 224862 240292
rect 206428 240252 206434 240264
rect 213178 240184 213184 240236
rect 213236 240224 213242 240236
rect 214834 240224 214840 240236
rect 213236 240196 214840 240224
rect 213236 240184 213242 240196
rect 214834 240184 214840 240196
rect 214892 240184 214898 240236
rect 216030 240184 216036 240236
rect 216088 240224 216094 240236
rect 219066 240224 219072 240236
rect 216088 240196 219072 240224
rect 216088 240184 216094 240196
rect 219066 240184 219072 240196
rect 219124 240184 219130 240236
rect 219342 240184 219348 240236
rect 219400 240224 219406 240236
rect 219400 240196 223666 240224
rect 219400 240184 219406 240196
rect 217870 240048 217876 240100
rect 217928 240088 217934 240100
rect 219526 240088 219532 240100
rect 217928 240060 219532 240088
rect 217928 240048 217934 240060
rect 219526 240048 219532 240060
rect 219584 240048 219590 240100
rect 222286 240048 222292 240100
rect 222344 240088 222350 240100
rect 222344 240060 223574 240088
rect 222344 240048 222350 240060
rect 217962 239980 217968 240032
rect 218020 240020 218026 240032
rect 222102 240020 222108 240032
rect 218020 239992 222108 240020
rect 218020 239980 218026 239992
rect 222102 239980 222108 239992
rect 222160 240020 222166 240032
rect 222160 239992 222654 240020
rect 222160 239980 222166 239992
rect 222626 239964 222654 239992
rect 223270 239992 223390 240020
rect 215202 239912 215208 239964
rect 215260 239952 215266 239964
rect 222516 239952 222522 239964
rect 215260 239924 222522 239952
rect 215260 239912 215266 239924
rect 222516 239912 222522 239924
rect 222574 239912 222580 239964
rect 222608 239912 222614 239964
rect 222666 239912 222672 239964
rect 222700 239912 222706 239964
rect 222758 239912 222764 239964
rect 223068 239952 223074 239964
rect 222810 239924 223074 239952
rect 210418 239844 210424 239896
rect 210476 239884 210482 239896
rect 221274 239884 221280 239896
rect 210476 239856 221280 239884
rect 210476 239844 210482 239856
rect 221274 239844 221280 239856
rect 221332 239844 221338 239896
rect 221550 239844 221556 239896
rect 221608 239884 221614 239896
rect 222378 239884 222384 239896
rect 221608 239856 222384 239884
rect 221608 239844 221614 239856
rect 222378 239844 222384 239856
rect 222436 239884 222442 239896
rect 222718 239884 222746 239912
rect 222436 239856 222746 239884
rect 222436 239844 222442 239856
rect 216674 239776 216680 239828
rect 216732 239816 216738 239828
rect 222810 239816 222838 239924
rect 223068 239912 223074 239924
rect 223126 239912 223132 239964
rect 223160 239912 223166 239964
rect 223218 239912 223224 239964
rect 222884 239844 222890 239896
rect 222942 239884 222948 239896
rect 222942 239844 222976 239884
rect 216732 239788 222838 239816
rect 216732 239776 216738 239788
rect 163498 239708 163504 239760
rect 163556 239748 163562 239760
rect 222838 239748 222844 239760
rect 163556 239720 222844 239748
rect 163556 239708 163562 239720
rect 222838 239708 222844 239720
rect 222896 239708 222902 239760
rect 198918 239640 198924 239692
rect 198976 239680 198982 239692
rect 218790 239680 218796 239692
rect 198976 239652 218796 239680
rect 198976 239640 198982 239652
rect 218790 239640 218796 239652
rect 218848 239640 218854 239692
rect 218974 239640 218980 239692
rect 219032 239680 219038 239692
rect 222194 239680 222200 239692
rect 219032 239652 222200 239680
rect 219032 239640 219038 239652
rect 222194 239640 222200 239652
rect 222252 239680 222258 239692
rect 222948 239680 222976 239844
rect 223178 239828 223206 239912
rect 223114 239776 223120 239828
rect 223172 239788 223206 239828
rect 223172 239776 223178 239788
rect 222252 239652 222976 239680
rect 222252 239640 222258 239652
rect 186498 239572 186504 239624
rect 186556 239612 186562 239624
rect 220078 239612 220084 239624
rect 186556 239584 220084 239612
rect 186556 239572 186562 239584
rect 220078 239572 220084 239584
rect 220136 239572 220142 239624
rect 221090 239572 221096 239624
rect 221148 239612 221154 239624
rect 223270 239612 223298 239992
rect 223362 239964 223390 239992
rect 223546 239964 223574 240060
rect 223638 240020 223666 240196
rect 224834 240156 224862 240264
rect 224834 240128 225046 240156
rect 223638 239992 224034 240020
rect 223344 239912 223350 239964
rect 223402 239912 223408 239964
rect 223436 239912 223442 239964
rect 223494 239912 223500 239964
rect 223528 239912 223534 239964
rect 223586 239912 223592 239964
rect 223620 239912 223626 239964
rect 223678 239912 223684 239964
rect 223712 239912 223718 239964
rect 223770 239912 223776 239964
rect 223896 239912 223902 239964
rect 223954 239912 223960 239964
rect 223454 239884 223482 239912
rect 223408 239856 223482 239884
rect 223408 239760 223436 239856
rect 223638 239828 223666 239912
rect 223730 239884 223758 239912
rect 223730 239856 223804 239884
rect 223638 239788 223672 239828
rect 223666 239776 223672 239788
rect 223724 239776 223730 239828
rect 223390 239708 223396 239760
rect 223448 239708 223454 239760
rect 223482 239708 223488 239760
rect 223540 239748 223546 239760
rect 223776 239748 223804 239856
rect 223540 239720 223804 239748
rect 223540 239708 223546 239720
rect 223666 239640 223672 239692
rect 223724 239680 223730 239692
rect 223914 239680 223942 239912
rect 223724 239652 223942 239680
rect 223724 239640 223730 239652
rect 221148 239584 223298 239612
rect 221148 239572 221154 239584
rect 159726 239504 159732 239556
rect 159784 239544 159790 239556
rect 205082 239544 205088 239556
rect 159784 239516 205088 239544
rect 159784 239504 159790 239516
rect 205082 239504 205088 239516
rect 205140 239544 205146 239556
rect 205450 239544 205456 239556
rect 205140 239516 205456 239544
rect 205140 239504 205146 239516
rect 205450 239504 205456 239516
rect 205508 239504 205514 239556
rect 215110 239504 215116 239556
rect 215168 239544 215174 239556
rect 224006 239544 224034 239992
rect 225018 239964 225046 240128
rect 224172 239912 224178 239964
rect 224230 239912 224236 239964
rect 224264 239912 224270 239964
rect 224322 239912 224328 239964
rect 224356 239912 224362 239964
rect 224414 239952 224420 239964
rect 224414 239912 224448 239952
rect 224632 239912 224638 239964
rect 224690 239912 224696 239964
rect 224816 239912 224822 239964
rect 224874 239912 224880 239964
rect 224908 239912 224914 239964
rect 224966 239912 224972 239964
rect 225000 239912 225006 239964
rect 225058 239912 225064 239964
rect 224080 239844 224086 239896
rect 224138 239844 224144 239896
rect 224098 239624 224126 239844
rect 224190 239828 224218 239912
rect 224282 239884 224310 239912
rect 224282 239856 224356 239884
rect 224328 239828 224356 239856
rect 224190 239788 224224 239828
rect 224218 239776 224224 239788
rect 224276 239776 224282 239828
rect 224310 239776 224316 239828
rect 224368 239776 224374 239828
rect 224098 239584 224132 239624
rect 224126 239572 224132 239584
rect 224184 239572 224190 239624
rect 224420 239612 224448 239912
rect 224540 239884 224546 239896
rect 224512 239844 224546 239884
rect 224598 239844 224604 239896
rect 224512 239680 224540 239844
rect 224650 239816 224678 239912
rect 224724 239844 224730 239896
rect 224782 239844 224788 239896
rect 224604 239788 224678 239816
rect 224604 239760 224632 239788
rect 224742 239760 224770 239844
rect 224834 239828 224862 239912
rect 224926 239884 224954 239912
rect 224926 239856 225000 239884
rect 224834 239788 224868 239828
rect 224862 239776 224868 239788
rect 224920 239776 224926 239828
rect 224586 239708 224592 239760
rect 224644 239708 224650 239760
rect 224678 239708 224684 239760
rect 224736 239720 224770 239760
rect 224736 239708 224742 239720
rect 224972 239692 225000 239856
rect 224770 239680 224776 239692
rect 224512 239652 224776 239680
rect 224770 239640 224776 239652
rect 224828 239640 224834 239692
rect 224954 239640 224960 239692
rect 225012 239640 225018 239692
rect 225110 239680 225138 240400
rect 225386 240156 225414 240468
rect 229434 240156 229462 240468
rect 225294 240128 225414 240156
rect 229250 240134 229462 240156
rect 229158 240128 229462 240134
rect 229802 240156 229830 240808
rect 229940 240700 229968 240876
rect 230124 240768 230152 241012
rect 230584 240836 230612 241148
rect 230584 240808 230704 240836
rect 230124 240740 230612 240768
rect 229940 240672 230244 240700
rect 229802 240128 230014 240156
rect 225294 239952 225322 240128
rect 229158 240106 229278 240128
rect 227042 240060 228450 240088
rect 227042 239964 227070 240060
rect 228422 240020 228450 240060
rect 227456 239992 228082 240020
rect 228422 239992 228634 240020
rect 225552 239952 225558 239964
rect 225294 239924 225558 239952
rect 225552 239912 225558 239924
rect 225610 239912 225616 239964
rect 225736 239952 225742 239964
rect 225708 239912 225742 239952
rect 225794 239912 225800 239964
rect 225828 239912 225834 239964
rect 225886 239952 225892 239964
rect 225886 239912 225920 239952
rect 226104 239912 226110 239964
rect 226162 239912 226168 239964
rect 226380 239912 226386 239964
rect 226438 239912 226444 239964
rect 226472 239912 226478 239964
rect 226530 239912 226536 239964
rect 226840 239912 226846 239964
rect 226898 239952 226904 239964
rect 226898 239912 226932 239952
rect 227024 239912 227030 239964
rect 227082 239912 227088 239964
rect 227300 239912 227306 239964
rect 227358 239952 227364 239964
rect 227358 239912 227392 239952
rect 225184 239844 225190 239896
rect 225242 239844 225248 239896
rect 225460 239884 225466 239896
rect 225432 239844 225466 239884
rect 225518 239844 225524 239896
rect 225202 239760 225230 239844
rect 225202 239720 225236 239760
rect 225230 239708 225236 239720
rect 225288 239708 225294 239760
rect 225110 239652 225184 239680
rect 224494 239612 224500 239624
rect 224420 239584 224500 239612
rect 224494 239572 224500 239584
rect 224552 239572 224558 239624
rect 215168 239516 223804 239544
rect 224006 239516 224816 239544
rect 215168 239504 215174 239516
rect 158530 239436 158536 239488
rect 158588 239476 158594 239488
rect 220538 239476 220544 239488
rect 158588 239448 220544 239476
rect 158588 239436 158594 239448
rect 220538 239436 220544 239448
rect 220596 239476 220602 239488
rect 221274 239476 221280 239488
rect 220596 239448 221280 239476
rect 220596 239436 220602 239448
rect 221274 239436 221280 239448
rect 221332 239436 221338 239488
rect 221366 239436 221372 239488
rect 221424 239476 221430 239488
rect 223482 239476 223488 239488
rect 221424 239448 223488 239476
rect 221424 239436 221430 239448
rect 223482 239436 223488 239448
rect 223540 239436 223546 239488
rect 223776 239476 223804 239516
rect 224402 239476 224408 239488
rect 223776 239448 224408 239476
rect 224402 239436 224408 239448
rect 224460 239436 224466 239488
rect 3326 239368 3332 239420
rect 3384 239408 3390 239420
rect 198918 239408 198924 239420
rect 3384 239380 198924 239408
rect 3384 239368 3390 239380
rect 198918 239368 198924 239380
rect 198976 239368 198982 239420
rect 223298 239408 223304 239420
rect 213886 239380 223304 239408
rect 212166 239300 212172 239352
rect 212224 239340 212230 239352
rect 213886 239340 213914 239380
rect 223298 239368 223304 239380
rect 223356 239408 223362 239420
rect 224678 239408 224684 239420
rect 223356 239380 224684 239408
rect 223356 239368 223362 239380
rect 224678 239368 224684 239380
rect 224736 239368 224742 239420
rect 224788 239408 224816 239516
rect 225156 239488 225184 239652
rect 225432 239624 225460 239844
rect 225414 239572 225420 239624
rect 225472 239572 225478 239624
rect 225708 239544 225736 239912
rect 225782 239776 225788 239828
rect 225840 239816 225846 239828
rect 225892 239816 225920 239912
rect 225840 239788 225920 239816
rect 225840 239776 225846 239788
rect 225966 239640 225972 239692
rect 226024 239680 226030 239692
rect 226122 239680 226150 239912
rect 226024 239652 226150 239680
rect 226398 239692 226426 239912
rect 226490 239760 226518 239912
rect 226748 239844 226754 239896
rect 226806 239844 226812 239896
rect 226766 239760 226794 239844
rect 226490 239720 226524 239760
rect 226518 239708 226524 239720
rect 226576 239708 226582 239760
rect 226766 239720 226800 239760
rect 226794 239708 226800 239720
rect 226852 239708 226858 239760
rect 226398 239652 226432 239692
rect 226024 239640 226030 239652
rect 226426 239640 226432 239652
rect 226484 239640 226490 239692
rect 226904 239612 226932 239912
rect 227208 239844 227214 239896
rect 227266 239844 227272 239896
rect 227226 239760 227254 239844
rect 227162 239708 227168 239760
rect 227220 239720 227254 239760
rect 227220 239708 227226 239720
rect 227070 239640 227076 239692
rect 227128 239680 227134 239692
rect 227364 239680 227392 239912
rect 227128 239652 227392 239680
rect 227128 239640 227134 239652
rect 227456 239624 227484 239992
rect 228054 239964 228082 239992
rect 227668 239912 227674 239964
rect 227726 239912 227732 239964
rect 227944 239952 227950 239964
rect 227824 239924 227950 239952
rect 227686 239760 227714 239912
rect 227824 239760 227852 239924
rect 227944 239912 227950 239924
rect 228002 239912 228008 239964
rect 228036 239912 228042 239964
rect 228094 239912 228100 239964
rect 228496 239952 228502 239964
rect 228146 239924 228502 239952
rect 228146 239884 228174 239924
rect 228496 239912 228502 239924
rect 228554 239912 228560 239964
rect 227916 239856 228174 239884
rect 227622 239708 227628 239760
rect 227680 239720 227714 239760
rect 227680 239708 227686 239720
rect 227806 239708 227812 239760
rect 227864 239708 227870 239760
rect 227346 239612 227352 239624
rect 226904 239584 227352 239612
rect 227346 239572 227352 239584
rect 227404 239572 227410 239624
rect 227438 239572 227444 239624
rect 227496 239572 227502 239624
rect 227916 239612 227944 239856
rect 228220 239844 228226 239896
rect 228278 239844 228284 239896
rect 228312 239844 228318 239896
rect 228370 239844 228376 239896
rect 227990 239776 227996 239828
rect 228048 239816 228054 239828
rect 228238 239816 228266 239844
rect 228048 239788 228266 239816
rect 228048 239776 228054 239788
rect 228330 239680 228358 239844
rect 228330 239652 228496 239680
rect 228468 239624 228496 239652
rect 228606 239624 228634 239992
rect 229158 239964 229186 240106
rect 228864 239952 228870 239964
rect 228836 239912 228870 239952
rect 228922 239912 228928 239964
rect 229140 239912 229146 239964
rect 229198 239912 229204 239964
rect 229232 239912 229238 239964
rect 229290 239912 229296 239964
rect 229324 239912 229330 239964
rect 229382 239912 229388 239964
rect 229416 239912 229422 239964
rect 229474 239912 229480 239964
rect 229876 239912 229882 239964
rect 229934 239912 229940 239964
rect 228680 239844 228686 239896
rect 228738 239884 228744 239896
rect 228738 239844 228772 239884
rect 228744 239624 228772 239844
rect 228836 239624 228864 239912
rect 229250 239624 229278 239912
rect 229342 239828 229370 239912
rect 229434 239884 229462 239912
rect 229784 239884 229790 239896
rect 229434 239856 229508 239884
rect 229342 239788 229376 239828
rect 229370 239776 229376 239788
rect 229428 239776 229434 239828
rect 228174 239612 228180 239624
rect 227916 239584 228180 239612
rect 228174 239572 228180 239584
rect 228232 239572 228238 239624
rect 228450 239572 228456 239624
rect 228508 239572 228514 239624
rect 228542 239572 228548 239624
rect 228600 239584 228634 239624
rect 228600 239572 228606 239584
rect 228726 239572 228732 239624
rect 228784 239572 228790 239624
rect 228818 239572 228824 239624
rect 228876 239572 228882 239624
rect 229250 239584 229284 239624
rect 229278 239572 229284 239584
rect 229336 239572 229342 239624
rect 225248 239516 225736 239544
rect 225248 239488 225276 239516
rect 229094 239504 229100 239556
rect 229152 239544 229158 239556
rect 229480 239544 229508 239856
rect 229664 239856 229790 239884
rect 229664 239624 229692 239856
rect 229784 239844 229790 239856
rect 229842 239844 229848 239896
rect 229894 239760 229922 239912
rect 229830 239708 229836 239760
rect 229888 239720 229922 239760
rect 229986 239760 230014 240128
rect 230060 239912 230066 239964
rect 230118 239952 230124 239964
rect 230118 239912 230152 239952
rect 229986 239720 230020 239760
rect 229888 239708 229894 239720
rect 230014 239708 230020 239720
rect 230072 239708 230078 239760
rect 229646 239572 229652 239624
rect 229704 239572 229710 239624
rect 229152 239516 229508 239544
rect 229152 239504 229158 239516
rect 225138 239436 225144 239488
rect 225196 239436 225202 239488
rect 225230 239436 225236 239488
rect 225288 239436 225294 239488
rect 225506 239436 225512 239488
rect 225564 239476 225570 239488
rect 226058 239476 226064 239488
rect 225564 239448 226064 239476
rect 225564 239436 225570 239448
rect 226058 239436 226064 239448
rect 226116 239436 226122 239488
rect 226610 239436 226616 239488
rect 226668 239476 226674 239488
rect 229738 239476 229744 239488
rect 226668 239448 229744 239476
rect 226668 239436 226674 239448
rect 229738 239436 229744 239448
rect 229796 239436 229802 239488
rect 230124 239420 230152 239912
rect 230216 239476 230244 240672
rect 230584 240020 230612 240740
rect 230676 240088 230704 240808
rect 233758 240224 233786 241420
rect 233758 240196 233878 240224
rect 230676 240060 233602 240088
rect 230584 239992 232314 240020
rect 232286 239964 232314 239992
rect 233574 239964 233602 240060
rect 233850 239964 233878 240196
rect 234218 239964 234246 241488
rect 270218 241476 270224 241528
rect 270276 241516 270282 241528
rect 273346 241516 273352 241528
rect 270276 241488 273352 241516
rect 270276 241476 270282 241488
rect 273346 241476 273352 241488
rect 273404 241476 273410 241528
rect 321002 241476 321008 241528
rect 321060 241516 321066 241528
rect 321462 241516 321468 241528
rect 321060 241488 321468 241516
rect 321060 241476 321066 241488
rect 321462 241476 321468 241488
rect 321520 241516 321526 241528
rect 488534 241516 488540 241528
rect 321520 241488 488540 241516
rect 321520 241476 321526 241488
rect 488534 241476 488540 241488
rect 488592 241476 488598 241528
rect 271414 241380 271420 241392
rect 258046 241352 271420 241380
rect 258046 241312 258074 241352
rect 271414 241340 271420 241352
rect 271472 241340 271478 241392
rect 271322 241312 271328 241324
rect 247006 241284 258074 241312
rect 266326 241284 271328 241312
rect 247006 241108 247034 241284
rect 266326 241244 266354 241284
rect 271322 241272 271328 241284
rect 271380 241272 271386 241324
rect 273254 241272 273260 241324
rect 273312 241312 273318 241324
rect 273898 241312 273904 241324
rect 273312 241284 273904 241312
rect 273312 241272 273318 241284
rect 273898 241272 273904 241284
rect 273956 241272 273962 241324
rect 283558 241244 283564 241256
rect 234862 241080 247034 241108
rect 251146 241216 266354 241244
rect 271156 241216 283564 241244
rect 234862 239964 234890 241080
rect 251146 240836 251174 241216
rect 271046 241176 271052 241188
rect 239140 240808 251174 240836
rect 252526 241148 271052 241176
rect 239140 240496 239168 240808
rect 238910 240468 239168 240496
rect 237622 240128 238478 240156
rect 234954 239992 236086 240020
rect 230520 239952 230526 239964
rect 230446 239924 230526 239952
rect 230446 239544 230474 239924
rect 230520 239912 230526 239924
rect 230578 239912 230584 239964
rect 230980 239952 230986 239964
rect 230722 239924 230986 239952
rect 230722 239680 230750 239924
rect 230980 239912 230986 239924
rect 231038 239912 231044 239964
rect 231256 239912 231262 239964
rect 231314 239912 231320 239964
rect 231716 239952 231722 239964
rect 231642 239924 231722 239952
rect 230796 239844 230802 239896
rect 230854 239844 230860 239896
rect 231274 239884 231302 239912
rect 231044 239856 231302 239884
rect 230676 239652 230750 239680
rect 230676 239624 230704 239652
rect 230814 239624 230842 239844
rect 230658 239572 230664 239624
rect 230716 239572 230722 239624
rect 230750 239572 230756 239624
rect 230808 239584 230842 239624
rect 231044 239612 231072 239856
rect 231440 239844 231446 239896
rect 231498 239844 231504 239896
rect 231118 239708 231124 239760
rect 231176 239748 231182 239760
rect 231458 239748 231486 239844
rect 231176 239720 231486 239748
rect 231176 239708 231182 239720
rect 231394 239640 231400 239692
rect 231452 239680 231458 239692
rect 231642 239680 231670 239924
rect 231716 239912 231722 239924
rect 231774 239912 231780 239964
rect 232268 239912 232274 239964
rect 232326 239912 232332 239964
rect 232452 239952 232458 239964
rect 232424 239912 232458 239952
rect 232510 239912 232516 239964
rect 232636 239952 232642 239964
rect 232608 239912 232642 239952
rect 232694 239912 232700 239964
rect 232912 239912 232918 239964
rect 232970 239952 232976 239964
rect 232970 239912 233004 239952
rect 233372 239912 233378 239964
rect 233430 239912 233436 239964
rect 233464 239912 233470 239964
rect 233522 239912 233528 239964
rect 233556 239912 233562 239964
rect 233614 239912 233620 239964
rect 233648 239912 233654 239964
rect 233706 239912 233712 239964
rect 233740 239912 233746 239964
rect 233798 239912 233804 239964
rect 233832 239912 233838 239964
rect 233890 239912 233896 239964
rect 233924 239912 233930 239964
rect 233982 239912 233988 239964
rect 234200 239912 234206 239964
rect 234258 239912 234264 239964
rect 234292 239912 234298 239964
rect 234350 239912 234356 239964
rect 234752 239912 234758 239964
rect 234810 239912 234816 239964
rect 234844 239912 234850 239964
rect 234902 239912 234908 239964
rect 231900 239884 231906 239896
rect 231872 239844 231906 239884
rect 231958 239844 231964 239896
rect 231872 239760 231900 239844
rect 231854 239708 231860 239760
rect 231912 239708 231918 239760
rect 232424 239692 232452 239912
rect 232608 239692 232636 239912
rect 231452 239652 231670 239680
rect 231452 239640 231458 239652
rect 232406 239640 232412 239692
rect 232464 239640 232470 239692
rect 232590 239640 232596 239692
rect 232648 239640 232654 239692
rect 232976 239680 233004 239912
rect 233280 239844 233286 239896
rect 233338 239844 233344 239896
rect 233298 239760 233326 239844
rect 233390 239828 233418 239912
rect 233482 239884 233510 239912
rect 233482 239856 233556 239884
rect 233528 239828 233556 239856
rect 233390 239788 233424 239828
rect 233418 239776 233424 239788
rect 233476 239776 233482 239828
rect 233510 239776 233516 239828
rect 233568 239776 233574 239828
rect 233666 239760 233694 239912
rect 233758 239828 233786 239912
rect 233942 239884 233970 239912
rect 234310 239884 234338 239912
rect 233896 239856 233970 239884
rect 234264 239856 234338 239884
rect 233896 239828 233924 239856
rect 234264 239828 234292 239856
rect 234568 239844 234574 239896
rect 234626 239844 234632 239896
rect 233758 239788 233792 239828
rect 233786 239776 233792 239788
rect 233844 239776 233850 239828
rect 233878 239776 233884 239828
rect 233936 239776 233942 239828
rect 234246 239776 234252 239828
rect 234304 239776 234310 239828
rect 234586 239760 234614 239844
rect 233298 239720 233332 239760
rect 233326 239708 233332 239720
rect 233384 239708 233390 239760
rect 233666 239720 233700 239760
rect 233694 239708 233700 239720
rect 233752 239708 233758 239760
rect 234586 239720 234620 239760
rect 234614 239708 234620 239720
rect 234672 239708 234678 239760
rect 233234 239680 233240 239692
rect 232976 239652 233240 239680
rect 233234 239640 233240 239652
rect 233292 239640 233298 239692
rect 234770 239680 234798 239912
rect 234080 239652 234798 239680
rect 231118 239612 231124 239624
rect 231044 239584 231124 239612
rect 230808 239572 230814 239584
rect 231118 239572 231124 239584
rect 231176 239572 231182 239624
rect 231946 239544 231952 239556
rect 230446 239516 231952 239544
rect 231946 239504 231952 239516
rect 232004 239504 232010 239556
rect 233234 239504 233240 239556
rect 233292 239544 233298 239556
rect 233418 239544 233424 239556
rect 233292 239516 233424 239544
rect 233292 239504 233298 239516
rect 233418 239504 233424 239516
rect 233476 239504 233482 239556
rect 232774 239476 232780 239488
rect 230216 239448 232780 239476
rect 232774 239436 232780 239448
rect 232832 239436 232838 239488
rect 232866 239436 232872 239488
rect 232924 239476 232930 239488
rect 233050 239476 233056 239488
rect 232924 239448 233056 239476
rect 232924 239436 232930 239448
rect 233050 239436 233056 239448
rect 233108 239436 233114 239488
rect 233142 239436 233148 239488
rect 233200 239476 233206 239488
rect 234080 239476 234108 239652
rect 234246 239572 234252 239624
rect 234304 239612 234310 239624
rect 234430 239612 234436 239624
rect 234304 239584 234436 239612
rect 234304 239572 234310 239584
rect 234430 239572 234436 239584
rect 234488 239572 234494 239624
rect 234614 239572 234620 239624
rect 234672 239612 234678 239624
rect 234954 239612 234982 239992
rect 236058 239964 236086 239992
rect 236196 239992 236454 240020
rect 235028 239912 235034 239964
rect 235086 239912 235092 239964
rect 235396 239912 235402 239964
rect 235454 239912 235460 239964
rect 235580 239912 235586 239964
rect 235638 239912 235644 239964
rect 235672 239912 235678 239964
rect 235730 239912 235736 239964
rect 236040 239912 236046 239964
rect 236098 239912 236104 239964
rect 234672 239584 234982 239612
rect 234672 239572 234678 239584
rect 233200 239448 234108 239476
rect 233200 239436 233206 239448
rect 234338 239436 234344 239488
rect 234396 239476 234402 239488
rect 234522 239476 234528 239488
rect 234396 239448 234528 239476
rect 234396 239436 234402 239448
rect 234522 239436 234528 239448
rect 234580 239436 234586 239488
rect 235046 239476 235074 239912
rect 235414 239760 235442 239912
rect 235598 239760 235626 239912
rect 235690 239816 235718 239912
rect 235856 239844 235862 239896
rect 235914 239884 235920 239896
rect 235914 239844 235948 239884
rect 235690 239788 235764 239816
rect 235414 239720 235448 239760
rect 235442 239708 235448 239720
rect 235500 239708 235506 239760
rect 235598 239720 235632 239760
rect 235626 239708 235632 239720
rect 235684 239708 235690 239760
rect 235258 239572 235264 239624
rect 235316 239612 235322 239624
rect 235736 239612 235764 239788
rect 235920 239760 235948 239844
rect 236196 239760 236224 239992
rect 236426 239964 236454 239992
rect 237162 239992 237558 240020
rect 236316 239952 236322 239964
rect 236288 239912 236322 239952
rect 236374 239912 236380 239964
rect 236408 239912 236414 239964
rect 236466 239912 236472 239964
rect 236592 239912 236598 239964
rect 236650 239912 236656 239964
rect 236960 239912 236966 239964
rect 237018 239912 237024 239964
rect 237052 239912 237058 239964
rect 237110 239912 237116 239964
rect 236288 239760 236316 239912
rect 235902 239708 235908 239760
rect 235960 239708 235966 239760
rect 236178 239708 236184 239760
rect 236236 239708 236242 239760
rect 236270 239708 236276 239760
rect 236328 239708 236334 239760
rect 236454 239680 236460 239692
rect 235316 239584 235764 239612
rect 236104 239652 236460 239680
rect 235316 239572 235322 239584
rect 235810 239476 235816 239488
rect 235046 239448 235816 239476
rect 235810 239436 235816 239448
rect 235868 239436 235874 239488
rect 224788 239380 225460 239408
rect 212224 239312 213914 239340
rect 212224 239300 212230 239312
rect 217778 239300 217784 239352
rect 217836 239340 217842 239352
rect 224494 239340 224500 239352
rect 217836 239312 224500 239340
rect 217836 239300 217842 239312
rect 224494 239300 224500 239312
rect 224552 239300 224558 239352
rect 225138 239300 225144 239352
rect 225196 239340 225202 239352
rect 225432 239340 225460 239380
rect 225690 239368 225696 239420
rect 225748 239408 225754 239420
rect 227990 239408 227996 239420
rect 225748 239380 227996 239408
rect 225748 239368 225754 239380
rect 227990 239368 227996 239380
rect 228048 239368 228054 239420
rect 230106 239368 230112 239420
rect 230164 239368 230170 239420
rect 230658 239368 230664 239420
rect 230716 239408 230722 239420
rect 236104 239408 236132 239652
rect 236454 239640 236460 239652
rect 236512 239680 236518 239692
rect 236610 239680 236638 239912
rect 236868 239884 236874 239896
rect 236512 239652 236638 239680
rect 236748 239856 236874 239884
rect 236748 239680 236776 239856
rect 236868 239844 236874 239856
rect 236926 239844 236932 239896
rect 236978 239828 237006 239912
rect 236960 239776 236966 239828
rect 237018 239776 237024 239828
rect 236822 239708 236828 239760
rect 236880 239748 236886 239760
rect 237070 239748 237098 239912
rect 236880 239720 237098 239748
rect 236880 239708 236886 239720
rect 236914 239680 236920 239692
rect 236748 239652 236920 239680
rect 236512 239640 236518 239652
rect 236914 239640 236920 239652
rect 236972 239640 236978 239692
rect 236178 239572 236184 239624
rect 236236 239612 236242 239624
rect 237162 239612 237190 239992
rect 237530 239964 237558 239992
rect 237328 239952 237334 239964
rect 236236 239584 237190 239612
rect 237300 239912 237334 239952
rect 237386 239912 237392 239964
rect 237512 239912 237518 239964
rect 237570 239912 237576 239964
rect 236236 239572 236242 239584
rect 237098 239504 237104 239556
rect 237156 239544 237162 239556
rect 237300 239544 237328 239912
rect 237622 239884 237650 240128
rect 237806 240060 238386 240088
rect 237696 239912 237702 239964
rect 237754 239912 237760 239964
rect 237484 239856 237650 239884
rect 237484 239624 237512 239856
rect 237714 239816 237742 239912
rect 237576 239788 237742 239816
rect 237576 239760 237604 239788
rect 237558 239708 237564 239760
rect 237616 239708 237622 239760
rect 237466 239572 237472 239624
rect 237524 239572 237530 239624
rect 237156 239516 237328 239544
rect 237156 239504 237162 239516
rect 237806 239476 237834 240060
rect 238358 239964 238386 240060
rect 238450 239964 238478 240128
rect 237880 239912 237886 239964
rect 237938 239912 237944 239964
rect 238248 239952 238254 239964
rect 237990 239924 238254 239952
rect 237898 239556 237926 239912
rect 237990 239612 238018 239924
rect 238248 239912 238254 239924
rect 238306 239912 238312 239964
rect 238340 239912 238346 239964
rect 238398 239912 238404 239964
rect 238432 239912 238438 239964
rect 238490 239912 238496 239964
rect 238910 239896 238938 240468
rect 252526 240292 252554 241148
rect 271046 241136 271052 241148
rect 271104 241136 271110 241188
rect 268102 240864 268108 240916
rect 268160 240904 268166 240916
rect 271156 240904 271184 241216
rect 283558 241204 283564 241216
rect 283616 241244 283622 241256
rect 308582 241244 308588 241256
rect 283616 241216 308588 241244
rect 283616 241204 283622 241216
rect 308582 241204 308588 241216
rect 308640 241204 308646 241256
rect 282270 241176 282276 241188
rect 268160 240876 271184 240904
rect 271248 241148 282276 241176
rect 268160 240864 268166 240876
rect 271248 240836 271276 241148
rect 282270 241136 282276 241148
rect 282328 241176 282334 241188
rect 307294 241176 307300 241188
rect 282328 241148 307300 241176
rect 282328 241136 282334 241148
rect 307294 241136 307300 241148
rect 307352 241136 307358 241188
rect 271506 241068 271512 241120
rect 271564 241108 271570 241120
rect 303154 241108 303160 241120
rect 271564 241080 303160 241108
rect 271564 241068 271570 241080
rect 303154 241068 303160 241080
rect 303212 241068 303218 241120
rect 272058 241000 272064 241052
rect 272116 241040 272122 241052
rect 320082 241040 320088 241052
rect 272116 241012 320088 241040
rect 272116 241000 272122 241012
rect 320082 241000 320088 241012
rect 320140 241000 320146 241052
rect 271690 240932 271696 240984
rect 271748 240972 271754 240984
rect 321002 240972 321008 240984
rect 271748 240944 321008 240972
rect 271748 240932 271754 240944
rect 321002 240932 321008 240944
rect 321060 240932 321066 240984
rect 271414 240864 271420 240916
rect 271472 240904 271478 240916
rect 294966 240904 294972 240916
rect 271472 240876 294972 240904
rect 271472 240864 271478 240876
rect 294966 240864 294972 240876
rect 295024 240864 295030 240916
rect 240106 240264 252554 240292
rect 253952 240808 271276 240836
rect 240106 240224 240134 240264
rect 253952 240224 253980 240808
rect 271322 240796 271328 240848
rect 271380 240836 271386 240848
rect 299106 240836 299112 240848
rect 271380 240808 299112 240836
rect 271380 240796 271386 240808
rect 299106 240796 299112 240808
rect 299164 240796 299170 240848
rect 239646 240196 240134 240224
rect 247374 240196 253980 240224
rect 260484 240740 264284 240768
rect 239076 239912 239082 239964
rect 239134 239912 239140 239964
rect 239536 239952 239542 239964
rect 239324 239924 239542 239952
rect 238064 239844 238070 239896
rect 238122 239884 238128 239896
rect 238524 239884 238530 239896
rect 238122 239856 238248 239884
rect 238122 239844 238128 239856
rect 238220 239816 238248 239856
rect 238496 239844 238530 239884
rect 238582 239844 238588 239896
rect 238616 239844 238622 239896
rect 238674 239844 238680 239896
rect 238800 239884 238806 239896
rect 238772 239844 238806 239884
rect 238858 239844 238864 239896
rect 238892 239844 238898 239896
rect 238950 239844 238956 239896
rect 238294 239816 238300 239828
rect 238220 239788 238300 239816
rect 238294 239776 238300 239788
rect 238352 239776 238358 239828
rect 238496 239760 238524 239844
rect 238634 239760 238662 239844
rect 238772 239760 238800 239844
rect 238478 239708 238484 239760
rect 238536 239708 238542 239760
rect 238570 239708 238576 239760
rect 238628 239720 238662 239760
rect 238628 239708 238634 239720
rect 238754 239708 238760 239760
rect 238812 239708 238818 239760
rect 238110 239640 238116 239692
rect 238168 239680 238174 239692
rect 238910 239680 238938 239844
rect 238168 239652 238938 239680
rect 238168 239640 238174 239652
rect 238202 239612 238208 239624
rect 237990 239584 238208 239612
rect 238202 239572 238208 239584
rect 238260 239572 238266 239624
rect 239094 239612 239122 239912
rect 238772 239584 239122 239612
rect 237898 239516 237932 239556
rect 237926 239504 237932 239516
rect 237984 239504 237990 239556
rect 238772 239488 238800 239584
rect 238018 239476 238024 239488
rect 237806 239448 238024 239476
rect 238018 239436 238024 239448
rect 238076 239436 238082 239488
rect 238754 239436 238760 239488
rect 238812 239436 238818 239488
rect 230716 239380 236132 239408
rect 230716 239368 230722 239380
rect 236730 239368 236736 239420
rect 236788 239408 236794 239420
rect 237006 239408 237012 239420
rect 236788 239380 237012 239408
rect 236788 239368 236794 239380
rect 237006 239368 237012 239380
rect 237064 239368 237070 239420
rect 238846 239368 238852 239420
rect 238904 239408 238910 239420
rect 239324 239408 239352 239924
rect 239536 239912 239542 239924
rect 239594 239912 239600 239964
rect 239646 239760 239674 240196
rect 243418 239992 244044 240020
rect 243418 239964 243446 239992
rect 239904 239912 239910 239964
rect 239962 239912 239968 239964
rect 240088 239952 240094 239964
rect 240060 239912 240094 239952
rect 240146 239912 240152 239964
rect 240364 239912 240370 239964
rect 240422 239912 240428 239964
rect 240824 239912 240830 239964
rect 240882 239912 240888 239964
rect 240916 239912 240922 239964
rect 240974 239912 240980 239964
rect 241008 239912 241014 239964
rect 241066 239952 241072 239964
rect 241192 239952 241198 239964
rect 241066 239912 241100 239952
rect 239720 239844 239726 239896
rect 239778 239844 239784 239896
rect 239582 239708 239588 239760
rect 239640 239720 239674 239760
rect 239640 239708 239646 239720
rect 239490 239436 239496 239488
rect 239548 239476 239554 239488
rect 239738 239476 239766 239844
rect 239922 239624 239950 239912
rect 239858 239572 239864 239624
rect 239916 239584 239950 239624
rect 240060 239612 240088 239912
rect 240382 239816 240410 239912
rect 240548 239884 240554 239896
rect 240520 239844 240554 239884
rect 240606 239844 240612 239896
rect 240382 239788 240456 239816
rect 240134 239612 240140 239624
rect 240060 239584 240140 239612
rect 239916 239572 239922 239584
rect 240134 239572 240140 239584
rect 240192 239572 240198 239624
rect 240428 239612 240456 239788
rect 240520 239692 240548 239844
rect 240502 239640 240508 239692
rect 240560 239640 240566 239692
rect 240686 239612 240692 239624
rect 240428 239584 240692 239612
rect 240686 239572 240692 239584
rect 240744 239572 240750 239624
rect 240842 239556 240870 239912
rect 240934 239748 240962 239912
rect 240934 239720 241008 239748
rect 240842 239516 240876 239556
rect 240870 239504 240876 239516
rect 240928 239504 240934 239556
rect 239548 239448 239766 239476
rect 239548 239436 239554 239448
rect 240778 239436 240784 239488
rect 240836 239476 240842 239488
rect 240980 239476 241008 239720
rect 241072 239692 241100 239912
rect 241164 239912 241198 239952
rect 241250 239912 241256 239964
rect 241468 239912 241474 239964
rect 241526 239912 241532 239964
rect 241928 239912 241934 239964
rect 241986 239912 241992 239964
rect 242020 239912 242026 239964
rect 242078 239952 242084 239964
rect 242078 239912 242112 239952
rect 242388 239912 242394 239964
rect 242446 239912 242452 239964
rect 242756 239952 242762 239964
rect 242728 239912 242762 239952
rect 242814 239912 242820 239964
rect 242848 239912 242854 239964
rect 242906 239912 242912 239964
rect 242940 239912 242946 239964
rect 242998 239912 243004 239964
rect 243124 239912 243130 239964
rect 243182 239912 243188 239964
rect 243308 239912 243314 239964
rect 243366 239912 243372 239964
rect 243400 239912 243406 239964
rect 243458 239912 243464 239964
rect 243676 239912 243682 239964
rect 243734 239912 243740 239964
rect 243860 239912 243866 239964
rect 243918 239912 243924 239964
rect 241054 239640 241060 239692
rect 241112 239640 241118 239692
rect 240836 239448 241008 239476
rect 241164 239476 241192 239912
rect 241284 239844 241290 239896
rect 241342 239844 241348 239896
rect 241302 239624 241330 239844
rect 241486 239692 241514 239912
rect 241836 239844 241842 239896
rect 241894 239844 241900 239896
rect 241854 239816 241882 239844
rect 241808 239788 241882 239816
rect 241486 239652 241520 239692
rect 241514 239640 241520 239652
rect 241572 239640 241578 239692
rect 241808 239680 241836 239788
rect 241946 239760 241974 239912
rect 242084 239760 242112 239912
rect 241882 239708 241888 239760
rect 241940 239720 241974 239760
rect 241940 239708 241946 239720
rect 242066 239708 242072 239760
rect 242124 239708 242130 239760
rect 241974 239680 241980 239692
rect 241808 239652 241980 239680
rect 241974 239640 241980 239652
rect 242032 239640 242038 239692
rect 241238 239572 241244 239624
rect 241296 239584 241330 239624
rect 241296 239572 241302 239584
rect 241330 239476 241336 239488
rect 241164 239448 241336 239476
rect 240836 239436 240842 239448
rect 238904 239380 239352 239408
rect 238904 239368 238910 239380
rect 239398 239368 239404 239420
rect 239456 239408 239462 239420
rect 241164 239408 241192 239448
rect 241330 239436 241336 239448
rect 241388 239436 241394 239488
rect 241790 239436 241796 239488
rect 241848 239476 241854 239488
rect 242406 239476 242434 239912
rect 242728 239692 242756 239912
rect 242866 239692 242894 239912
rect 242710 239640 242716 239692
rect 242768 239640 242774 239692
rect 242802 239640 242808 239692
rect 242860 239652 242894 239692
rect 242958 239692 242986 239912
rect 243032 239844 243038 239896
rect 243090 239844 243096 239896
rect 243050 239748 243078 239844
rect 243142 239816 243170 239912
rect 243326 239884 243354 239912
rect 243326 239856 243492 239884
rect 243142 239788 243308 239816
rect 243050 239720 243124 239748
rect 243096 239692 243124 239720
rect 243280 239692 243308 239788
rect 242958 239652 242992 239692
rect 242860 239640 242866 239652
rect 242986 239640 242992 239652
rect 243044 239640 243050 239692
rect 243078 239640 243084 239692
rect 243136 239640 243142 239692
rect 243262 239640 243268 239692
rect 243320 239640 243326 239692
rect 243464 239624 243492 239856
rect 243446 239572 243452 239624
rect 243504 239572 243510 239624
rect 243354 239504 243360 239556
rect 243412 239544 243418 239556
rect 243694 239544 243722 239912
rect 243878 239760 243906 239912
rect 243814 239708 243820 239760
rect 243872 239720 243906 239760
rect 243872 239708 243878 239720
rect 244016 239692 244044 239992
rect 247374 239964 247402 240196
rect 260484 240156 260512 240740
rect 264256 240700 264284 240740
rect 271046 240728 271052 240780
rect 271104 240768 271110 240780
rect 292758 240768 292764 240780
rect 271104 240740 292764 240768
rect 271104 240728 271110 240740
rect 292758 240728 292764 240740
rect 292816 240728 292822 240780
rect 264256 240672 276014 240700
rect 247696 240128 260512 240156
rect 262922 240604 263226 240632
rect 244412 239912 244418 239964
rect 244470 239912 244476 239964
rect 244688 239912 244694 239964
rect 244746 239952 244752 239964
rect 244746 239912 244780 239952
rect 244964 239912 244970 239964
rect 245022 239952 245028 239964
rect 245332 239952 245338 239964
rect 245022 239924 245148 239952
rect 245022 239912 245028 239924
rect 244136 239884 244142 239896
rect 244108 239844 244142 239884
rect 244194 239844 244200 239896
rect 244228 239844 244234 239896
rect 244286 239844 244292 239896
rect 244108 239760 244136 239844
rect 244090 239708 244096 239760
rect 244148 239708 244154 239760
rect 244246 239748 244274 239844
rect 244430 239816 244458 239912
rect 244504 239844 244510 239896
rect 244562 239884 244568 239896
rect 244562 239856 244688 239884
rect 244562 239844 244568 239856
rect 244430 239788 244596 239816
rect 244200 239720 244274 239748
rect 244200 239692 244228 239720
rect 244568 239692 244596 239788
rect 243998 239640 244004 239692
rect 244056 239640 244062 239692
rect 244182 239640 244188 239692
rect 244240 239640 244246 239692
rect 244550 239640 244556 239692
rect 244608 239640 244614 239692
rect 244458 239572 244464 239624
rect 244516 239612 244522 239624
rect 244660 239612 244688 239856
rect 244752 239760 244780 239912
rect 244734 239708 244740 239760
rect 244792 239708 244798 239760
rect 245010 239748 245016 239760
rect 244844 239720 245016 239748
rect 244516 239584 244688 239612
rect 244516 239572 244522 239584
rect 243412 239516 243722 239544
rect 243412 239504 243418 239516
rect 243998 239504 244004 239556
rect 244056 239544 244062 239556
rect 244366 239544 244372 239556
rect 244056 239516 244372 239544
rect 244056 239504 244062 239516
rect 244366 239504 244372 239516
rect 244424 239504 244430 239556
rect 241848 239448 242434 239476
rect 241848 239436 241854 239448
rect 239456 239380 241192 239408
rect 239456 239368 239462 239380
rect 244366 239368 244372 239420
rect 244424 239408 244430 239420
rect 244844 239408 244872 239720
rect 245010 239708 245016 239720
rect 245068 239708 245074 239760
rect 244918 239572 244924 239624
rect 244976 239612 244982 239624
rect 245120 239612 245148 239924
rect 245212 239924 245338 239952
rect 245212 239624 245240 239924
rect 245332 239912 245338 239924
rect 245390 239912 245396 239964
rect 245516 239952 245522 239964
rect 245488 239912 245522 239952
rect 245574 239912 245580 239964
rect 245608 239912 245614 239964
rect 245666 239912 245672 239964
rect 245976 239952 245982 239964
rect 245948 239912 245982 239952
rect 246034 239912 246040 239964
rect 246528 239912 246534 239964
rect 246586 239912 246592 239964
rect 246620 239912 246626 239964
rect 246678 239912 246684 239964
rect 246804 239912 246810 239964
rect 246862 239912 246868 239964
rect 246988 239912 246994 239964
rect 247046 239912 247052 239964
rect 247080 239912 247086 239964
rect 247138 239912 247144 239964
rect 247264 239912 247270 239964
rect 247322 239912 247328 239964
rect 247356 239912 247362 239964
rect 247414 239912 247420 239964
rect 245488 239624 245516 239912
rect 245626 239624 245654 239912
rect 245700 239844 245706 239896
rect 245758 239844 245764 239896
rect 244976 239584 245148 239612
rect 244976 239572 244982 239584
rect 245194 239572 245200 239624
rect 245252 239572 245258 239624
rect 245470 239572 245476 239624
rect 245528 239572 245534 239624
rect 245562 239572 245568 239624
rect 245620 239584 245654 239624
rect 245620 239572 245626 239584
rect 245718 239544 245746 239844
rect 245304 239516 245746 239544
rect 244424 239380 244872 239408
rect 244424 239368 244430 239380
rect 245010 239368 245016 239420
rect 245068 239408 245074 239420
rect 245304 239408 245332 239516
rect 245948 239476 245976 239912
rect 246068 239844 246074 239896
rect 246126 239844 246132 239896
rect 246160 239844 246166 239896
rect 246218 239844 246224 239896
rect 246252 239844 246258 239896
rect 246310 239844 246316 239896
rect 246344 239844 246350 239896
rect 246402 239884 246408 239896
rect 246402 239844 246436 239884
rect 246086 239816 246114 239844
rect 246040 239788 246114 239816
rect 246040 239760 246068 239788
rect 246178 239760 246206 239844
rect 246022 239708 246028 239760
rect 246080 239708 246086 239760
rect 246114 239708 246120 239760
rect 246172 239720 246206 239760
rect 246172 239708 246178 239720
rect 246270 239692 246298 239844
rect 246270 239652 246304 239692
rect 246298 239640 246304 239652
rect 246356 239640 246362 239692
rect 246408 239544 246436 239844
rect 246546 239816 246574 239912
rect 246500 239788 246574 239816
rect 246638 239816 246666 239912
rect 246638 239788 246712 239816
rect 246500 239692 246528 239788
rect 246684 239760 246712 239788
rect 246822 239760 246850 239912
rect 246666 239708 246672 239760
rect 246724 239708 246730 239760
rect 246822 239720 246856 239760
rect 246850 239708 246856 239720
rect 246908 239708 246914 239760
rect 247006 239692 247034 239912
rect 247098 239760 247126 239912
rect 247282 239760 247310 239912
rect 247540 239844 247546 239896
rect 247598 239844 247604 239896
rect 247098 239720 247132 239760
rect 247126 239708 247132 239720
rect 247184 239708 247190 239760
rect 247218 239708 247224 239760
rect 247276 239720 247310 239760
rect 247276 239708 247282 239720
rect 246482 239640 246488 239692
rect 246540 239640 246546 239692
rect 247006 239652 247040 239692
rect 247034 239640 247040 239652
rect 247092 239640 247098 239692
rect 247558 239624 247586 239844
rect 247494 239572 247500 239624
rect 247552 239584 247586 239624
rect 247552 239572 247558 239584
rect 246574 239544 246580 239556
rect 246408 239516 246580 239544
rect 246574 239504 246580 239516
rect 246632 239504 246638 239556
rect 247696 239488 247724 240128
rect 247788 240060 252048 240088
rect 247310 239476 247316 239488
rect 245948 239448 247316 239476
rect 247310 239436 247316 239448
rect 247368 239436 247374 239488
rect 247678 239436 247684 239488
rect 247736 239436 247742 239488
rect 245068 239380 245332 239408
rect 245068 239368 245074 239380
rect 246298 239368 246304 239420
rect 246356 239408 246362 239420
rect 247034 239408 247040 239420
rect 246356 239380 247040 239408
rect 246356 239368 246362 239380
rect 247034 239368 247040 239380
rect 247092 239368 247098 239420
rect 247402 239368 247408 239420
rect 247460 239408 247466 239420
rect 247788 239408 247816 240060
rect 248386 239992 248782 240020
rect 248000 239912 248006 239964
rect 248058 239912 248064 239964
rect 247862 239572 247868 239624
rect 247920 239612 247926 239624
rect 248018 239612 248046 239912
rect 248386 239680 248414 239992
rect 248754 239964 248782 239992
rect 248938 239992 250898 240020
rect 248938 239964 248966 239992
rect 248460 239912 248466 239964
rect 248518 239952 248524 239964
rect 248518 239912 248552 239952
rect 248644 239912 248650 239964
rect 248702 239912 248708 239964
rect 248736 239912 248742 239964
rect 248794 239912 248800 239964
rect 248828 239912 248834 239964
rect 248886 239912 248892 239964
rect 248920 239912 248926 239964
rect 248978 239912 248984 239964
rect 249012 239912 249018 239964
rect 249070 239912 249076 239964
rect 249196 239912 249202 239964
rect 249254 239912 249260 239964
rect 249380 239912 249386 239964
rect 249438 239912 249444 239964
rect 249472 239912 249478 239964
rect 249530 239912 249536 239964
rect 249932 239912 249938 239964
rect 249990 239912 249996 239964
rect 250116 239912 250122 239964
rect 250174 239912 250180 239964
rect 250300 239912 250306 239964
rect 250358 239912 250364 239964
rect 250484 239952 250490 239964
rect 250456 239912 250490 239952
rect 250542 239912 250548 239964
rect 250576 239912 250582 239964
rect 250634 239912 250640 239964
rect 250760 239912 250766 239964
rect 250818 239912 250824 239964
rect 248524 239760 248552 239912
rect 248662 239760 248690 239912
rect 248846 239760 248874 239912
rect 248506 239708 248512 239760
rect 248564 239708 248570 239760
rect 248662 239720 248696 239760
rect 248690 239708 248696 239720
rect 248748 239708 248754 239760
rect 248782 239708 248788 239760
rect 248840 239720 248874 239760
rect 248840 239708 248846 239720
rect 248874 239680 248880 239692
rect 248386 239652 248880 239680
rect 248874 239640 248880 239652
rect 248932 239640 248938 239692
rect 249030 239680 249058 239912
rect 249214 239816 249242 239912
rect 249288 239844 249294 239896
rect 249346 239844 249352 239896
rect 249168 239788 249242 239816
rect 249168 239760 249196 239788
rect 249306 239760 249334 239844
rect 249150 239708 249156 239760
rect 249208 239708 249214 239760
rect 249242 239708 249248 239760
rect 249300 239720 249334 239760
rect 249300 239708 249306 239720
rect 249398 239692 249426 239912
rect 249030 239652 249196 239680
rect 247920 239584 248046 239612
rect 247920 239572 247926 239584
rect 248874 239504 248880 239556
rect 248932 239544 248938 239556
rect 249168 239544 249196 239652
rect 249334 239640 249340 239692
rect 249392 239652 249426 239692
rect 249490 239680 249518 239912
rect 249656 239844 249662 239896
rect 249714 239844 249720 239896
rect 249840 239844 249846 239896
rect 249898 239844 249904 239896
rect 249674 239760 249702 239844
rect 249610 239708 249616 239760
rect 249668 239720 249702 239760
rect 249668 239708 249674 239720
rect 249490 239652 249610 239680
rect 249392 239640 249398 239652
rect 249582 239612 249610 239652
rect 249858 239624 249886 239844
rect 249702 239612 249708 239624
rect 249582 239584 249708 239612
rect 249702 239572 249708 239584
rect 249760 239572 249766 239624
rect 249794 239572 249800 239624
rect 249852 239584 249886 239624
rect 249852 239572 249858 239584
rect 249950 239556 249978 239912
rect 250134 239556 250162 239912
rect 250318 239760 250346 239912
rect 250456 239760 250484 239912
rect 250594 239760 250622 239912
rect 250778 239816 250806 239912
rect 250870 239884 250898 239992
rect 250962 239992 251772 240020
rect 250962 239964 250990 239992
rect 250944 239912 250950 239964
rect 251002 239912 251008 239964
rect 251128 239952 251134 239964
rect 251054 239924 251134 239952
rect 250870 239856 250944 239884
rect 250778 239788 250852 239816
rect 250824 239760 250852 239788
rect 250254 239708 250260 239760
rect 250312 239720 250346 239760
rect 250312 239708 250318 239720
rect 250438 239708 250444 239760
rect 250496 239708 250502 239760
rect 250594 239720 250628 239760
rect 250622 239708 250628 239720
rect 250680 239708 250686 239760
rect 250806 239708 250812 239760
rect 250864 239708 250870 239760
rect 250530 239640 250536 239692
rect 250588 239680 250594 239692
rect 250916 239680 250944 239856
rect 250588 239652 250944 239680
rect 250588 239640 250594 239652
rect 251054 239624 251082 239924
rect 251128 239912 251134 239924
rect 251186 239912 251192 239964
rect 251220 239844 251226 239896
rect 251278 239844 251284 239896
rect 251496 239844 251502 239896
rect 251554 239844 251560 239896
rect 251588 239844 251594 239896
rect 251646 239844 251652 239896
rect 251238 239692 251266 239844
rect 251174 239640 251180 239692
rect 251232 239652 251266 239692
rect 251232 239640 251238 239652
rect 251514 239624 251542 239844
rect 251054 239584 251088 239624
rect 251082 239572 251088 239584
rect 251140 239572 251146 239624
rect 251450 239572 251456 239624
rect 251508 239584 251542 239624
rect 251606 239624 251634 239844
rect 251744 239680 251772 239992
rect 251864 239912 251870 239964
rect 251922 239952 251928 239964
rect 251922 239912 251956 239952
rect 251744 239652 251864 239680
rect 251836 239624 251864 239652
rect 251606 239584 251640 239624
rect 251508 239572 251514 239584
rect 251634 239572 251640 239584
rect 251692 239572 251698 239624
rect 251818 239572 251824 239624
rect 251876 239572 251882 239624
rect 248932 239516 249196 239544
rect 248932 239504 248938 239516
rect 249886 239504 249892 239556
rect 249944 239516 249978 239556
rect 249944 239504 249950 239516
rect 250070 239504 250076 239556
rect 250128 239516 250162 239556
rect 250128 239504 250134 239516
rect 251358 239504 251364 239556
rect 251416 239544 251422 239556
rect 251928 239544 251956 239912
rect 252020 239624 252048 240060
rect 256482 240060 257154 240088
rect 253308 239992 253658 240020
rect 252508 239912 252514 239964
rect 252566 239952 252572 239964
rect 252566 239912 252600 239952
rect 252968 239912 252974 239964
rect 253026 239952 253032 239964
rect 253026 239912 253060 239952
rect 252140 239844 252146 239896
rect 252198 239844 252204 239896
rect 252324 239844 252330 239896
rect 252382 239844 252388 239896
rect 252002 239572 252008 239624
rect 252060 239572 252066 239624
rect 252158 239556 252186 239844
rect 252342 239760 252370 239844
rect 252342 239720 252376 239760
rect 252370 239708 252376 239720
rect 252428 239708 252434 239760
rect 251416 239516 251956 239544
rect 251416 239504 251422 239516
rect 252094 239504 252100 239556
rect 252152 239516 252186 239556
rect 252572 239544 252600 239912
rect 252692 239844 252698 239896
rect 252750 239844 252756 239896
rect 252710 239692 252738 239844
rect 253032 239692 253060 239912
rect 253152 239844 253158 239896
rect 253210 239884 253216 239896
rect 253210 239844 253244 239884
rect 253216 239692 253244 239844
rect 253308 239692 253336 239992
rect 253630 239964 253658 239992
rect 254918 239992 255130 240020
rect 253428 239952 253434 239964
rect 253400 239912 253434 239952
rect 253486 239912 253492 239964
rect 253520 239912 253526 239964
rect 253578 239912 253584 239964
rect 253612 239912 253618 239964
rect 253670 239912 253676 239964
rect 253888 239912 253894 239964
rect 253946 239912 253952 239964
rect 253980 239912 253986 239964
rect 254038 239912 254044 239964
rect 254256 239912 254262 239964
rect 254314 239912 254320 239964
rect 254440 239912 254446 239964
rect 254498 239912 254504 239964
rect 254808 239952 254814 239964
rect 254780 239912 254814 239952
rect 254866 239912 254872 239964
rect 252646 239640 252652 239692
rect 252704 239652 252738 239692
rect 252704 239640 252710 239652
rect 253014 239640 253020 239692
rect 253072 239640 253078 239692
rect 253198 239640 253204 239692
rect 253256 239640 253262 239692
rect 253290 239640 253296 239692
rect 253348 239640 253354 239692
rect 253400 239612 253428 239912
rect 253538 239680 253566 239912
rect 253658 239680 253664 239692
rect 253538 239652 253664 239680
rect 253658 239640 253664 239652
rect 253716 239640 253722 239692
rect 253750 239640 253756 239692
rect 253808 239680 253814 239692
rect 253906 239680 253934 239912
rect 253808 239652 253934 239680
rect 253808 239640 253814 239652
rect 253998 239624 254026 239912
rect 254274 239760 254302 239912
rect 254274 239720 254308 239760
rect 254302 239708 254308 239720
rect 254360 239708 254366 239760
rect 254458 239680 254486 239912
rect 254624 239844 254630 239896
rect 254682 239844 254688 239896
rect 253566 239612 253572 239624
rect 253400 239584 253572 239612
rect 253566 239572 253572 239584
rect 253624 239572 253630 239624
rect 253934 239572 253940 239624
rect 253992 239584 254026 239624
rect 254136 239652 254486 239680
rect 253992 239572 253998 239584
rect 252830 239544 252836 239556
rect 252572 239516 252836 239544
rect 252152 239504 252158 239516
rect 252830 239504 252836 239516
rect 252888 239504 252894 239556
rect 254136 239544 254164 239652
rect 254210 239572 254216 239624
rect 254268 239612 254274 239624
rect 254642 239612 254670 239844
rect 254780 239692 254808 239912
rect 254918 239884 254946 239992
rect 255102 239964 255130 239992
rect 255194 239992 256418 240020
rect 254992 239912 254998 239964
rect 255050 239912 255056 239964
rect 255084 239912 255090 239964
rect 255142 239912 255148 239964
rect 254872 239856 254946 239884
rect 254762 239640 254768 239692
rect 254820 239640 254826 239692
rect 254268 239584 254670 239612
rect 254872 239612 254900 239856
rect 255010 239760 255038 239912
rect 255194 239760 255222 239992
rect 256390 239964 256418 239992
rect 255268 239912 255274 239964
rect 255326 239912 255332 239964
rect 255452 239912 255458 239964
rect 255510 239912 255516 239964
rect 256004 239912 256010 239964
rect 256062 239912 256068 239964
rect 256096 239912 256102 239964
rect 256154 239912 256160 239964
rect 256372 239912 256378 239964
rect 256430 239912 256436 239964
rect 254946 239708 254952 239760
rect 255004 239720 255038 239760
rect 255004 239708 255010 239720
rect 255130 239708 255136 239760
rect 255188 239720 255222 239760
rect 255286 239748 255314 239912
rect 255470 239816 255498 239912
rect 255728 239844 255734 239896
rect 255786 239844 255792 239896
rect 255820 239844 255826 239896
rect 255878 239844 255884 239896
rect 255470 239788 255636 239816
rect 255498 239748 255504 239760
rect 255286 239720 255504 239748
rect 255188 239708 255194 239720
rect 255498 239708 255504 239720
rect 255556 239708 255562 239760
rect 255222 239612 255228 239624
rect 254872 239584 255228 239612
rect 254268 239572 254274 239584
rect 255222 239572 255228 239584
rect 255280 239572 255286 239624
rect 255608 239556 255636 239788
rect 255746 239624 255774 239844
rect 255838 239692 255866 239844
rect 255838 239652 255872 239692
rect 255866 239640 255872 239652
rect 255924 239640 255930 239692
rect 256022 239624 256050 239912
rect 255746 239584 255780 239624
rect 255774 239572 255780 239584
rect 255832 239572 255838 239624
rect 255958 239572 255964 239624
rect 256016 239584 256050 239624
rect 256114 239624 256142 239912
rect 256280 239884 256286 239896
rect 256252 239844 256286 239884
rect 256338 239844 256344 239896
rect 256252 239692 256280 239844
rect 256234 239640 256240 239692
rect 256292 239640 256298 239692
rect 256326 239640 256332 239692
rect 256384 239680 256390 239692
rect 256482 239680 256510 240060
rect 256666 239992 257062 240020
rect 256666 239964 256694 239992
rect 256556 239912 256562 239964
rect 256614 239912 256620 239964
rect 256648 239912 256654 239964
rect 256706 239912 256712 239964
rect 256924 239952 256930 239964
rect 256804 239924 256930 239952
rect 256384 239652 256510 239680
rect 256384 239640 256390 239652
rect 256114 239584 256148 239624
rect 256016 239572 256022 239584
rect 256142 239572 256148 239584
rect 256200 239572 256206 239624
rect 256574 239556 256602 239912
rect 254486 239544 254492 239556
rect 254136 239516 254492 239544
rect 254486 239504 254492 239516
rect 254544 239504 254550 239556
rect 255130 239504 255136 239556
rect 255188 239544 255194 239556
rect 255406 239544 255412 239556
rect 255188 239516 255412 239544
rect 255188 239504 255194 239516
rect 255406 239504 255412 239516
rect 255464 239504 255470 239556
rect 255590 239504 255596 239556
rect 255648 239504 255654 239556
rect 256510 239504 256516 239556
rect 256568 239516 256602 239556
rect 256804 239544 256832 239924
rect 256924 239912 256930 239924
rect 256982 239912 256988 239964
rect 257034 239884 257062 239992
rect 257126 239964 257154 240060
rect 257310 239992 259270 240020
rect 257310 239964 257338 239992
rect 257108 239912 257114 239964
rect 257166 239912 257172 239964
rect 257292 239912 257298 239964
rect 257350 239912 257356 239964
rect 257476 239912 257482 239964
rect 257534 239912 257540 239964
rect 257568 239912 257574 239964
rect 257626 239912 257632 239964
rect 257752 239912 257758 239964
rect 257810 239912 257816 239964
rect 257844 239912 257850 239964
rect 257902 239912 257908 239964
rect 258396 239952 258402 239964
rect 258368 239912 258402 239952
rect 258454 239912 258460 239964
rect 258488 239912 258494 239964
rect 258546 239912 258552 239964
rect 258672 239912 258678 239964
rect 258730 239912 258736 239964
rect 258856 239912 258862 239964
rect 258914 239912 258920 239964
rect 259132 239912 259138 239964
rect 259190 239912 259196 239964
rect 256896 239856 257062 239884
rect 256896 239624 256924 239856
rect 257200 239844 257206 239896
rect 257258 239844 257264 239896
rect 257218 239760 257246 239844
rect 257154 239708 257160 239760
rect 257212 239720 257246 239760
rect 257212 239708 257218 239720
rect 257494 239624 257522 239912
rect 257586 239748 257614 239912
rect 257586 239720 257660 239748
rect 257632 239692 257660 239720
rect 257770 239692 257798 239912
rect 257614 239640 257620 239692
rect 257672 239640 257678 239692
rect 257706 239640 257712 239692
rect 257764 239652 257798 239692
rect 257764 239640 257770 239652
rect 256878 239572 256884 239624
rect 256936 239572 256942 239624
rect 257494 239584 257528 239624
rect 257522 239572 257528 239584
rect 257580 239572 257586 239624
rect 257862 239612 257890 239912
rect 258212 239844 258218 239896
rect 258270 239844 258276 239896
rect 258230 239680 258258 239844
rect 258368 239760 258396 239912
rect 258506 239828 258534 239912
rect 258442 239776 258448 239828
rect 258500 239788 258534 239828
rect 258500 239776 258506 239788
rect 258350 239708 258356 239760
rect 258408 239708 258414 239760
rect 258534 239680 258540 239692
rect 258230 239652 258540 239680
rect 258534 239640 258540 239652
rect 258592 239640 258598 239692
rect 258258 239612 258264 239624
rect 257862 239584 258264 239612
rect 258258 239572 258264 239584
rect 258316 239572 258322 239624
rect 257062 239544 257068 239556
rect 256804 239516 257068 239544
rect 256568 239504 256574 239516
rect 257062 239504 257068 239516
rect 257120 239544 257126 239556
rect 257798 239544 257804 239556
rect 257120 239516 257804 239544
rect 257120 239504 257126 239516
rect 257798 239504 257804 239516
rect 257856 239504 257862 239556
rect 257982 239504 257988 239556
rect 258040 239544 258046 239556
rect 258690 239544 258718 239912
rect 258874 239760 258902 239912
rect 259150 239816 259178 239912
rect 258810 239708 258816 239760
rect 258868 239720 258902 239760
rect 259104 239788 259178 239816
rect 258868 239708 258874 239720
rect 259104 239624 259132 239788
rect 259242 239760 259270 239992
rect 260530 239992 260880 240020
rect 260530 239964 260558 239992
rect 259316 239912 259322 239964
rect 259374 239912 259380 239964
rect 259684 239912 259690 239964
rect 259742 239912 259748 239964
rect 260052 239912 260058 239964
rect 260110 239912 260116 239964
rect 260420 239912 260426 239964
rect 260478 239912 260484 239964
rect 260512 239912 260518 239964
rect 260570 239912 260576 239964
rect 260604 239912 260610 239964
rect 260662 239912 260668 239964
rect 260696 239912 260702 239964
rect 260754 239912 260760 239964
rect 259334 239816 259362 239912
rect 259334 239788 259500 239816
rect 259178 239708 259184 239760
rect 259236 239720 259270 239760
rect 259236 239708 259242 239720
rect 259472 239692 259500 239788
rect 259454 239640 259460 239692
rect 259512 239640 259518 239692
rect 259702 239624 259730 239912
rect 259086 239572 259092 239624
rect 259144 239572 259150 239624
rect 259638 239612 259644 239624
rect 259597 239584 259644 239612
rect 259638 239572 259644 239584
rect 259696 239612 259730 239624
rect 259914 239612 259920 239624
rect 259696 239584 259920 239612
rect 259696 239572 259702 239584
rect 259914 239572 259920 239584
rect 259972 239572 259978 239624
rect 260070 239612 260098 239912
rect 260438 239828 260466 239912
rect 260622 239828 260650 239912
rect 260438 239788 260472 239828
rect 260466 239776 260472 239788
rect 260524 239776 260530 239828
rect 260558 239776 260564 239828
rect 260616 239788 260650 239828
rect 260616 239776 260622 239788
rect 260714 239760 260742 239912
rect 260650 239708 260656 239760
rect 260708 239720 260742 239760
rect 260708 239708 260714 239720
rect 260852 239692 260880 239992
rect 262922 239964 262950 240604
rect 263198 240360 263226 240604
rect 275986 240564 276014 240672
rect 278130 240564 278136 240576
rect 275986 240536 278136 240564
rect 278130 240524 278136 240536
rect 278188 240524 278194 240576
rect 267918 240456 267924 240508
rect 267976 240496 267982 240508
rect 267976 240468 270494 240496
rect 267976 240456 267982 240468
rect 270466 240428 270494 240468
rect 270466 240400 274634 240428
rect 271230 240360 271236 240372
rect 263198 240332 271236 240360
rect 271230 240320 271236 240332
rect 271288 240320 271294 240372
rect 267734 240292 267740 240304
rect 263290 240264 267740 240292
rect 263290 239964 263318 240264
rect 267734 240252 267740 240264
rect 267792 240252 267798 240304
rect 268102 240224 268108 240236
rect 265866 240196 268108 240224
rect 265866 240088 265894 240196
rect 268102 240184 268108 240196
rect 268160 240224 268166 240236
rect 273070 240224 273076 240236
rect 268160 240196 273076 240224
rect 268160 240184 268166 240196
rect 273070 240184 273076 240196
rect 273128 240184 273134 240236
rect 269206 240156 269212 240168
rect 266326 240128 269212 240156
rect 266326 240088 266354 240128
rect 269206 240116 269212 240128
rect 269264 240116 269270 240168
rect 274606 240156 274634 240400
rect 276014 240156 276020 240168
rect 274606 240128 276020 240156
rect 276014 240116 276020 240128
rect 276072 240116 276078 240168
rect 267918 240088 267924 240100
rect 264026 240060 265894 240088
rect 265958 240060 266354 240088
rect 266878 240060 267924 240088
rect 264026 239964 264054 240060
rect 265958 240020 265986 240060
rect 266878 240020 266906 240060
rect 267918 240048 267924 240060
rect 267976 240048 267982 240100
rect 270494 240020 270500 240032
rect 264118 239992 265986 240020
rect 266142 239992 266906 240020
rect 266970 239992 270500 240020
rect 260972 239912 260978 239964
rect 261030 239912 261036 239964
rect 261432 239912 261438 239964
rect 261490 239952 261496 239964
rect 261892 239952 261898 239964
rect 261490 239912 261524 239952
rect 260834 239640 260840 239692
rect 260892 239640 260898 239692
rect 260190 239612 260196 239624
rect 260070 239584 260196 239612
rect 260190 239572 260196 239584
rect 260248 239572 260254 239624
rect 258040 239516 258718 239544
rect 258040 239504 258046 239516
rect 260834 239504 260840 239556
rect 260892 239544 260898 239556
rect 260990 239544 261018 239912
rect 261248 239844 261254 239896
rect 261306 239844 261312 239896
rect 261340 239844 261346 239896
rect 261398 239884 261404 239896
rect 261398 239844 261432 239884
rect 261266 239692 261294 239844
rect 261266 239652 261300 239692
rect 261294 239640 261300 239652
rect 261352 239640 261358 239692
rect 261404 239556 261432 239844
rect 261496 239760 261524 239912
rect 261864 239912 261898 239952
rect 261950 239912 261956 239964
rect 261984 239912 261990 239964
rect 262042 239912 262048 239964
rect 262076 239912 262082 239964
rect 262134 239912 262140 239964
rect 262168 239912 262174 239964
rect 262226 239952 262232 239964
rect 262352 239952 262358 239964
rect 262226 239912 262260 239952
rect 261616 239884 261622 239896
rect 261588 239844 261622 239884
rect 261674 239844 261680 239896
rect 261708 239844 261714 239896
rect 261766 239844 261772 239896
rect 261588 239760 261616 239844
rect 261726 239760 261754 239844
rect 261478 239708 261484 239760
rect 261536 239708 261542 239760
rect 261570 239708 261576 239760
rect 261628 239708 261634 239760
rect 261662 239708 261668 239760
rect 261720 239720 261754 239760
rect 261864 239748 261892 239912
rect 262002 239828 262030 239912
rect 262094 239884 262122 239912
rect 262094 239856 262168 239884
rect 262140 239828 262168 239856
rect 261938 239776 261944 239828
rect 261996 239788 262030 239828
rect 261996 239776 262002 239788
rect 262122 239776 262128 239828
rect 262180 239776 262186 239828
rect 262030 239748 262036 239760
rect 261864 239720 262036 239748
rect 261720 239708 261726 239720
rect 262030 239708 262036 239720
rect 262088 239708 262094 239760
rect 262232 239692 262260 239912
rect 262324 239912 262358 239952
rect 262410 239912 262416 239964
rect 262444 239912 262450 239964
rect 262502 239912 262508 239964
rect 262812 239912 262818 239964
rect 262870 239912 262876 239964
rect 262904 239912 262910 239964
rect 262962 239912 262968 239964
rect 262996 239912 263002 239964
rect 263054 239912 263060 239964
rect 263272 239912 263278 239964
rect 263330 239912 263336 239964
rect 263364 239912 263370 239964
rect 263422 239912 263428 239964
rect 263824 239912 263830 239964
rect 263882 239912 263888 239964
rect 264008 239912 264014 239964
rect 264066 239912 264072 239964
rect 262214 239640 262220 239692
rect 262272 239640 262278 239692
rect 262324 239612 262352 239912
rect 262462 239828 262490 239912
rect 262398 239776 262404 239828
rect 262456 239788 262490 239828
rect 262456 239776 262462 239788
rect 262830 239748 262858 239912
rect 263014 239884 263042 239912
rect 262968 239856 263042 239884
rect 262968 239828 262996 239856
rect 263180 239844 263186 239896
rect 263238 239844 263244 239896
rect 262950 239776 262956 239828
rect 263008 239776 263014 239828
rect 263042 239748 263048 239760
rect 262830 239720 263048 239748
rect 263042 239708 263048 239720
rect 263100 239708 263106 239760
rect 263198 239748 263226 239844
rect 263152 239720 263226 239748
rect 262858 239640 262864 239692
rect 262916 239680 262922 239692
rect 263152 239680 263180 239720
rect 263290 239692 263318 239912
rect 262916 239652 263180 239680
rect 262916 239640 262922 239652
rect 263226 239640 263232 239692
rect 263284 239652 263318 239692
rect 263382 239680 263410 239912
rect 263842 239884 263870 239912
rect 264118 239884 264146 239992
rect 266142 239964 266170 239992
rect 266970 239964 266998 239992
rect 270494 239980 270500 239992
rect 270552 239980 270558 240032
rect 264284 239912 264290 239964
rect 264342 239912 264348 239964
rect 264376 239912 264382 239964
rect 264434 239952 264440 239964
rect 264434 239912 264468 239952
rect 264652 239912 264658 239964
rect 264710 239912 264716 239964
rect 265020 239952 265026 239964
rect 264946 239924 265026 239952
rect 263842 239856 264146 239884
rect 263888 239692 263916 239856
rect 264302 239828 264330 239912
rect 264302 239788 264336 239828
rect 264330 239776 264336 239788
rect 264388 239776 264394 239828
rect 264440 239692 264468 239912
rect 264514 239708 264520 239760
rect 264572 239748 264578 239760
rect 264670 239748 264698 239912
rect 264836 239844 264842 239896
rect 264894 239844 264900 239896
rect 264572 239720 264698 239748
rect 264572 239708 264578 239720
rect 264854 239692 264882 239844
rect 263502 239680 263508 239692
rect 263382 239652 263508 239680
rect 263284 239640 263290 239652
rect 263502 239640 263508 239652
rect 263560 239640 263566 239692
rect 263870 239640 263876 239692
rect 263928 239640 263934 239692
rect 264422 239640 264428 239692
rect 264480 239640 264486 239692
rect 264790 239640 264796 239692
rect 264848 239652 264882 239692
rect 264848 239640 264854 239652
rect 264946 239624 264974 239924
rect 265020 239912 265026 239924
rect 265078 239912 265084 239964
rect 265572 239912 265578 239964
rect 265630 239912 265636 239964
rect 265756 239952 265762 239964
rect 265728 239912 265762 239952
rect 265814 239912 265820 239964
rect 266124 239912 266130 239964
rect 266182 239912 266188 239964
rect 266308 239912 266314 239964
rect 266366 239912 266372 239964
rect 266676 239952 266682 239964
rect 266648 239912 266682 239952
rect 266734 239912 266740 239964
rect 266952 239912 266958 239964
rect 267010 239912 267016 239964
rect 267044 239912 267050 239964
rect 267102 239952 267108 239964
rect 268010 239952 268016 239964
rect 267102 239924 268016 239952
rect 267102 239912 267108 239924
rect 268010 239912 268016 239924
rect 268068 239912 268074 239964
rect 268470 239912 268476 239964
rect 268528 239952 268534 239964
rect 269206 239952 269212 239964
rect 268528 239924 269212 239952
rect 268528 239912 268534 239924
rect 269206 239912 269212 239924
rect 269264 239912 269270 239964
rect 265112 239844 265118 239896
rect 265170 239844 265176 239896
rect 265204 239844 265210 239896
rect 265262 239844 265268 239896
rect 265296 239844 265302 239896
rect 265354 239844 265360 239896
rect 265130 239692 265158 239844
rect 265066 239640 265072 239692
rect 265124 239652 265158 239692
rect 265124 239640 265130 239652
rect 263134 239612 263140 239624
rect 262324 239584 263140 239612
rect 263134 239572 263140 239584
rect 263192 239572 263198 239624
rect 264882 239572 264888 239624
rect 264940 239584 264974 239624
rect 264940 239572 264946 239584
rect 261386 239544 261392 239556
rect 260892 239516 261018 239544
rect 261299 239516 261392 239544
rect 260892 239504 260898 239516
rect 261386 239504 261392 239516
rect 261444 239544 261450 239556
rect 262674 239544 262680 239556
rect 261444 239516 262680 239544
rect 261444 239504 261450 239516
rect 262674 239504 262680 239516
rect 262732 239504 262738 239556
rect 265222 239488 265250 239844
rect 265314 239544 265342 239844
rect 265590 239612 265618 239912
rect 265728 239748 265756 239912
rect 265940 239844 265946 239896
rect 265998 239884 266004 239896
rect 265998 239844 266032 239884
rect 266004 239760 266032 239844
rect 266326 239816 266354 239912
rect 266400 239844 266406 239896
rect 266458 239844 266464 239896
rect 266492 239844 266498 239896
rect 266550 239844 266556 239896
rect 266280 239788 266354 239816
rect 266280 239760 266308 239788
rect 266418 239760 266446 239844
rect 265894 239748 265900 239760
rect 265728 239720 265900 239748
rect 265894 239708 265900 239720
rect 265952 239708 265958 239760
rect 265986 239708 265992 239760
rect 266044 239708 266050 239760
rect 266262 239708 266268 239760
rect 266320 239708 266326 239760
rect 266354 239708 266360 239760
rect 266412 239720 266446 239760
rect 266510 239760 266538 239844
rect 266648 239760 266676 239912
rect 267062 239828 267090 239912
rect 267136 239844 267142 239896
rect 267194 239884 267200 239896
rect 267826 239884 267832 239896
rect 267194 239856 267832 239884
rect 267194 239844 267200 239856
rect 267826 239844 267832 239856
rect 267884 239844 267890 239896
rect 266998 239776 267004 239828
rect 267056 239788 267090 239828
rect 267056 239776 267062 239788
rect 266510 239720 266544 239760
rect 266412 239708 266418 239720
rect 266538 239708 266544 239720
rect 266596 239708 266602 239760
rect 266630 239708 266636 239760
rect 266688 239708 266694 239760
rect 266814 239708 266820 239760
rect 266872 239748 266878 239760
rect 267154 239748 267182 239844
rect 266872 239720 267182 239748
rect 266872 239708 266878 239720
rect 270954 239708 270960 239760
rect 271012 239748 271018 239760
rect 271012 239720 278084 239748
rect 271012 239708 271018 239720
rect 266906 239640 266912 239692
rect 266964 239680 266970 239692
rect 269114 239680 269120 239692
rect 266964 239652 269120 239680
rect 266964 239640 266970 239652
rect 269114 239640 269120 239652
rect 269172 239640 269178 239692
rect 266170 239612 266176 239624
rect 265590 239584 266176 239612
rect 266170 239572 266176 239584
rect 266228 239572 266234 239624
rect 267366 239572 267372 239624
rect 267424 239612 267430 239624
rect 269298 239612 269304 239624
rect 267424 239584 269304 239612
rect 267424 239572 267430 239584
rect 269298 239572 269304 239584
rect 269356 239572 269362 239624
rect 278056 239612 278084 239720
rect 278406 239708 278412 239760
rect 278464 239748 278470 239760
rect 299290 239748 299296 239760
rect 278464 239720 299296 239748
rect 278464 239708 278470 239720
rect 299290 239708 299296 239720
rect 299348 239708 299354 239760
rect 278130 239640 278136 239692
rect 278188 239680 278194 239692
rect 292206 239680 292212 239692
rect 278188 239652 292212 239680
rect 278188 239640 278194 239652
rect 292206 239640 292212 239652
rect 292264 239640 292270 239692
rect 278406 239612 278412 239624
rect 278056 239584 278412 239612
rect 278406 239572 278412 239584
rect 278464 239572 278470 239624
rect 265802 239544 265808 239556
rect 265314 239516 265808 239544
rect 265802 239504 265808 239516
rect 265860 239504 265866 239556
rect 266078 239504 266084 239556
rect 266136 239544 266142 239556
rect 268194 239544 268200 239556
rect 266136 239516 268200 239544
rect 266136 239504 266142 239516
rect 268194 239504 268200 239516
rect 268252 239504 268258 239556
rect 286962 239504 286968 239556
rect 287020 239544 287026 239556
rect 311434 239544 311440 239556
rect 287020 239516 311440 239544
rect 287020 239504 287026 239516
rect 311434 239504 311440 239516
rect 311492 239504 311498 239556
rect 248322 239436 248328 239488
rect 248380 239476 248386 239488
rect 260742 239476 260748 239488
rect 248380 239448 260748 239476
rect 248380 239436 248386 239448
rect 260742 239436 260748 239448
rect 260800 239436 260806 239488
rect 263594 239436 263600 239488
rect 263652 239476 263658 239488
rect 264974 239476 264980 239488
rect 263652 239448 264980 239476
rect 263652 239436 263658 239448
rect 264974 239436 264980 239448
rect 265032 239436 265038 239488
rect 265222 239448 265256 239488
rect 265250 239436 265256 239448
rect 265308 239436 265314 239488
rect 266630 239436 266636 239488
rect 266688 239476 266694 239488
rect 273254 239476 273260 239488
rect 266688 239448 273260 239476
rect 266688 239436 266694 239448
rect 273254 239436 273260 239448
rect 273312 239436 273318 239488
rect 278130 239436 278136 239488
rect 278188 239476 278194 239488
rect 305822 239476 305828 239488
rect 278188 239448 305828 239476
rect 278188 239436 278194 239448
rect 305822 239436 305828 239448
rect 305880 239436 305886 239488
rect 247460 239380 247816 239408
rect 247460 239368 247466 239380
rect 249058 239368 249064 239420
rect 249116 239408 249122 239420
rect 285306 239408 285312 239420
rect 249116 239380 285312 239408
rect 249116 239368 249122 239380
rect 285306 239368 285312 239380
rect 285364 239368 285370 239420
rect 302142 239368 302148 239420
rect 302200 239408 302206 239420
rect 348786 239408 348792 239420
rect 302200 239380 348792 239408
rect 302200 239368 302206 239380
rect 348786 239368 348792 239380
rect 348844 239408 348850 239420
rect 558914 239408 558920 239420
rect 348844 239380 558920 239408
rect 348844 239368 348850 239380
rect 558914 239368 558920 239380
rect 558972 239368 558978 239420
rect 227438 239340 227444 239352
rect 225196 239312 225368 239340
rect 225432 239312 227444 239340
rect 225196 239300 225202 239312
rect 152918 239232 152924 239284
rect 152976 239272 152982 239284
rect 152976 239244 224770 239272
rect 152976 239232 152982 239244
rect 154114 239164 154120 239216
rect 154172 239204 154178 239216
rect 224218 239204 224224 239216
rect 154172 239176 224224 239204
rect 154172 239164 154178 239176
rect 224218 239164 224224 239176
rect 224276 239204 224282 239216
rect 224402 239204 224408 239216
rect 224276 239176 224408 239204
rect 224276 239164 224282 239176
rect 224402 239164 224408 239176
rect 224460 239164 224466 239216
rect 224742 239204 224770 239244
rect 224954 239232 224960 239284
rect 225012 239272 225018 239284
rect 225230 239272 225236 239284
rect 225012 239244 225236 239272
rect 225012 239232 225018 239244
rect 225230 239232 225236 239244
rect 225288 239232 225294 239284
rect 225340 239272 225368 239312
rect 227438 239300 227444 239312
rect 227496 239300 227502 239352
rect 232222 239300 232228 239352
rect 232280 239340 232286 239352
rect 280706 239340 280712 239352
rect 232280 239312 280712 239340
rect 232280 239300 232286 239312
rect 280706 239300 280712 239312
rect 280764 239300 280770 239352
rect 226610 239272 226616 239284
rect 225340 239244 226616 239272
rect 226610 239232 226616 239244
rect 226668 239232 226674 239284
rect 227162 239232 227168 239284
rect 227220 239272 227226 239284
rect 228542 239272 228548 239284
rect 227220 239244 228548 239272
rect 227220 239232 227226 239244
rect 228542 239232 228548 239244
rect 228600 239232 228606 239284
rect 229278 239232 229284 239284
rect 229336 239272 229342 239284
rect 231302 239272 231308 239284
rect 229336 239244 231308 239272
rect 229336 239232 229342 239244
rect 231302 239232 231308 239244
rect 231360 239232 231366 239284
rect 231670 239232 231676 239284
rect 231728 239272 231734 239284
rect 248046 239272 248052 239284
rect 231728 239244 248052 239272
rect 231728 239232 231734 239244
rect 248046 239232 248052 239244
rect 248104 239232 248110 239284
rect 250530 239232 250536 239284
rect 250588 239272 250594 239284
rect 282086 239272 282092 239284
rect 250588 239244 282092 239272
rect 250588 239232 250594 239244
rect 282086 239232 282092 239244
rect 282144 239232 282150 239284
rect 224742 239176 227714 239204
rect 221476 239108 223758 239136
rect 212994 239028 213000 239080
rect 213052 239068 213058 239080
rect 216214 239068 216220 239080
rect 213052 239040 216220 239068
rect 213052 239028 213058 239040
rect 216214 239028 216220 239040
rect 216272 239068 216278 239080
rect 221476 239068 221504 239108
rect 216272 239040 221504 239068
rect 223730 239068 223758 239108
rect 224678 239096 224684 239148
rect 224736 239136 224742 239148
rect 225874 239136 225880 239148
rect 224736 239108 225880 239136
rect 224736 239096 224742 239108
rect 225874 239096 225880 239108
rect 225932 239096 225938 239148
rect 227686 239136 227714 239176
rect 227990 239164 227996 239216
rect 228048 239204 228054 239216
rect 282914 239204 282920 239216
rect 228048 239176 282920 239204
rect 228048 239164 228054 239176
rect 282914 239164 282920 239176
rect 282972 239164 282978 239216
rect 228818 239136 228824 239148
rect 227686 239108 228824 239136
rect 228818 239096 228824 239108
rect 228876 239136 228882 239148
rect 231670 239136 231676 239148
rect 228876 239108 231676 239136
rect 228876 239096 228882 239108
rect 231670 239096 231676 239108
rect 231728 239096 231734 239148
rect 233050 239096 233056 239148
rect 233108 239136 233114 239148
rect 233108 239108 234844 239136
rect 233108 239096 233114 239108
rect 234706 239068 234712 239080
rect 223730 239040 234712 239068
rect 216272 239028 216278 239040
rect 234706 239028 234712 239040
rect 234764 239028 234770 239080
rect 234816 239068 234844 239108
rect 234982 239096 234988 239148
rect 235040 239136 235046 239148
rect 248322 239136 248328 239148
rect 235040 239108 248328 239136
rect 235040 239096 235046 239108
rect 248322 239096 248328 239108
rect 248380 239096 248386 239148
rect 248506 239096 248512 239148
rect 248564 239136 248570 239148
rect 292666 239136 292672 239148
rect 248564 239108 292672 239136
rect 248564 239096 248570 239108
rect 292666 239096 292672 239108
rect 292724 239096 292730 239148
rect 237006 239068 237012 239080
rect 234816 239040 237012 239068
rect 237006 239028 237012 239040
rect 237064 239028 237070 239080
rect 237834 239028 237840 239080
rect 237892 239068 237898 239080
rect 297818 239068 297824 239080
rect 237892 239040 297824 239068
rect 237892 239028 237898 239040
rect 297818 239028 297824 239040
rect 297876 239028 297882 239080
rect 215846 238960 215852 239012
rect 215904 239000 215910 239012
rect 225138 239000 225144 239012
rect 215904 238972 225144 239000
rect 215904 238960 215910 238972
rect 225138 238960 225144 238972
rect 225196 238960 225202 239012
rect 226058 238960 226064 239012
rect 226116 239000 226122 239012
rect 228082 239000 228088 239012
rect 226116 238972 228088 239000
rect 226116 238960 226122 238972
rect 228082 238960 228088 238972
rect 228140 238960 228146 239012
rect 229738 238960 229744 239012
rect 229796 239000 229802 239012
rect 229796 238972 235120 239000
rect 229796 238960 229802 238972
rect 220262 238892 220268 238944
rect 220320 238932 220326 238944
rect 230658 238932 230664 238944
rect 220320 238904 230664 238932
rect 220320 238892 220326 238904
rect 230658 238892 230664 238904
rect 230716 238892 230722 238944
rect 230842 238892 230848 238944
rect 230900 238932 230906 238944
rect 231486 238932 231492 238944
rect 230900 238904 231492 238932
rect 230900 238892 230906 238904
rect 231486 238892 231492 238904
rect 231544 238892 231550 238944
rect 232406 238892 232412 238944
rect 232464 238932 232470 238944
rect 234982 238932 234988 238944
rect 232464 238904 234988 238932
rect 232464 238892 232470 238904
rect 234982 238892 234988 238904
rect 235040 238892 235046 238944
rect 235092 238932 235120 238972
rect 237558 238960 237564 239012
rect 237616 239000 237622 239012
rect 297634 239000 297640 239012
rect 237616 238972 297640 239000
rect 237616 238960 237622 238972
rect 297634 238960 297640 238972
rect 297692 238960 297698 239012
rect 238754 238932 238760 238944
rect 235092 238904 238760 238932
rect 238754 238892 238760 238904
rect 238812 238932 238818 238944
rect 240594 238932 240600 238944
rect 238812 238904 240600 238932
rect 238812 238892 238818 238904
rect 240594 238892 240600 238904
rect 240652 238892 240658 238944
rect 248506 238932 248512 238944
rect 242452 238904 248512 238932
rect 217594 238824 217600 238876
rect 217652 238864 217658 238876
rect 220722 238864 220728 238876
rect 217652 238836 220728 238864
rect 217652 238824 217658 238836
rect 220722 238824 220728 238836
rect 220780 238824 220786 238876
rect 222102 238824 222108 238876
rect 222160 238864 222166 238876
rect 240226 238864 240232 238876
rect 222160 238836 240232 238864
rect 222160 238824 222166 238836
rect 240226 238824 240232 238836
rect 240284 238824 240290 238876
rect 220354 238756 220360 238808
rect 220412 238796 220418 238808
rect 233050 238796 233056 238808
rect 220412 238768 233056 238796
rect 220412 238756 220418 238768
rect 233050 238756 233056 238768
rect 233108 238756 233114 238808
rect 233234 238756 233240 238808
rect 233292 238796 233298 238808
rect 242452 238796 242480 238904
rect 248506 238892 248512 238904
rect 248564 238892 248570 238944
rect 249242 238892 249248 238944
rect 249300 238932 249306 238944
rect 305914 238932 305920 238944
rect 249300 238904 305920 238932
rect 249300 238892 249306 238904
rect 305914 238892 305920 238904
rect 305972 238892 305978 238944
rect 246482 238824 246488 238876
rect 246540 238864 246546 238876
rect 262766 238864 262772 238876
rect 246540 238836 262772 238864
rect 246540 238824 246546 238836
rect 262766 238824 262772 238836
rect 262824 238824 262830 238876
rect 269574 238864 269580 238876
rect 263612 238836 269580 238864
rect 233292 238768 242480 238796
rect 233292 238756 233298 238768
rect 245286 238756 245292 238808
rect 245344 238796 245350 238808
rect 245838 238796 245844 238808
rect 245344 238768 245844 238796
rect 245344 238756 245350 238768
rect 245838 238756 245844 238768
rect 245896 238756 245902 238808
rect 247310 238756 247316 238808
rect 247368 238796 247374 238808
rect 262950 238796 262956 238808
rect 247368 238768 262956 238796
rect 247368 238756 247374 238768
rect 262950 238756 262956 238768
rect 263008 238756 263014 238808
rect 209222 238688 209228 238740
rect 209280 238728 209286 238740
rect 223758 238728 223764 238740
rect 209280 238700 223764 238728
rect 209280 238688 209286 238700
rect 223758 238688 223764 238700
rect 223816 238688 223822 238740
rect 224218 238688 224224 238740
rect 224276 238728 224282 238740
rect 226702 238728 226708 238740
rect 224276 238700 226708 238728
rect 224276 238688 224282 238700
rect 226702 238688 226708 238700
rect 226760 238688 226766 238740
rect 230014 238688 230020 238740
rect 230072 238728 230078 238740
rect 230072 238700 232544 238728
rect 230072 238688 230078 238700
rect 222838 238620 222844 238672
rect 222896 238660 222902 238672
rect 232406 238660 232412 238672
rect 222896 238632 232412 238660
rect 222896 238620 222902 238632
rect 232406 238620 232412 238632
rect 232464 238620 232470 238672
rect 232516 238660 232544 238700
rect 233510 238688 233516 238740
rect 233568 238728 233574 238740
rect 233786 238728 233792 238740
rect 233568 238700 233792 238728
rect 233568 238688 233574 238700
rect 233786 238688 233792 238700
rect 233844 238688 233850 238740
rect 236178 238728 236184 238740
rect 233896 238700 236184 238728
rect 233896 238660 233924 238700
rect 236178 238688 236184 238700
rect 236236 238688 236242 238740
rect 240962 238728 240968 238740
rect 237024 238700 240968 238728
rect 232516 238632 233924 238660
rect 234982 238620 234988 238672
rect 235040 238660 235046 238672
rect 237024 238660 237052 238700
rect 240962 238688 240968 238700
rect 241020 238688 241026 238740
rect 245194 238688 245200 238740
rect 245252 238728 245258 238740
rect 249242 238728 249248 238740
rect 245252 238700 249248 238728
rect 245252 238688 245258 238700
rect 249242 238688 249248 238700
rect 249300 238688 249306 238740
rect 250898 238688 250904 238740
rect 250956 238728 250962 238740
rect 251174 238728 251180 238740
rect 250956 238700 251180 238728
rect 250956 238688 250962 238700
rect 251174 238688 251180 238700
rect 251232 238688 251238 238740
rect 257154 238688 257160 238740
rect 257212 238728 257218 238740
rect 257890 238728 257896 238740
rect 257212 238700 257896 238728
rect 257212 238688 257218 238700
rect 257890 238688 257896 238700
rect 257948 238688 257954 238740
rect 260466 238688 260472 238740
rect 260524 238728 260530 238740
rect 263612 238728 263640 238836
rect 269574 238824 269580 238836
rect 269632 238824 269638 238876
rect 296622 238824 296628 238876
rect 296680 238864 296686 238876
rect 506474 238864 506480 238876
rect 296680 238836 506480 238864
rect 296680 238824 296686 238836
rect 506474 238824 506480 238836
rect 506532 238824 506538 238876
rect 264974 238756 264980 238808
rect 265032 238796 265038 238808
rect 278130 238796 278136 238808
rect 265032 238768 278136 238796
rect 265032 238756 265038 238768
rect 278130 238756 278136 238768
rect 278188 238756 278194 238808
rect 296530 238756 296536 238808
rect 296588 238796 296594 238808
rect 540974 238796 540980 238808
rect 296588 238768 540980 238796
rect 296588 238756 296594 238768
rect 540974 238756 540980 238768
rect 541032 238756 541038 238808
rect 260524 238700 263640 238728
rect 260524 238688 260530 238700
rect 264422 238688 264428 238740
rect 264480 238728 264486 238740
rect 269206 238728 269212 238740
rect 264480 238700 269212 238728
rect 264480 238688 264486 238700
rect 269206 238688 269212 238700
rect 269264 238688 269270 238740
rect 235040 238632 237052 238660
rect 235040 238620 235046 238632
rect 240226 238620 240232 238672
rect 240284 238660 240290 238672
rect 249058 238660 249064 238672
rect 240284 238632 249064 238660
rect 240284 238620 240290 238632
rect 249058 238620 249064 238632
rect 249116 238620 249122 238672
rect 249426 238620 249432 238672
rect 249484 238660 249490 238672
rect 251450 238660 251456 238672
rect 249484 238632 251456 238660
rect 249484 238620 249490 238632
rect 251450 238620 251456 238632
rect 251508 238620 251514 238672
rect 251818 238620 251824 238672
rect 251876 238660 251882 238672
rect 258810 238660 258816 238672
rect 251876 238632 258816 238660
rect 251876 238620 251882 238632
rect 258810 238620 258816 238632
rect 258868 238620 258874 238672
rect 270954 238660 270960 238672
rect 258920 238632 270960 238660
rect 207750 238552 207756 238604
rect 207808 238592 207814 238604
rect 231854 238592 231860 238604
rect 207808 238564 231860 238592
rect 207808 238552 207814 238564
rect 231854 238552 231860 238564
rect 231912 238552 231918 238604
rect 232774 238552 232780 238604
rect 232832 238592 232838 238604
rect 239582 238592 239588 238604
rect 232832 238564 239588 238592
rect 232832 238552 232838 238564
rect 239582 238552 239588 238564
rect 239640 238552 239646 238604
rect 250162 238552 250168 238604
rect 250220 238592 250226 238604
rect 251266 238592 251272 238604
rect 250220 238564 251272 238592
rect 250220 238552 250226 238564
rect 251266 238552 251272 238564
rect 251324 238552 251330 238604
rect 252002 238552 252008 238604
rect 252060 238592 252066 238604
rect 258920 238592 258948 238632
rect 270954 238620 270960 238632
rect 271012 238620 271018 238672
rect 271046 238620 271052 238672
rect 271104 238660 271110 238672
rect 312446 238660 312452 238672
rect 271104 238632 312452 238660
rect 271104 238620 271110 238632
rect 312446 238620 312452 238632
rect 312504 238620 312510 238672
rect 252060 238564 258948 238592
rect 252060 238552 252066 238564
rect 261294 238552 261300 238604
rect 261352 238592 261358 238604
rect 264422 238592 264428 238604
rect 261352 238564 264428 238592
rect 261352 238552 261358 238564
rect 264422 238552 264428 238564
rect 264480 238552 264486 238604
rect 265986 238552 265992 238604
rect 266044 238592 266050 238604
rect 270862 238592 270868 238604
rect 266044 238564 270868 238592
rect 266044 238552 266050 238564
rect 270862 238552 270868 238564
rect 270920 238552 270926 238604
rect 210326 238484 210332 238536
rect 210384 238524 210390 238536
rect 226518 238524 226524 238536
rect 210384 238496 226524 238524
rect 210384 238484 210390 238496
rect 226518 238484 226524 238496
rect 226576 238484 226582 238536
rect 228818 238484 228824 238536
rect 228876 238524 228882 238536
rect 231210 238524 231216 238536
rect 228876 238496 231216 238524
rect 228876 238484 228882 238496
rect 231210 238484 231216 238496
rect 231268 238484 231274 238536
rect 232130 238484 232136 238536
rect 232188 238524 232194 238536
rect 233050 238524 233056 238536
rect 232188 238496 233056 238524
rect 232188 238484 232194 238496
rect 233050 238484 233056 238496
rect 233108 238484 233114 238536
rect 233234 238484 233240 238536
rect 233292 238524 233298 238536
rect 268562 238524 268568 238536
rect 233292 238496 268568 238524
rect 233292 238484 233298 238496
rect 268562 238484 268568 238496
rect 268620 238484 268626 238536
rect 209314 238416 209320 238468
rect 209372 238456 209378 238468
rect 222562 238456 222568 238468
rect 209372 238428 222568 238456
rect 209372 238416 209378 238428
rect 222562 238416 222568 238428
rect 222620 238416 222626 238468
rect 222838 238416 222844 238468
rect 222896 238456 222902 238468
rect 230198 238456 230204 238468
rect 222896 238428 230204 238456
rect 222896 238416 222902 238428
rect 230198 238416 230204 238428
rect 230256 238416 230262 238468
rect 230658 238416 230664 238468
rect 230716 238456 230722 238468
rect 267274 238456 267280 238468
rect 230716 238428 267280 238456
rect 230716 238416 230722 238428
rect 267274 238416 267280 238428
rect 267332 238416 267338 238468
rect 269298 238416 269304 238468
rect 269356 238456 269362 238468
rect 271506 238456 271512 238468
rect 269356 238428 271512 238456
rect 269356 238416 269362 238428
rect 271506 238416 271512 238428
rect 271564 238416 271570 238468
rect 192478 238348 192484 238400
rect 192536 238388 192542 238400
rect 223574 238388 223580 238400
rect 192536 238360 223580 238388
rect 192536 238348 192542 238360
rect 223574 238348 223580 238360
rect 223632 238348 223638 238400
rect 225322 238348 225328 238400
rect 225380 238388 225386 238400
rect 225782 238388 225788 238400
rect 225380 238360 225788 238388
rect 225380 238348 225386 238360
rect 225782 238348 225788 238360
rect 225840 238348 225846 238400
rect 226518 238348 226524 238400
rect 226576 238388 226582 238400
rect 227346 238388 227352 238400
rect 226576 238360 227352 238388
rect 226576 238348 226582 238360
rect 227346 238348 227352 238360
rect 227404 238348 227410 238400
rect 228450 238348 228456 238400
rect 228508 238388 228514 238400
rect 229094 238388 229100 238400
rect 228508 238360 229100 238388
rect 228508 238348 228514 238360
rect 229094 238348 229100 238360
rect 229152 238348 229158 238400
rect 231946 238348 231952 238400
rect 232004 238388 232010 238400
rect 237098 238388 237104 238400
rect 232004 238360 237104 238388
rect 232004 238348 232010 238360
rect 237098 238348 237104 238360
rect 237156 238348 237162 238400
rect 239214 238348 239220 238400
rect 239272 238388 239278 238400
rect 239582 238388 239588 238400
rect 239272 238360 239588 238388
rect 239272 238348 239278 238360
rect 239582 238348 239588 238360
rect 239640 238348 239646 238400
rect 270770 238388 270776 238400
rect 239692 238360 270776 238388
rect 191650 238280 191656 238332
rect 191708 238320 191714 238332
rect 222746 238320 222752 238332
rect 191708 238292 222752 238320
rect 191708 238280 191714 238292
rect 222746 238280 222752 238292
rect 222804 238280 222810 238332
rect 225414 238320 225420 238332
rect 223546 238292 225420 238320
rect 194318 238212 194324 238264
rect 194376 238252 194382 238264
rect 223546 238252 223574 238292
rect 225414 238280 225420 238292
rect 225472 238280 225478 238332
rect 227438 238280 227444 238332
rect 227496 238320 227502 238332
rect 229830 238320 229836 238332
rect 227496 238292 229836 238320
rect 227496 238280 227502 238292
rect 229830 238280 229836 238292
rect 229888 238280 229894 238332
rect 230382 238280 230388 238332
rect 230440 238320 230446 238332
rect 233234 238320 233240 238332
rect 230440 238292 233240 238320
rect 230440 238280 230446 238292
rect 233234 238280 233240 238292
rect 233292 238280 233298 238332
rect 233418 238280 233424 238332
rect 233476 238320 233482 238332
rect 239692 238320 239720 238360
rect 270770 238348 270776 238360
rect 270828 238348 270834 238400
rect 268838 238320 268844 238332
rect 233476 238292 239720 238320
rect 239784 238292 268844 238320
rect 233476 238280 233482 238292
rect 194376 238224 223574 238252
rect 194376 238212 194382 238224
rect 225322 238212 225328 238264
rect 225380 238252 225386 238264
rect 227898 238252 227904 238264
rect 225380 238224 227904 238252
rect 225380 238212 225386 238224
rect 227898 238212 227904 238224
rect 227956 238212 227962 238264
rect 229186 238212 229192 238264
rect 229244 238252 229250 238264
rect 229646 238252 229652 238264
rect 229244 238224 229652 238252
rect 229244 238212 229250 238224
rect 229646 238212 229652 238224
rect 229704 238212 229710 238264
rect 231486 238212 231492 238264
rect 231544 238252 231550 238264
rect 239784 238252 239812 238292
rect 268838 238280 268844 238292
rect 268896 238280 268902 238332
rect 267366 238252 267372 238264
rect 231544 238224 239812 238252
rect 252526 238224 264100 238252
rect 231544 238212 231550 238224
rect 182910 238144 182916 238196
rect 182968 238184 182974 238196
rect 218974 238184 218980 238196
rect 182968 238156 218980 238184
rect 182968 238144 182974 238156
rect 218974 238144 218980 238156
rect 219032 238144 219038 238196
rect 222562 238144 222568 238196
rect 222620 238184 222626 238196
rect 225690 238184 225696 238196
rect 222620 238156 225696 238184
rect 222620 238144 222626 238156
rect 225690 238144 225696 238156
rect 225748 238144 225754 238196
rect 225874 238144 225880 238196
rect 225932 238184 225938 238196
rect 226978 238184 226984 238196
rect 225932 238156 226984 238184
rect 225932 238144 225938 238156
rect 226978 238144 226984 238156
rect 227036 238144 227042 238196
rect 227806 238144 227812 238196
rect 227864 238184 227870 238196
rect 231946 238184 231952 238196
rect 227864 238156 231952 238184
rect 227864 238144 227870 238156
rect 231946 238144 231952 238156
rect 232004 238144 232010 238196
rect 233050 238144 233056 238196
rect 233108 238184 233114 238196
rect 252526 238184 252554 238224
rect 233108 238156 252554 238184
rect 233108 238144 233114 238156
rect 259822 238144 259828 238196
rect 259880 238184 259886 238196
rect 263870 238184 263876 238196
rect 259880 238156 263876 238184
rect 259880 238144 259886 238156
rect 263870 238144 263876 238156
rect 263928 238144 263934 238196
rect 161290 238076 161296 238128
rect 161348 238116 161354 238128
rect 215938 238116 215944 238128
rect 161348 238088 215944 238116
rect 161348 238076 161354 238088
rect 215938 238076 215944 238088
rect 215996 238116 216002 238128
rect 216582 238116 216588 238128
rect 215996 238088 216588 238116
rect 215996 238076 216002 238088
rect 216582 238076 216588 238088
rect 216640 238076 216646 238128
rect 225598 238076 225604 238128
rect 225656 238116 225662 238128
rect 231670 238116 231676 238128
rect 225656 238088 231676 238116
rect 225656 238076 225662 238088
rect 231670 238076 231676 238088
rect 231728 238076 231734 238128
rect 231762 238076 231768 238128
rect 231820 238116 231826 238128
rect 247678 238116 247684 238128
rect 231820 238088 247684 238116
rect 231820 238076 231826 238088
rect 247678 238076 247684 238088
rect 247736 238076 247742 238128
rect 264072 238116 264100 238224
rect 265728 238224 267372 238252
rect 265728 238116 265756 238224
rect 267366 238212 267372 238224
rect 267424 238212 267430 238264
rect 267734 238212 267740 238264
rect 267792 238252 267798 238264
rect 268378 238252 268384 238264
rect 267792 238224 268384 238252
rect 267792 238212 267798 238224
rect 268378 238212 268384 238224
rect 268436 238212 268442 238264
rect 268470 238144 268476 238196
rect 268528 238184 268534 238196
rect 319622 238184 319628 238196
rect 268528 238156 319628 238184
rect 268528 238144 268534 238156
rect 319622 238144 319628 238156
rect 319680 238144 319686 238196
rect 264072 238088 265756 238116
rect 265802 238076 265808 238128
rect 265860 238116 265866 238128
rect 322934 238116 322940 238128
rect 265860 238088 322940 238116
rect 265860 238076 265866 238088
rect 322934 238076 322940 238088
rect 322992 238076 322998 238128
rect 161198 238008 161204 238060
rect 161256 238048 161262 238060
rect 238478 238048 238484 238060
rect 161256 238020 238484 238048
rect 161256 238008 161262 238020
rect 238478 238008 238484 238020
rect 238536 238008 238542 238060
rect 239214 238008 239220 238060
rect 239272 238048 239278 238060
rect 239398 238048 239404 238060
rect 239272 238020 239404 238048
rect 239272 238008 239278 238020
rect 239398 238008 239404 238020
rect 239456 238008 239462 238060
rect 242894 238008 242900 238060
rect 242952 238048 242958 238060
rect 245010 238048 245016 238060
rect 242952 238020 245016 238048
rect 242952 238008 242958 238020
rect 245010 238008 245016 238020
rect 245068 238048 245074 238060
rect 246574 238048 246580 238060
rect 245068 238020 246580 238048
rect 245068 238008 245074 238020
rect 246574 238008 246580 238020
rect 246632 238008 246638 238060
rect 268010 238008 268016 238060
rect 268068 238048 268074 238060
rect 335538 238048 335544 238060
rect 268068 238020 335544 238048
rect 268068 238008 268074 238020
rect 335538 238008 335544 238020
rect 335596 238008 335602 238060
rect 221458 237940 221464 237992
rect 221516 237980 221522 237992
rect 232314 237980 232320 237992
rect 221516 237952 232320 237980
rect 221516 237940 221522 237952
rect 232314 237940 232320 237952
rect 232372 237940 232378 237992
rect 236270 237940 236276 237992
rect 236328 237980 236334 237992
rect 236914 237980 236920 237992
rect 236328 237952 236920 237980
rect 236328 237940 236334 237952
rect 236914 237940 236920 237952
rect 236972 237940 236978 237992
rect 238496 237980 238524 238008
rect 246390 237980 246396 237992
rect 238496 237952 246396 237980
rect 246390 237940 246396 237952
rect 246448 237940 246454 237992
rect 247126 237940 247132 237992
rect 247184 237980 247190 237992
rect 262030 237980 262036 237992
rect 247184 237952 262036 237980
rect 247184 237940 247190 237952
rect 262030 237940 262036 237952
rect 262088 237940 262094 237992
rect 266630 237940 266636 237992
rect 266688 237980 266694 237992
rect 266814 237980 266820 237992
rect 266688 237952 266820 237980
rect 266688 237940 266694 237952
rect 266814 237940 266820 237952
rect 266872 237940 266878 237992
rect 267550 237940 267556 237992
rect 267608 237980 267614 237992
rect 268562 237980 268568 237992
rect 267608 237952 268568 237980
rect 267608 237940 267614 237952
rect 268562 237940 268568 237952
rect 268620 237940 268626 237992
rect 268746 237940 268752 237992
rect 268804 237980 268810 237992
rect 304718 237980 304724 237992
rect 268804 237952 304724 237980
rect 268804 237940 268810 237952
rect 304718 237940 304724 237952
rect 304776 237940 304782 237992
rect 225138 237872 225144 237924
rect 225196 237912 225202 237924
rect 238938 237912 238944 237924
rect 225196 237884 238944 237912
rect 225196 237872 225202 237884
rect 238938 237872 238944 237884
rect 238996 237872 239002 237924
rect 239858 237872 239864 237924
rect 239916 237912 239922 237924
rect 241606 237912 241612 237924
rect 239916 237884 241612 237912
rect 239916 237872 239922 237884
rect 241606 237872 241612 237884
rect 241664 237872 241670 237924
rect 243722 237872 243728 237924
rect 243780 237912 243786 237924
rect 258902 237912 258908 237924
rect 243780 237884 258908 237912
rect 243780 237872 243786 237884
rect 258902 237872 258908 237884
rect 258960 237872 258966 237924
rect 259730 237872 259736 237924
rect 259788 237912 259794 237924
rect 269114 237912 269120 237924
rect 259788 237884 269120 237912
rect 259788 237872 259794 237884
rect 269114 237872 269120 237884
rect 269172 237872 269178 237924
rect 270310 237872 270316 237924
rect 270368 237912 270374 237924
rect 275738 237912 275744 237924
rect 270368 237884 275744 237912
rect 270368 237872 270374 237884
rect 275738 237872 275744 237884
rect 275796 237872 275802 237924
rect 216582 237804 216588 237856
rect 216640 237844 216646 237856
rect 229094 237844 229100 237856
rect 216640 237816 229100 237844
rect 216640 237804 216646 237816
rect 229094 237804 229100 237816
rect 229152 237804 229158 237856
rect 235718 237844 235724 237856
rect 229848 237816 235724 237844
rect 216306 237736 216312 237788
rect 216364 237776 216370 237788
rect 229848 237776 229876 237816
rect 235718 237804 235724 237816
rect 235776 237804 235782 237856
rect 236270 237804 236276 237856
rect 236328 237844 236334 237856
rect 236454 237844 236460 237856
rect 236328 237816 236460 237844
rect 236328 237804 236334 237816
rect 236454 237804 236460 237816
rect 236512 237804 236518 237856
rect 254302 237804 254308 237856
rect 254360 237844 254366 237856
rect 260466 237844 260472 237856
rect 254360 237816 260472 237844
rect 254360 237804 254366 237816
rect 260466 237804 260472 237816
rect 260524 237804 260530 237856
rect 263870 237804 263876 237856
rect 263928 237844 263934 237856
rect 270586 237844 270592 237856
rect 263928 237816 270592 237844
rect 263928 237804 263934 237816
rect 270586 237804 270592 237816
rect 270644 237844 270650 237856
rect 272058 237844 272064 237856
rect 270644 237816 272064 237844
rect 270644 237804 270650 237816
rect 272058 237804 272064 237816
rect 272116 237804 272122 237856
rect 216364 237748 229876 237776
rect 216364 237736 216370 237748
rect 229922 237736 229928 237788
rect 229980 237776 229986 237788
rect 233418 237776 233424 237788
rect 229980 237748 233424 237776
rect 229980 237736 229986 237748
rect 233418 237736 233424 237748
rect 233476 237736 233482 237788
rect 253934 237736 253940 237788
rect 253992 237776 253998 237788
rect 271230 237776 271236 237788
rect 253992 237748 271236 237776
rect 253992 237736 253998 237748
rect 271230 237736 271236 237748
rect 271288 237736 271294 237788
rect 231854 237668 231860 237720
rect 231912 237708 231918 237720
rect 231912 237680 237374 237708
rect 231912 237668 231918 237680
rect 224494 237600 224500 237652
rect 224552 237640 224558 237652
rect 235166 237640 235172 237652
rect 224552 237612 235172 237640
rect 224552 237600 224558 237612
rect 235166 237600 235172 237612
rect 235224 237600 235230 237652
rect 237346 237640 237374 237680
rect 257982 237668 257988 237720
rect 258040 237708 258046 237720
rect 259914 237708 259920 237720
rect 258040 237680 259920 237708
rect 258040 237668 258046 237680
rect 259914 237668 259920 237680
rect 259972 237668 259978 237720
rect 264054 237668 264060 237720
rect 264112 237708 264118 237720
rect 270310 237708 270316 237720
rect 264112 237680 270316 237708
rect 264112 237668 264118 237680
rect 270310 237668 270316 237680
rect 270368 237668 270374 237720
rect 271598 237640 271604 237652
rect 237346 237612 271604 237640
rect 271598 237600 271604 237612
rect 271656 237600 271662 237652
rect 231578 237572 231584 237584
rect 227686 237544 231584 237572
rect 162302 237396 162308 237448
rect 162360 237436 162366 237448
rect 227686 237436 227714 237544
rect 231578 237532 231584 237544
rect 231636 237532 231642 237584
rect 231670 237532 231676 237584
rect 231728 237572 231734 237584
rect 269482 237572 269488 237584
rect 231728 237544 269488 237572
rect 231728 237532 231734 237544
rect 269482 237532 269488 237544
rect 269540 237532 269546 237584
rect 230566 237464 230572 237516
rect 230624 237504 230630 237516
rect 269390 237504 269396 237516
rect 230624 237476 269396 237504
rect 230624 237464 230630 237476
rect 269390 237464 269396 237476
rect 269448 237464 269454 237516
rect 162360 237408 227714 237436
rect 162360 237396 162366 237408
rect 229370 237396 229376 237448
rect 229428 237436 229434 237448
rect 229554 237436 229560 237448
rect 229428 237408 229560 237436
rect 229428 237396 229434 237408
rect 229554 237396 229560 237408
rect 229612 237436 229618 237448
rect 229922 237436 229928 237448
rect 229612 237408 229928 237436
rect 229612 237396 229618 237408
rect 229922 237396 229928 237408
rect 229980 237396 229986 237448
rect 231302 237396 231308 237448
rect 231360 237436 231366 237448
rect 231486 237436 231492 237448
rect 231360 237408 231492 237436
rect 231360 237396 231366 237408
rect 231486 237396 231492 237408
rect 231544 237396 231550 237448
rect 231578 237396 231584 237448
rect 231636 237436 231642 237448
rect 236914 237436 236920 237448
rect 231636 237408 236920 237436
rect 231636 237396 231642 237408
rect 236914 237396 236920 237408
rect 236972 237396 236978 237448
rect 252278 237396 252284 237448
rect 252336 237436 252342 237448
rect 252646 237436 252652 237448
rect 252336 237408 252652 237436
rect 252336 237396 252342 237408
rect 252646 237396 252652 237408
rect 252704 237436 252710 237448
rect 271046 237436 271052 237448
rect 252704 237408 271052 237436
rect 252704 237396 252710 237408
rect 271046 237396 271052 237408
rect 271104 237396 271110 237448
rect 281534 237396 281540 237448
rect 281592 237436 281598 237448
rect 284478 237436 284484 237448
rect 281592 237408 284484 237436
rect 281592 237396 281598 237408
rect 284478 237396 284484 237408
rect 284536 237396 284542 237448
rect 231946 237328 231952 237380
rect 232004 237368 232010 237380
rect 232222 237368 232228 237380
rect 232004 237340 232228 237368
rect 232004 237328 232010 237340
rect 232222 237328 232228 237340
rect 232280 237328 232286 237380
rect 267550 237328 267556 237380
rect 267608 237368 267614 237380
rect 267826 237368 267832 237380
rect 267608 237340 267832 237368
rect 267608 237328 267614 237340
rect 267826 237328 267832 237340
rect 267884 237328 267890 237380
rect 269114 237328 269120 237380
rect 269172 237368 269178 237380
rect 270402 237368 270408 237380
rect 269172 237340 270408 237368
rect 269172 237328 269178 237340
rect 270402 237328 270408 237340
rect 270460 237368 270466 237380
rect 281350 237368 281356 237380
rect 270460 237340 281356 237368
rect 270460 237328 270466 237340
rect 281350 237328 281356 237340
rect 281408 237328 281414 237380
rect 213454 237260 213460 237312
rect 213512 237300 213518 237312
rect 221642 237300 221648 237312
rect 213512 237272 221648 237300
rect 213512 237260 213518 237272
rect 221642 237260 221648 237272
rect 221700 237300 221706 237312
rect 255682 237300 255688 237312
rect 221700 237272 255688 237300
rect 221700 237260 221706 237272
rect 255682 237260 255688 237272
rect 255740 237260 255746 237312
rect 261478 237260 261484 237312
rect 261536 237300 261542 237312
rect 274634 237300 274640 237312
rect 261536 237272 274640 237300
rect 261536 237260 261542 237272
rect 274634 237260 274640 237272
rect 274692 237260 274698 237312
rect 276290 237260 276296 237312
rect 276348 237300 276354 237312
rect 277118 237300 277124 237312
rect 276348 237272 277124 237300
rect 276348 237260 276354 237272
rect 277118 237260 277124 237272
rect 277176 237260 277182 237312
rect 277394 237260 277400 237312
rect 277452 237300 277458 237312
rect 278498 237300 278504 237312
rect 277452 237272 278504 237300
rect 277452 237260 277458 237272
rect 278498 237260 278504 237272
rect 278556 237260 278562 237312
rect 205542 237192 205548 237244
rect 205600 237232 205606 237244
rect 224310 237232 224316 237244
rect 205600 237204 224316 237232
rect 205600 237192 205606 237204
rect 224310 237192 224316 237204
rect 224368 237192 224374 237244
rect 234890 237192 234896 237244
rect 234948 237232 234954 237244
rect 253290 237232 253296 237244
rect 234948 237204 253296 237232
rect 234948 237192 234954 237204
rect 253290 237192 253296 237204
rect 253348 237192 253354 237244
rect 254394 237192 254400 237244
rect 254452 237232 254458 237244
rect 294782 237232 294788 237244
rect 254452 237204 294788 237232
rect 254452 237192 254458 237204
rect 294782 237192 294788 237204
rect 294840 237192 294846 237244
rect 239858 237124 239864 237176
rect 239916 237164 239922 237176
rect 240042 237164 240048 237176
rect 239916 237136 240048 237164
rect 239916 237124 239922 237136
rect 240042 237124 240048 237136
rect 240100 237124 240106 237176
rect 252646 237124 252652 237176
rect 252704 237164 252710 237176
rect 253658 237164 253664 237176
rect 252704 237136 253664 237164
rect 252704 237124 252710 237136
rect 253658 237124 253664 237136
rect 253716 237124 253722 237176
rect 286594 237164 286600 237176
rect 258736 237136 286600 237164
rect 234798 237056 234804 237108
rect 234856 237096 234862 237108
rect 235626 237096 235632 237108
rect 234856 237068 235632 237096
rect 234856 237056 234862 237068
rect 235626 237056 235632 237068
rect 235684 237056 235690 237108
rect 237282 237056 237288 237108
rect 237340 237096 237346 237108
rect 241146 237096 241152 237108
rect 237340 237068 241152 237096
rect 237340 237056 237346 237068
rect 241146 237056 241152 237068
rect 241204 237056 241210 237108
rect 245654 237056 245660 237108
rect 245712 237096 245718 237108
rect 253290 237096 253296 237108
rect 245712 237068 253296 237096
rect 245712 237056 245718 237068
rect 253290 237056 253296 237068
rect 253348 237056 253354 237108
rect 253400 237068 258074 237096
rect 235902 237028 235908 237040
rect 215266 237000 235908 237028
rect 214834 236920 214840 236972
rect 214892 236960 214898 236972
rect 215266 236960 215294 237000
rect 235902 236988 235908 237000
rect 235960 236988 235966 237040
rect 239858 236988 239864 237040
rect 239916 237028 239922 237040
rect 240686 237028 240692 237040
rect 239916 237000 240692 237028
rect 239916 236988 239922 237000
rect 240686 236988 240692 237000
rect 240744 236988 240750 237040
rect 240778 236988 240784 237040
rect 240836 237028 240842 237040
rect 241054 237028 241060 237040
rect 240836 237000 241060 237028
rect 240836 236988 240842 237000
rect 241054 236988 241060 237000
rect 241112 236988 241118 237040
rect 246574 236988 246580 237040
rect 246632 237028 246638 237040
rect 253400 237028 253428 237068
rect 246632 237000 253428 237028
rect 246632 236988 246638 237000
rect 254394 236988 254400 237040
rect 254452 237028 254458 237040
rect 254854 237028 254860 237040
rect 254452 237000 254860 237028
rect 254452 236988 254458 237000
rect 254854 236988 254860 237000
rect 254912 236988 254918 237040
rect 258046 237028 258074 237068
rect 258736 237028 258764 237136
rect 286594 237124 286600 237136
rect 286652 237124 286658 237176
rect 277026 237096 277032 237108
rect 258046 237000 258764 237028
rect 258828 237068 277032 237096
rect 214892 236932 215294 236960
rect 214892 236920 214898 236932
rect 232498 236920 232504 236972
rect 232556 236960 232562 236972
rect 232682 236960 232688 236972
rect 232556 236932 232688 236960
rect 232556 236920 232562 236932
rect 232682 236920 232688 236932
rect 232740 236920 232746 236972
rect 235626 236920 235632 236972
rect 235684 236960 235690 236972
rect 252278 236960 252284 236972
rect 235684 236932 252284 236960
rect 235684 236920 235690 236932
rect 252278 236920 252284 236932
rect 252336 236920 252342 236972
rect 253290 236920 253296 236972
rect 253348 236960 253354 236972
rect 258828 236960 258856 237068
rect 277026 237056 277032 237068
rect 277084 237056 277090 237108
rect 259546 236988 259552 237040
rect 259604 237028 259610 237040
rect 260282 237028 260288 237040
rect 259604 237000 260288 237028
rect 259604 236988 259610 237000
rect 260282 236988 260288 237000
rect 260340 236988 260346 237040
rect 260466 236988 260472 237040
rect 260524 237028 260530 237040
rect 285858 237028 285864 237040
rect 260524 237000 285864 237028
rect 260524 236988 260530 237000
rect 285858 236988 285864 237000
rect 285916 236988 285922 237040
rect 253348 236932 258856 236960
rect 253348 236920 253354 236932
rect 258902 236920 258908 236972
rect 258960 236960 258966 236972
rect 268378 236960 268384 236972
rect 258960 236932 268384 236960
rect 258960 236920 258966 236932
rect 268378 236920 268384 236932
rect 268436 236920 268442 236972
rect 212166 236852 212172 236904
rect 212224 236892 212230 236904
rect 238110 236892 238116 236904
rect 212224 236864 238116 236892
rect 212224 236852 212230 236864
rect 238110 236852 238116 236864
rect 238168 236852 238174 236904
rect 240686 236852 240692 236904
rect 240744 236892 240750 236904
rect 241422 236892 241428 236904
rect 240744 236864 241428 236892
rect 240744 236852 240750 236864
rect 241422 236852 241428 236864
rect 241480 236852 241486 236904
rect 244550 236852 244556 236904
rect 244608 236892 244614 236904
rect 267826 236892 267832 236904
rect 244608 236864 267832 236892
rect 244608 236852 244614 236864
rect 267826 236852 267832 236864
rect 267884 236892 267890 236904
rect 287698 236892 287704 236904
rect 267884 236864 287704 236892
rect 267884 236852 267890 236864
rect 287698 236852 287704 236864
rect 287756 236852 287762 236904
rect 161382 236784 161388 236836
rect 161440 236824 161446 236836
rect 213270 236824 213276 236836
rect 161440 236796 213276 236824
rect 161440 236784 161446 236796
rect 213270 236784 213276 236796
rect 213328 236784 213334 236836
rect 214926 236784 214932 236836
rect 214984 236824 214990 236836
rect 253014 236824 253020 236836
rect 214984 236796 253020 236824
rect 214984 236784 214990 236796
rect 253014 236784 253020 236796
rect 253072 236824 253078 236836
rect 255866 236824 255872 236836
rect 253072 236796 255872 236824
rect 253072 236784 253078 236796
rect 255866 236784 255872 236796
rect 255924 236784 255930 236836
rect 276014 236784 276020 236836
rect 276072 236824 276078 236836
rect 296070 236824 296076 236836
rect 276072 236796 296076 236824
rect 276072 236784 276078 236796
rect 296070 236784 296076 236796
rect 296128 236824 296134 236836
rect 296128 236796 296714 236824
rect 296128 236784 296134 236796
rect 150342 236716 150348 236768
rect 150400 236756 150406 236768
rect 215110 236756 215116 236768
rect 150400 236728 215116 236756
rect 150400 236716 150406 236728
rect 215110 236716 215116 236728
rect 215168 236716 215174 236768
rect 221550 236716 221556 236768
rect 221608 236756 221614 236768
rect 244090 236756 244096 236768
rect 221608 236728 244096 236756
rect 221608 236716 221614 236728
rect 244090 236716 244096 236728
rect 244148 236756 244154 236768
rect 278774 236756 278780 236768
rect 244148 236728 278780 236756
rect 244148 236716 244154 236728
rect 278774 236716 278780 236728
rect 278832 236716 278838 236768
rect 296686 236756 296714 236796
rect 332870 236756 332876 236768
rect 296686 236728 332876 236756
rect 332870 236716 332876 236728
rect 332928 236716 332934 236768
rect 159818 236648 159824 236700
rect 159876 236688 159882 236700
rect 231946 236688 231952 236700
rect 159876 236660 231952 236688
rect 159876 236648 159882 236660
rect 231946 236648 231952 236660
rect 232004 236648 232010 236700
rect 242526 236648 242532 236700
rect 242584 236688 242590 236700
rect 243078 236688 243084 236700
rect 242584 236660 243084 236688
rect 242584 236648 242590 236660
rect 243078 236648 243084 236660
rect 243136 236648 243142 236700
rect 245194 236648 245200 236700
rect 245252 236688 245258 236700
rect 299658 236688 299664 236700
rect 245252 236660 299664 236688
rect 245252 236648 245258 236660
rect 299658 236648 299664 236660
rect 299716 236648 299722 236700
rect 307662 236648 307668 236700
rect 307720 236688 307726 236700
rect 321554 236688 321560 236700
rect 307720 236660 321560 236688
rect 307720 236648 307726 236660
rect 321554 236648 321560 236660
rect 321612 236648 321618 236700
rect 213362 236580 213368 236632
rect 213420 236620 213426 236632
rect 223666 236620 223672 236632
rect 213420 236592 223672 236620
rect 213420 236580 213426 236592
rect 223666 236580 223672 236592
rect 223724 236580 223730 236632
rect 241330 236580 241336 236632
rect 241388 236620 241394 236632
rect 242986 236620 242992 236632
rect 241388 236592 242992 236620
rect 241388 236580 241394 236592
rect 242986 236580 242992 236592
rect 243044 236580 243050 236632
rect 244826 236580 244832 236632
rect 244884 236620 244890 236632
rect 245286 236620 245292 236632
rect 244884 236592 245292 236620
rect 244884 236580 244890 236592
rect 245286 236580 245292 236592
rect 245344 236580 245350 236632
rect 247218 236580 247224 236632
rect 247276 236620 247282 236632
rect 247678 236620 247684 236632
rect 247276 236592 247684 236620
rect 247276 236580 247282 236592
rect 247678 236580 247684 236592
rect 247736 236580 247742 236632
rect 248230 236580 248236 236632
rect 248288 236620 248294 236632
rect 248966 236620 248972 236632
rect 248288 236592 248972 236620
rect 248288 236580 248294 236592
rect 248966 236580 248972 236592
rect 249024 236580 249030 236632
rect 266354 236580 266360 236632
rect 266412 236620 266418 236632
rect 330018 236620 330024 236632
rect 266412 236592 330024 236620
rect 266412 236580 266418 236592
rect 330018 236580 330024 236592
rect 330076 236580 330082 236632
rect 217594 236512 217600 236564
rect 217652 236552 217658 236564
rect 219986 236552 219992 236564
rect 217652 236524 219992 236552
rect 217652 236512 217658 236524
rect 219986 236512 219992 236524
rect 220044 236552 220050 236564
rect 254578 236552 254584 236564
rect 220044 236524 254584 236552
rect 220044 236512 220050 236524
rect 254578 236512 254584 236524
rect 254636 236512 254642 236564
rect 255774 236512 255780 236564
rect 255832 236552 255838 236564
rect 256418 236552 256424 236564
rect 255832 236524 256424 236552
rect 255832 236512 255838 236524
rect 256418 236512 256424 236524
rect 256476 236512 256482 236564
rect 259178 236512 259184 236564
rect 259236 236552 259242 236564
rect 276290 236552 276296 236564
rect 259236 236524 276296 236552
rect 259236 236512 259242 236524
rect 276290 236512 276296 236524
rect 276348 236512 276354 236564
rect 244826 236444 244832 236496
rect 244884 236484 244890 236496
rect 245470 236484 245476 236496
rect 244884 236456 245476 236484
rect 244884 236444 244890 236456
rect 245470 236444 245476 236456
rect 245528 236444 245534 236496
rect 253934 236444 253940 236496
rect 253992 236484 253998 236496
rect 255038 236484 255044 236496
rect 253992 236456 255044 236484
rect 253992 236444 253998 236456
rect 255038 236444 255044 236456
rect 255096 236444 255102 236496
rect 268378 236444 268384 236496
rect 268436 236484 268442 236496
rect 277394 236484 277400 236496
rect 268436 236456 277400 236484
rect 268436 236444 268442 236456
rect 277394 236444 277400 236456
rect 277452 236444 277458 236496
rect 244550 236376 244556 236428
rect 244608 236416 244614 236428
rect 249610 236416 249616 236428
rect 244608 236388 249616 236416
rect 244608 236376 244614 236388
rect 249610 236376 249616 236388
rect 249668 236416 249674 236428
rect 310146 236416 310152 236428
rect 249668 236388 310152 236416
rect 249668 236376 249674 236388
rect 310146 236376 310152 236388
rect 310204 236376 310210 236428
rect 252554 236308 252560 236360
rect 252612 236348 252618 236360
rect 261202 236348 261208 236360
rect 252612 236320 261208 236348
rect 252612 236308 252618 236320
rect 261202 236308 261208 236320
rect 261260 236308 261266 236360
rect 263502 236308 263508 236360
rect 263560 236348 263566 236360
rect 270770 236348 270776 236360
rect 263560 236320 270776 236348
rect 263560 236308 263566 236320
rect 270770 236308 270776 236320
rect 270828 236308 270834 236360
rect 233970 236104 233976 236156
rect 234028 236144 234034 236156
rect 244918 236144 244924 236156
rect 234028 236116 244924 236144
rect 234028 236104 234034 236116
rect 244918 236104 244924 236116
rect 244976 236144 244982 236156
rect 245654 236144 245660 236156
rect 244976 236116 245660 236144
rect 244976 236104 244982 236116
rect 245654 236104 245660 236116
rect 245712 236104 245718 236156
rect 237466 236036 237472 236088
rect 237524 236076 237530 236088
rect 238662 236076 238668 236088
rect 237524 236048 238668 236076
rect 237524 236036 237530 236048
rect 238662 236036 238668 236048
rect 238720 236036 238726 236088
rect 242066 236036 242072 236088
rect 242124 236076 242130 236088
rect 242124 236048 251174 236076
rect 242124 236036 242130 236048
rect 212350 235968 212356 236020
rect 212408 236008 212414 236020
rect 214834 236008 214840 236020
rect 212408 235980 214840 236008
rect 212408 235968 212414 235980
rect 214024 235952 214052 235980
rect 214834 235968 214840 235980
rect 214892 235968 214898 236020
rect 217502 235968 217508 236020
rect 217560 236008 217566 236020
rect 246298 236008 246304 236020
rect 217560 235980 246304 236008
rect 217560 235968 217566 235980
rect 246298 235968 246304 235980
rect 246356 236008 246362 236020
rect 246942 236008 246948 236020
rect 246356 235980 246948 236008
rect 246356 235968 246362 235980
rect 246942 235968 246948 235980
rect 247000 235968 247006 236020
rect 247126 235968 247132 236020
rect 247184 236008 247190 236020
rect 248414 236008 248420 236020
rect 247184 235980 248420 236008
rect 247184 235968 247190 235980
rect 248414 235968 248420 235980
rect 248472 235968 248478 236020
rect 214006 235900 214012 235952
rect 214064 235900 214070 235952
rect 224402 235900 224408 235952
rect 224460 235940 224466 235952
rect 224862 235940 224868 235952
rect 224460 235912 224868 235940
rect 224460 235900 224466 235912
rect 224862 235900 224868 235912
rect 224920 235900 224926 235952
rect 236914 235900 236920 235952
rect 236972 235940 236978 235952
rect 242066 235940 242072 235952
rect 236972 235912 242072 235940
rect 236972 235900 236978 235912
rect 242066 235900 242072 235912
rect 242124 235900 242130 235952
rect 207014 235832 207020 235884
rect 207072 235872 207078 235884
rect 208026 235872 208032 235884
rect 207072 235844 208032 235872
rect 207072 235832 207078 235844
rect 208026 235832 208032 235844
rect 208084 235872 208090 235884
rect 224218 235872 224224 235884
rect 208084 235844 224224 235872
rect 208084 235832 208090 235844
rect 224218 235832 224224 235844
rect 224276 235832 224282 235884
rect 242158 235832 242164 235884
rect 242216 235872 242222 235884
rect 243722 235872 243728 235884
rect 242216 235844 243728 235872
rect 242216 235832 242222 235844
rect 243722 235832 243728 235844
rect 243780 235832 243786 235884
rect 251146 235872 251174 236048
rect 256970 236036 256976 236088
rect 257028 236076 257034 236088
rect 267182 236076 267188 236088
rect 257028 236048 267188 236076
rect 257028 236036 257034 236048
rect 267182 236036 267188 236048
rect 267240 236036 267246 236088
rect 256050 235968 256056 236020
rect 256108 236008 256114 236020
rect 261478 236008 261484 236020
rect 256108 235980 261484 236008
rect 256108 235968 256114 235980
rect 261478 235968 261484 235980
rect 261536 235968 261542 236020
rect 265250 235968 265256 236020
rect 265308 236008 265314 236020
rect 265986 236008 265992 236020
rect 265308 235980 265992 236008
rect 265308 235968 265314 235980
rect 265986 235968 265992 235980
rect 266044 235968 266050 236020
rect 266170 235968 266176 236020
rect 266228 236008 266234 236020
rect 269022 236008 269028 236020
rect 266228 235980 269028 236008
rect 266228 235968 266234 235980
rect 269022 235968 269028 235980
rect 269080 236008 269086 236020
rect 272702 236008 272708 236020
rect 269080 235980 272708 236008
rect 269080 235968 269086 235980
rect 272702 235968 272708 235980
rect 272760 235968 272766 236020
rect 299658 235968 299664 236020
rect 299716 236008 299722 236020
rect 300394 236008 300400 236020
rect 299716 235980 300400 236008
rect 299716 235968 299722 235980
rect 300394 235968 300400 235980
rect 300452 235968 300458 236020
rect 288342 235900 288348 235952
rect 288400 235940 288406 235952
rect 329926 235940 329932 235952
rect 288400 235912 329932 235940
rect 288400 235900 288406 235912
rect 329926 235900 329932 235912
rect 329984 235900 329990 235952
rect 276934 235872 276940 235884
rect 251146 235844 276940 235872
rect 276934 235832 276940 235844
rect 276992 235832 276998 235884
rect 278774 235832 278780 235884
rect 278832 235872 278838 235884
rect 301958 235872 301964 235884
rect 278832 235844 301964 235872
rect 278832 235832 278838 235844
rect 301958 235832 301964 235844
rect 302016 235832 302022 235884
rect 242802 235764 242808 235816
rect 242860 235804 242866 235816
rect 244918 235804 244924 235816
rect 242860 235776 244924 235804
rect 242860 235764 242866 235776
rect 244918 235764 244924 235776
rect 244976 235764 244982 235816
rect 250346 235764 250352 235816
rect 250404 235804 250410 235816
rect 284846 235804 284852 235816
rect 250404 235776 284852 235804
rect 250404 235764 250410 235776
rect 284846 235764 284852 235776
rect 284904 235764 284910 235816
rect 210602 235696 210608 235748
rect 210660 235736 210666 235748
rect 245194 235736 245200 235748
rect 210660 235708 245200 235736
rect 210660 235696 210666 235708
rect 245194 235696 245200 235708
rect 245252 235696 245258 235748
rect 263318 235696 263324 235748
rect 263376 235736 263382 235748
rect 268930 235736 268936 235748
rect 263376 235708 268936 235736
rect 263376 235696 263382 235708
rect 268930 235696 268936 235708
rect 268988 235696 268994 235748
rect 269022 235696 269028 235748
rect 269080 235736 269086 235748
rect 277854 235736 277860 235748
rect 269080 235708 277860 235736
rect 269080 235696 269086 235708
rect 277854 235696 277860 235708
rect 277912 235696 277918 235748
rect 211614 235628 211620 235680
rect 211672 235668 211678 235680
rect 244550 235668 244556 235680
rect 211672 235640 244556 235668
rect 211672 235628 211678 235640
rect 244550 235628 244556 235640
rect 244608 235628 244614 235680
rect 266170 235628 266176 235680
rect 266228 235668 266234 235680
rect 267458 235668 267464 235680
rect 266228 235640 267464 235668
rect 266228 235628 266234 235640
rect 267458 235628 267464 235640
rect 267516 235628 267522 235680
rect 209222 235560 209228 235612
rect 209280 235600 209286 235612
rect 239398 235600 239404 235612
rect 209280 235572 239404 235600
rect 209280 235560 209286 235572
rect 239398 235560 239404 235572
rect 239456 235560 239462 235612
rect 252278 235560 252284 235612
rect 252336 235600 252342 235612
rect 252922 235600 252928 235612
rect 252336 235572 252928 235600
rect 252336 235560 252342 235572
rect 252922 235560 252928 235572
rect 252980 235560 252986 235612
rect 260190 235560 260196 235612
rect 260248 235600 260254 235612
rect 270218 235600 270224 235612
rect 260248 235572 270224 235600
rect 260248 235560 260254 235572
rect 270218 235560 270224 235572
rect 270276 235600 270282 235612
rect 281258 235600 281264 235612
rect 270276 235572 281264 235600
rect 270276 235560 270282 235572
rect 281258 235560 281264 235572
rect 281316 235560 281322 235612
rect 214834 235492 214840 235544
rect 214892 235532 214898 235544
rect 244734 235532 244740 235544
rect 214892 235504 244740 235532
rect 214892 235492 214898 235504
rect 244734 235492 244740 235504
rect 244792 235532 244798 235544
rect 285674 235532 285680 235544
rect 244792 235504 285680 235532
rect 244792 235492 244798 235504
rect 285674 235492 285680 235504
rect 285732 235492 285738 235544
rect 159634 235424 159640 235476
rect 159692 235464 159698 235476
rect 207014 235464 207020 235476
rect 159692 235436 207020 235464
rect 159692 235424 159698 235436
rect 207014 235424 207020 235436
rect 207072 235424 207078 235476
rect 210694 235424 210700 235476
rect 210752 235464 210758 235476
rect 256418 235464 256424 235476
rect 210752 235436 256424 235464
rect 210752 235424 210758 235436
rect 256418 235424 256424 235436
rect 256476 235424 256482 235476
rect 264698 235424 264704 235476
rect 264756 235464 264762 235476
rect 282454 235464 282460 235476
rect 264756 235436 282460 235464
rect 264756 235424 264762 235436
rect 282454 235424 282460 235436
rect 282512 235464 282518 235476
rect 331490 235464 331496 235476
rect 282512 235436 331496 235464
rect 282512 235424 282518 235436
rect 331490 235424 331496 235436
rect 331548 235424 331554 235476
rect 161014 235356 161020 235408
rect 161072 235396 161078 235408
rect 216674 235396 216680 235408
rect 161072 235368 216680 235396
rect 161072 235356 161078 235368
rect 216674 235356 216680 235368
rect 216732 235356 216738 235408
rect 225966 235396 225972 235408
rect 220096 235368 225972 235396
rect 155770 235288 155776 235340
rect 155828 235328 155834 235340
rect 216490 235328 216496 235340
rect 155828 235300 216496 235328
rect 155828 235288 155834 235300
rect 216490 235288 216496 235300
rect 216548 235328 216554 235340
rect 220096 235328 220124 235368
rect 225966 235356 225972 235368
rect 226024 235356 226030 235408
rect 229738 235356 229744 235408
rect 229796 235396 229802 235408
rect 230382 235396 230388 235408
rect 229796 235368 230388 235396
rect 229796 235356 229802 235368
rect 230382 235356 230388 235368
rect 230440 235356 230446 235408
rect 245470 235356 245476 235408
rect 245528 235396 245534 235408
rect 246482 235396 246488 235408
rect 245528 235368 246488 235396
rect 245528 235356 245534 235368
rect 246482 235356 246488 235368
rect 246540 235356 246546 235408
rect 260558 235356 260564 235408
rect 260616 235396 260622 235408
rect 273898 235396 273904 235408
rect 260616 235368 273904 235396
rect 260616 235356 260622 235368
rect 273898 235356 273904 235368
rect 273956 235396 273962 235408
rect 328638 235396 328644 235408
rect 273956 235368 328644 235396
rect 273956 235356 273962 235368
rect 328638 235356 328644 235368
rect 328696 235356 328702 235408
rect 216548 235300 220124 235328
rect 216548 235288 216554 235300
rect 220170 235288 220176 235340
rect 220228 235328 220234 235340
rect 237098 235328 237104 235340
rect 220228 235300 237104 235328
rect 220228 235288 220234 235300
rect 237098 235288 237104 235300
rect 237156 235288 237162 235340
rect 243446 235288 243452 235340
rect 243504 235328 243510 235340
rect 243906 235328 243912 235340
rect 243504 235300 243912 235328
rect 243504 235288 243510 235300
rect 243906 235288 243912 235300
rect 243964 235288 243970 235340
rect 261662 235288 261668 235340
rect 261720 235328 261726 235340
rect 267918 235328 267924 235340
rect 261720 235300 267924 235328
rect 261720 235288 261726 235300
rect 267918 235288 267924 235300
rect 267976 235288 267982 235340
rect 268930 235288 268936 235340
rect 268988 235328 268994 235340
rect 271230 235328 271236 235340
rect 268988 235300 271236 235328
rect 268988 235288 268994 235300
rect 271230 235288 271236 235300
rect 271288 235328 271294 235340
rect 329098 235328 329104 235340
rect 271288 235300 329104 235328
rect 271288 235288 271294 235300
rect 329098 235288 329104 235300
rect 329156 235288 329162 235340
rect 158438 235220 158444 235272
rect 158496 235260 158502 235272
rect 233142 235260 233148 235272
rect 158496 235232 233148 235260
rect 158496 235220 158502 235232
rect 233142 235220 233148 235232
rect 233200 235220 233206 235272
rect 234706 235220 234712 235272
rect 234764 235260 234770 235272
rect 235718 235260 235724 235272
rect 234764 235232 235724 235260
rect 234764 235220 234770 235232
rect 235718 235220 235724 235232
rect 235776 235220 235782 235272
rect 258350 235260 258356 235272
rect 244246 235232 258356 235260
rect 207014 235152 207020 235204
rect 207072 235192 207078 235204
rect 207842 235192 207848 235204
rect 207072 235164 207848 235192
rect 207072 235152 207078 235164
rect 207842 235152 207848 235164
rect 207900 235192 207906 235204
rect 227714 235192 227720 235204
rect 207900 235164 227720 235192
rect 207900 235152 207906 235164
rect 227714 235152 227720 235164
rect 227772 235152 227778 235204
rect 236638 235152 236644 235204
rect 236696 235192 236702 235204
rect 244246 235192 244274 235232
rect 258350 235220 258356 235232
rect 258408 235260 258414 235272
rect 259454 235260 259460 235272
rect 258408 235232 259460 235260
rect 258408 235220 258414 235232
rect 259454 235220 259460 235232
rect 259512 235220 259518 235272
rect 260926 235220 260932 235272
rect 260984 235260 260990 235272
rect 269114 235260 269120 235272
rect 260984 235232 269120 235260
rect 260984 235220 260990 235232
rect 269114 235220 269120 235232
rect 269172 235260 269178 235272
rect 331582 235260 331588 235272
rect 269172 235232 331588 235260
rect 269172 235220 269178 235232
rect 331582 235220 331588 235232
rect 331640 235220 331646 235272
rect 236696 235164 244274 235192
rect 236696 235152 236702 235164
rect 254026 235152 254032 235204
rect 254084 235192 254090 235204
rect 254670 235192 254676 235204
rect 254084 235164 254676 235192
rect 254084 235152 254090 235164
rect 254670 235152 254676 235164
rect 254728 235152 254734 235204
rect 257614 235152 257620 235204
rect 257672 235192 257678 235204
rect 266446 235192 266452 235204
rect 257672 235164 266452 235192
rect 257672 235152 257678 235164
rect 266446 235152 266452 235164
rect 266504 235152 266510 235204
rect 239398 235084 239404 235136
rect 239456 235124 239462 235136
rect 250806 235124 250812 235136
rect 239456 235096 250812 235124
rect 239456 235084 239462 235096
rect 250806 235084 250812 235096
rect 250864 235124 250870 235136
rect 263870 235124 263876 235136
rect 250864 235096 263876 235124
rect 250864 235084 250870 235096
rect 263870 235084 263876 235096
rect 263928 235084 263934 235136
rect 266354 235084 266360 235136
rect 266412 235124 266418 235136
rect 266998 235124 267004 235136
rect 266412 235096 267004 235124
rect 266412 235084 266418 235096
rect 266998 235084 267004 235096
rect 267056 235084 267062 235136
rect 222562 235016 222568 235068
rect 222620 235056 222626 235068
rect 226150 235056 226156 235068
rect 222620 235028 226156 235056
rect 222620 235016 222626 235028
rect 226150 235016 226156 235028
rect 226208 235016 226214 235068
rect 256878 235016 256884 235068
rect 256936 235056 256942 235068
rect 257246 235056 257252 235068
rect 256936 235028 257252 235056
rect 256936 235016 256942 235028
rect 257246 235016 257252 235028
rect 257304 235016 257310 235068
rect 259454 235016 259460 235068
rect 259512 235056 259518 235068
rect 270126 235056 270132 235068
rect 259512 235028 270132 235056
rect 259512 235016 259518 235028
rect 270126 235016 270132 235028
rect 270184 235016 270190 235068
rect 244642 234948 244648 235000
rect 244700 234988 244706 235000
rect 245194 234988 245200 235000
rect 244700 234960 245200 234988
rect 244700 234948 244706 234960
rect 245194 234948 245200 234960
rect 245252 234948 245258 235000
rect 245654 234948 245660 235000
rect 245712 234988 245718 235000
rect 289078 234988 289084 235000
rect 245712 234960 289084 234988
rect 245712 234948 245718 234960
rect 289078 234948 289084 234960
rect 289136 234948 289142 235000
rect 237190 234880 237196 234932
rect 237248 234920 237254 234932
rect 240410 234920 240416 234932
rect 237248 234892 240416 234920
rect 237248 234880 237254 234892
rect 240410 234880 240416 234892
rect 240468 234880 240474 234932
rect 240870 234880 240876 234932
rect 240928 234920 240934 234932
rect 241054 234920 241060 234932
rect 240928 234892 241060 234920
rect 240928 234880 240934 234892
rect 241054 234880 241060 234892
rect 241112 234880 241118 234932
rect 262306 234880 262312 234932
rect 262364 234920 262370 234932
rect 269022 234920 269028 234932
rect 262364 234892 269028 234920
rect 262364 234880 262370 234892
rect 269022 234880 269028 234892
rect 269080 234880 269086 234932
rect 251910 234812 251916 234864
rect 251968 234852 251974 234864
rect 265802 234852 265808 234864
rect 251968 234824 265808 234852
rect 251968 234812 251974 234824
rect 265802 234812 265808 234824
rect 265860 234812 265866 234864
rect 232866 234744 232872 234796
rect 232924 234784 232930 234796
rect 238294 234784 238300 234796
rect 232924 234756 238300 234784
rect 232924 234744 232930 234756
rect 238294 234744 238300 234756
rect 238352 234744 238358 234796
rect 263042 234744 263048 234796
rect 263100 234784 263106 234796
rect 270126 234784 270132 234796
rect 263100 234756 270132 234784
rect 263100 234744 263106 234756
rect 270126 234744 270132 234756
rect 270184 234744 270190 234796
rect 245470 234716 245476 234728
rect 234586 234688 245476 234716
rect 215938 234608 215944 234660
rect 215996 234648 216002 234660
rect 234586 234648 234614 234688
rect 245470 234676 245476 234688
rect 245528 234676 245534 234728
rect 258350 234676 258356 234728
rect 258408 234716 258414 234728
rect 259270 234716 259276 234728
rect 258408 234688 259276 234716
rect 258408 234676 258414 234688
rect 259270 234676 259276 234688
rect 259328 234676 259334 234728
rect 260834 234676 260840 234728
rect 260892 234716 260898 234728
rect 261570 234716 261576 234728
rect 260892 234688 261576 234716
rect 260892 234676 260898 234688
rect 261570 234676 261576 234688
rect 261628 234676 261634 234728
rect 263502 234676 263508 234728
rect 263560 234716 263566 234728
rect 263778 234716 263784 234728
rect 263560 234688 263784 234716
rect 263560 234676 263566 234688
rect 263778 234676 263784 234688
rect 263836 234676 263842 234728
rect 265158 234676 265164 234728
rect 265216 234716 265222 234728
rect 265710 234716 265716 234728
rect 265216 234688 265716 234716
rect 265216 234676 265222 234688
rect 265710 234676 265716 234688
rect 265768 234676 265774 234728
rect 284294 234676 284300 234728
rect 284352 234716 284358 234728
rect 284846 234716 284852 234728
rect 284352 234688 284852 234716
rect 284352 234676 284358 234688
rect 284846 234676 284852 234688
rect 284904 234676 284910 234728
rect 215996 234620 234614 234648
rect 215996 234608 216002 234620
rect 247310 234608 247316 234660
rect 247368 234648 247374 234660
rect 291838 234648 291844 234660
rect 247368 234620 291844 234648
rect 247368 234608 247374 234620
rect 291838 234608 291844 234620
rect 291896 234608 291902 234660
rect 212534 234540 212540 234592
rect 212592 234580 212598 234592
rect 243354 234580 243360 234592
rect 212592 234552 243360 234580
rect 212592 234540 212598 234552
rect 243354 234540 243360 234552
rect 243412 234540 243418 234592
rect 243538 234540 243544 234592
rect 243596 234580 243602 234592
rect 303062 234580 303068 234592
rect 243596 234552 303068 234580
rect 243596 234540 243602 234552
rect 303062 234540 303068 234552
rect 303120 234540 303126 234592
rect 211890 234472 211896 234524
rect 211948 234512 211954 234524
rect 246666 234512 246672 234524
rect 211948 234484 246672 234512
rect 211948 234472 211954 234484
rect 246666 234472 246672 234484
rect 246724 234472 246730 234524
rect 247034 234472 247040 234524
rect 247092 234512 247098 234524
rect 305638 234512 305644 234524
rect 247092 234484 305644 234512
rect 247092 234472 247098 234484
rect 305638 234472 305644 234484
rect 305696 234472 305702 234524
rect 237650 234404 237656 234456
rect 237708 234444 237714 234456
rect 286870 234444 286876 234456
rect 237708 234416 286876 234444
rect 237708 234404 237714 234416
rect 286870 234404 286876 234416
rect 286928 234404 286934 234456
rect 223758 234336 223764 234388
rect 223816 234376 223822 234388
rect 226058 234376 226064 234388
rect 223816 234348 226064 234376
rect 223816 234336 223822 234348
rect 226058 234336 226064 234348
rect 226116 234336 226122 234388
rect 228174 234336 228180 234388
rect 228232 234376 228238 234388
rect 228450 234376 228456 234388
rect 228232 234348 228456 234376
rect 228232 234336 228238 234348
rect 228450 234336 228456 234348
rect 228508 234336 228514 234388
rect 237006 234336 237012 234388
rect 237064 234376 237070 234388
rect 279878 234376 279884 234388
rect 237064 234348 279884 234376
rect 237064 234336 237070 234348
rect 279878 234336 279884 234348
rect 279936 234336 279942 234388
rect 285674 234336 285680 234388
rect 285732 234376 285738 234388
rect 304626 234376 304632 234388
rect 285732 234348 304632 234376
rect 285732 234336 285738 234348
rect 304626 234336 304632 234348
rect 304684 234336 304690 234388
rect 249794 234268 249800 234320
rect 249852 234308 249858 234320
rect 293218 234308 293224 234320
rect 249852 234280 293224 234308
rect 249852 234268 249858 234280
rect 293218 234268 293224 234280
rect 293276 234268 293282 234320
rect 237558 234200 237564 234252
rect 237616 234240 237622 234252
rect 238294 234240 238300 234252
rect 237616 234212 238300 234240
rect 237616 234200 237622 234212
rect 238294 234200 238300 234212
rect 238352 234200 238358 234252
rect 239582 234200 239588 234252
rect 239640 234240 239646 234252
rect 282730 234240 282736 234252
rect 239640 234212 282736 234240
rect 239640 234200 239646 234212
rect 282730 234200 282736 234212
rect 282788 234200 282794 234252
rect 210786 234132 210792 234184
rect 210844 234172 210850 234184
rect 212534 234172 212540 234184
rect 210844 234144 212540 234172
rect 210844 234132 210850 234144
rect 212534 234132 212540 234144
rect 212592 234132 212598 234184
rect 219986 234132 219992 234184
rect 220044 234172 220050 234184
rect 220044 234144 223574 234172
rect 220044 234132 220050 234144
rect 153102 234064 153108 234116
rect 153160 234104 153166 234116
rect 211982 234104 211988 234116
rect 153160 234076 211988 234104
rect 153160 234064 153166 234076
rect 211982 234064 211988 234076
rect 212040 234064 212046 234116
rect 223546 234104 223574 234144
rect 237098 234132 237104 234184
rect 237156 234172 237162 234184
rect 240778 234172 240784 234184
rect 237156 234144 240784 234172
rect 237156 234132 237162 234144
rect 240778 234132 240784 234144
rect 240836 234172 240842 234184
rect 281902 234172 281908 234184
rect 240836 234144 281908 234172
rect 240836 234132 240842 234144
rect 281902 234132 281908 234144
rect 281960 234132 281966 234184
rect 238202 234104 238208 234116
rect 223546 234076 238208 234104
rect 238202 234064 238208 234076
rect 238260 234104 238266 234116
rect 277762 234104 277768 234116
rect 238260 234076 277768 234104
rect 238260 234064 238266 234076
rect 277762 234064 277768 234076
rect 277820 234064 277826 234116
rect 161106 233996 161112 234048
rect 161164 234036 161170 234048
rect 234890 234036 234896 234048
rect 161164 234008 234896 234036
rect 161164 233996 161170 234008
rect 234890 233996 234896 234008
rect 234948 233996 234954 234048
rect 236270 233996 236276 234048
rect 236328 234036 236334 234048
rect 276842 234036 276848 234048
rect 236328 234008 276848 234036
rect 236328 233996 236334 234008
rect 276842 233996 276848 234008
rect 276900 233996 276906 234048
rect 156966 233928 156972 233980
rect 157024 233968 157030 233980
rect 224862 233968 224868 233980
rect 157024 233940 224868 233968
rect 157024 233928 157030 233940
rect 224862 233928 224868 233940
rect 224920 233928 224926 233980
rect 240594 233928 240600 233980
rect 240652 233968 240658 233980
rect 279694 233968 279700 233980
rect 240652 233940 279700 233968
rect 240652 233928 240658 233940
rect 279694 233928 279700 233940
rect 279752 233928 279758 233980
rect 151630 233860 151636 233912
rect 151688 233900 151694 233912
rect 231210 233900 231216 233912
rect 151688 233872 231216 233900
rect 151688 233860 151694 233872
rect 231210 233860 231216 233872
rect 231268 233860 231274 233912
rect 273530 233900 273536 233912
rect 241532 233872 273536 233900
rect 216122 233588 216128 233640
rect 216180 233628 216186 233640
rect 217778 233628 217784 233640
rect 216180 233600 217784 233628
rect 216180 233588 216186 233600
rect 217778 233588 217784 233600
rect 217836 233588 217842 233640
rect 241422 233588 241428 233640
rect 241480 233628 241486 233640
rect 241532 233628 241560 233872
rect 273530 233860 273536 233872
rect 273588 233860 273594 233912
rect 243538 233792 243544 233844
rect 243596 233832 243602 233844
rect 244182 233832 244188 233844
rect 243596 233804 244188 233832
rect 243596 233792 243602 233804
rect 244182 233792 244188 233804
rect 244240 233792 244246 233844
rect 246114 233792 246120 233844
rect 246172 233832 246178 233844
rect 271782 233832 271788 233844
rect 246172 233804 271788 233832
rect 246172 233792 246178 233804
rect 271782 233792 271788 233804
rect 271840 233792 271846 233844
rect 272518 233792 272524 233844
rect 272576 233832 272582 233844
rect 272886 233832 272892 233844
rect 272576 233804 272892 233832
rect 272576 233792 272582 233804
rect 272886 233792 272892 233804
rect 272944 233792 272950 233844
rect 244918 233724 244924 233776
rect 244976 233764 244982 233776
rect 274358 233764 274364 233776
rect 244976 233736 274364 233764
rect 244976 233724 244982 233736
rect 274358 233724 274364 233736
rect 274416 233724 274422 233776
rect 272518 233696 272524 233708
rect 241480 233600 241560 233628
rect 253906 233668 272524 233696
rect 241480 233588 241486 233600
rect 247954 233520 247960 233572
rect 248012 233560 248018 233572
rect 253906 233560 253934 233668
rect 272518 233656 272524 233668
rect 272576 233656 272582 233708
rect 256694 233588 256700 233640
rect 256752 233628 256758 233640
rect 257430 233628 257436 233640
rect 256752 233600 257436 233628
rect 256752 233588 256758 233600
rect 257430 233588 257436 233600
rect 257488 233588 257494 233640
rect 260006 233588 260012 233640
rect 260064 233628 260070 233640
rect 260466 233628 260472 233640
rect 260064 233600 260472 233628
rect 260064 233588 260070 233600
rect 260466 233588 260472 233600
rect 260524 233588 260530 233640
rect 271782 233588 271788 233640
rect 271840 233628 271846 233640
rect 274818 233628 274824 233640
rect 271840 233600 274824 233628
rect 271840 233588 271846 233600
rect 274818 233588 274824 233600
rect 274876 233588 274882 233640
rect 248012 233532 253934 233560
rect 248012 233520 248018 233532
rect 263686 233520 263692 233572
rect 263744 233560 263750 233572
rect 264514 233560 264520 233572
rect 263744 233532 264520 233560
rect 263744 233520 263750 233532
rect 264514 233520 264520 233532
rect 264572 233520 264578 233572
rect 219526 233316 219532 233368
rect 219584 233356 219590 233368
rect 223850 233356 223856 233368
rect 219584 233328 223856 233356
rect 219584 233316 219590 233328
rect 223850 233316 223856 233328
rect 223908 233316 223914 233368
rect 248322 233316 248328 233368
rect 248380 233356 248386 233368
rect 249794 233356 249800 233368
rect 248380 233328 249800 233356
rect 248380 233316 248386 233328
rect 249794 233316 249800 233328
rect 249852 233316 249858 233368
rect 217410 233248 217416 233300
rect 217468 233288 217474 233300
rect 231854 233288 231860 233300
rect 217468 233260 231860 233288
rect 217468 233248 217474 233260
rect 231854 233248 231860 233260
rect 231912 233248 231918 233300
rect 258258 233248 258264 233300
rect 258316 233288 258322 233300
rect 259362 233288 259368 233300
rect 258316 233260 259368 233288
rect 258316 233248 258322 233260
rect 259362 233248 259368 233260
rect 259420 233248 259426 233300
rect 278038 233248 278044 233300
rect 278096 233288 278102 233300
rect 278096 233260 278452 233288
rect 278096 233248 278102 233260
rect 212442 233180 212448 233232
rect 212500 233220 212506 233232
rect 212500 233192 213914 233220
rect 212500 233180 212506 233192
rect 213886 233152 213914 233192
rect 219802 233180 219808 233232
rect 219860 233220 219866 233232
rect 226426 233220 226432 233232
rect 219860 233192 226432 233220
rect 219860 233180 219866 233192
rect 226426 233180 226432 233192
rect 226484 233220 226490 233232
rect 227162 233220 227168 233232
rect 226484 233192 227168 233220
rect 226484 233180 226490 233192
rect 227162 233180 227168 233192
rect 227220 233180 227226 233232
rect 276198 233180 276204 233232
rect 276256 233220 276262 233232
rect 278314 233220 278320 233232
rect 276256 233192 278320 233220
rect 276256 233180 276262 233192
rect 278314 233180 278320 233192
rect 278372 233180 278378 233232
rect 278424 233220 278452 233260
rect 579614 233220 579620 233232
rect 278424 233192 579620 233220
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 222562 233152 222568 233164
rect 213886 233124 222568 233152
rect 222562 233112 222568 233124
rect 222620 233112 222626 233164
rect 249426 233112 249432 233164
rect 249484 233152 249490 233164
rect 335446 233152 335452 233164
rect 249484 233124 335452 233152
rect 249484 233112 249490 233124
rect 335446 233112 335452 233124
rect 335504 233112 335510 233164
rect 219158 233044 219164 233096
rect 219216 233084 219222 233096
rect 223758 233084 223764 233096
rect 219216 233056 223764 233084
rect 219216 233044 219222 233056
rect 223758 233044 223764 233056
rect 223816 233044 223822 233096
rect 245194 233044 245200 233096
rect 245252 233084 245258 233096
rect 300302 233084 300308 233096
rect 245252 233056 300308 233084
rect 245252 233044 245258 233056
rect 300302 233044 300308 233056
rect 300360 233044 300366 233096
rect 219710 233016 219716 233028
rect 219406 232988 219716 233016
rect 194410 232840 194416 232892
rect 194468 232880 194474 232892
rect 219406 232880 219434 232988
rect 219710 232976 219716 232988
rect 219768 233016 219774 233028
rect 252554 233016 252560 233028
rect 219768 232988 252560 233016
rect 219768 232976 219774 232988
rect 252554 232976 252560 232988
rect 252612 232976 252618 233028
rect 253198 232976 253204 233028
rect 253256 233016 253262 233028
rect 304534 233016 304540 233028
rect 253256 232988 304540 233016
rect 253256 232976 253262 232988
rect 304534 232976 304540 232988
rect 304592 232976 304598 233028
rect 248874 232908 248880 232960
rect 248932 232948 248938 232960
rect 296254 232948 296260 232960
rect 248932 232920 296260 232948
rect 248932 232908 248938 232920
rect 296254 232908 296260 232920
rect 296312 232908 296318 232960
rect 194468 232852 219434 232880
rect 194468 232840 194474 232852
rect 252278 232840 252284 232892
rect 252336 232880 252342 232892
rect 297726 232880 297732 232892
rect 252336 232852 297732 232880
rect 252336 232840 252342 232852
rect 297726 232840 297732 232852
rect 297784 232840 297790 232892
rect 159542 232772 159548 232824
rect 159600 232812 159606 232824
rect 209406 232812 209412 232824
rect 159600 232784 209412 232812
rect 159600 232772 159606 232784
rect 209406 232772 209412 232784
rect 209464 232772 209470 232824
rect 235534 232772 235540 232824
rect 235592 232812 235598 232824
rect 274266 232812 274272 232824
rect 235592 232784 274272 232812
rect 235592 232772 235598 232784
rect 274266 232772 274272 232784
rect 274324 232772 274330 232824
rect 277854 232772 277860 232824
rect 277912 232812 277918 232824
rect 281074 232812 281080 232824
rect 277912 232784 281080 232812
rect 277912 232772 277918 232784
rect 281074 232772 281080 232784
rect 281132 232772 281138 232824
rect 156874 232704 156880 232756
rect 156932 232744 156938 232756
rect 207014 232744 207020 232756
rect 156932 232716 207020 232744
rect 156932 232704 156938 232716
rect 207014 232704 207020 232716
rect 207072 232704 207078 232756
rect 232498 232704 232504 232756
rect 232556 232744 232562 232756
rect 240962 232744 240968 232756
rect 232556 232716 240968 232744
rect 232556 232704 232562 232716
rect 240962 232704 240968 232716
rect 241020 232744 241026 232756
rect 275278 232744 275284 232756
rect 241020 232716 275284 232744
rect 241020 232704 241026 232716
rect 275278 232704 275284 232716
rect 275336 232704 275342 232756
rect 161474 232636 161480 232688
rect 161532 232676 161538 232688
rect 191650 232676 191656 232688
rect 161532 232648 191656 232676
rect 161532 232636 161538 232648
rect 191650 232636 191656 232648
rect 191708 232636 191714 232688
rect 195882 232636 195888 232688
rect 195940 232676 195946 232688
rect 256050 232676 256056 232688
rect 195940 232648 256056 232676
rect 195940 232636 195946 232648
rect 256050 232636 256056 232648
rect 256108 232636 256114 232688
rect 261202 232636 261208 232688
rect 261260 232676 261266 232688
rect 287146 232676 287152 232688
rect 261260 232648 287152 232676
rect 261260 232636 261266 232648
rect 287146 232636 287152 232648
rect 287204 232676 287210 232688
rect 287606 232676 287612 232688
rect 287204 232648 287612 232676
rect 287204 232636 287210 232648
rect 287606 232636 287612 232648
rect 287664 232636 287670 232688
rect 155678 232568 155684 232620
rect 155736 232608 155742 232620
rect 231670 232608 231676 232620
rect 155736 232580 231676 232608
rect 155736 232568 155742 232580
rect 231670 232568 231676 232580
rect 231728 232568 231734 232620
rect 240318 232568 240324 232620
rect 240376 232608 240382 232620
rect 240962 232608 240968 232620
rect 240376 232580 240968 232608
rect 240376 232568 240382 232580
rect 240962 232568 240968 232580
rect 241020 232568 241026 232620
rect 241698 232568 241704 232620
rect 241756 232608 241762 232620
rect 242710 232608 242716 232620
rect 241756 232580 242716 232608
rect 241756 232568 241762 232580
rect 242710 232568 242716 232580
rect 242768 232568 242774 232620
rect 249150 232568 249156 232620
rect 249208 232608 249214 232620
rect 278406 232608 278412 232620
rect 249208 232580 278412 232608
rect 249208 232568 249214 232580
rect 278406 232568 278412 232580
rect 278464 232608 278470 232620
rect 279234 232608 279240 232620
rect 278464 232580 279240 232608
rect 278464 232568 278470 232580
rect 279234 232568 279240 232580
rect 279292 232568 279298 232620
rect 157058 232500 157064 232552
rect 157116 232540 157122 232552
rect 234614 232540 234620 232552
rect 157116 232512 234620 232540
rect 157116 232500 157122 232512
rect 234614 232500 234620 232512
rect 234672 232500 234678 232552
rect 253566 232500 253572 232552
rect 253624 232540 253630 232552
rect 284018 232540 284024 232552
rect 253624 232512 284024 232540
rect 253624 232500 253630 232512
rect 284018 232500 284024 232512
rect 284076 232540 284082 232552
rect 328546 232540 328552 232552
rect 284076 232512 328552 232540
rect 284076 232500 284082 232512
rect 328546 232500 328552 232512
rect 328604 232500 328610 232552
rect 225690 232432 225696 232484
rect 225748 232472 225754 232484
rect 226794 232472 226800 232484
rect 225748 232444 226800 232472
rect 225748 232432 225754 232444
rect 226794 232432 226800 232444
rect 226852 232432 226858 232484
rect 233694 232432 233700 232484
rect 233752 232472 233758 232484
rect 234246 232472 234252 232484
rect 233752 232444 234252 232472
rect 233752 232432 233758 232444
rect 234246 232432 234252 232444
rect 234304 232432 234310 232484
rect 247494 232432 247500 232484
rect 247552 232472 247558 232484
rect 271138 232472 271144 232484
rect 247552 232444 271144 232472
rect 247552 232432 247558 232444
rect 271138 232432 271144 232444
rect 271196 232432 271202 232484
rect 280246 232432 280252 232484
rect 280304 232472 280310 232484
rect 282546 232472 282552 232484
rect 280304 232444 282552 232472
rect 280304 232432 280310 232444
rect 282546 232432 282552 232444
rect 282604 232432 282610 232484
rect 243170 232364 243176 232416
rect 243228 232404 243234 232416
rect 260190 232404 260196 232416
rect 243228 232376 260196 232404
rect 243228 232364 243234 232376
rect 260190 232364 260196 232376
rect 260248 232404 260254 232416
rect 269298 232404 269304 232416
rect 260248 232376 269304 232404
rect 260248 232364 260254 232376
rect 269298 232364 269304 232376
rect 269356 232364 269362 232416
rect 236730 232296 236736 232348
rect 236788 232336 236794 232348
rect 239674 232336 239680 232348
rect 236788 232308 239680 232336
rect 236788 232296 236794 232308
rect 239674 232296 239680 232308
rect 239732 232336 239738 232348
rect 280614 232336 280620 232348
rect 239732 232308 280620 232336
rect 239732 232296 239738 232308
rect 280614 232296 280620 232308
rect 280672 232296 280678 232348
rect 242066 232160 242072 232212
rect 242124 232200 242130 232212
rect 242434 232200 242440 232212
rect 242124 232172 242440 232200
rect 242124 232160 242130 232172
rect 242434 232160 242440 232172
rect 242492 232160 242498 232212
rect 229462 231888 229468 231940
rect 229520 231928 229526 231940
rect 230382 231928 230388 231940
rect 229520 231900 230388 231928
rect 229520 231888 229526 231900
rect 230382 231888 230388 231900
rect 230440 231888 230446 231940
rect 227990 231820 227996 231872
rect 228048 231860 228054 231872
rect 230750 231860 230756 231872
rect 228048 231832 230756 231860
rect 228048 231820 228054 231832
rect 230750 231820 230756 231832
rect 230808 231820 230814 231872
rect 254762 231820 254768 231872
rect 254820 231860 254826 231872
rect 264514 231860 264520 231872
rect 254820 231832 264520 231860
rect 254820 231820 254826 231832
rect 264514 231820 264520 231832
rect 264572 231820 264578 231872
rect 209498 231752 209504 231804
rect 209556 231792 209562 231804
rect 229646 231792 229652 231804
rect 209556 231764 229652 231792
rect 209556 231752 209562 231764
rect 229646 231752 229652 231764
rect 229704 231752 229710 231804
rect 242618 231752 242624 231804
rect 242676 231792 242682 231804
rect 243630 231792 243636 231804
rect 242676 231764 243636 231792
rect 242676 231752 242682 231764
rect 243630 231752 243636 231764
rect 243688 231752 243694 231804
rect 261570 231752 261576 231804
rect 261628 231792 261634 231804
rect 262398 231792 262404 231804
rect 261628 231764 262404 231792
rect 261628 231752 261634 231764
rect 262398 231752 262404 231764
rect 262456 231752 262462 231804
rect 262490 231752 262496 231804
rect 262548 231792 262554 231804
rect 269666 231792 269672 231804
rect 262548 231764 269672 231792
rect 262548 231752 262554 231764
rect 269666 231752 269672 231764
rect 269724 231752 269730 231804
rect 284386 231752 284392 231804
rect 284444 231792 284450 231804
rect 285122 231792 285128 231804
rect 284444 231764 285128 231792
rect 284444 231752 284450 231764
rect 285122 231752 285128 231764
rect 285180 231752 285186 231804
rect 291286 231752 291292 231804
rect 291344 231792 291350 231804
rect 291930 231792 291936 231804
rect 291344 231764 291936 231792
rect 291344 231752 291350 231764
rect 291930 231752 291936 231764
rect 291988 231752 291994 231804
rect 230750 231684 230756 231736
rect 230808 231724 230814 231736
rect 230934 231724 230940 231736
rect 230808 231696 230940 231724
rect 230808 231684 230814 231696
rect 230934 231684 230940 231696
rect 230992 231684 230998 231736
rect 240962 231684 240968 231736
rect 241020 231724 241026 231736
rect 300486 231724 300492 231736
rect 241020 231696 300492 231724
rect 241020 231684 241026 231696
rect 300486 231684 300492 231696
rect 300544 231684 300550 231736
rect 246758 231616 246764 231668
rect 246816 231656 246822 231668
rect 248782 231656 248788 231668
rect 246816 231628 248788 231656
rect 246816 231616 246822 231628
rect 248782 231616 248788 231628
rect 248840 231616 248846 231668
rect 256786 231616 256792 231668
rect 256844 231656 256850 231668
rect 316862 231656 316868 231668
rect 256844 231628 316868 231656
rect 256844 231616 256850 231628
rect 316862 231616 316868 231628
rect 316920 231616 316926 231668
rect 250070 231548 250076 231600
rect 250128 231588 250134 231600
rect 250806 231588 250812 231600
rect 250128 231560 250812 231588
rect 250128 231548 250134 231560
rect 250806 231548 250812 231560
rect 250864 231588 250870 231600
rect 294874 231588 294880 231600
rect 250864 231560 294880 231588
rect 250864 231548 250870 231560
rect 294874 231548 294880 231560
rect 294932 231548 294938 231600
rect 234522 231480 234528 231532
rect 234580 231520 234586 231532
rect 261754 231520 261760 231532
rect 234580 231492 261760 231520
rect 234580 231480 234586 231492
rect 261754 231480 261760 231492
rect 261812 231480 261818 231532
rect 262398 231480 262404 231532
rect 262456 231520 262462 231532
rect 305178 231520 305184 231532
rect 262456 231492 305184 231520
rect 262456 231480 262462 231492
rect 305178 231480 305184 231492
rect 305236 231480 305242 231532
rect 252370 231412 252376 231464
rect 252428 231452 252434 231464
rect 284386 231452 284392 231464
rect 252428 231424 284392 231452
rect 252428 231412 252434 231424
rect 284386 231412 284392 231424
rect 284444 231412 284450 231464
rect 291194 231412 291200 231464
rect 291252 231452 291258 231464
rect 292298 231452 292304 231464
rect 291252 231424 292304 231452
rect 291252 231412 291258 231424
rect 292298 231412 292304 231424
rect 292356 231412 292362 231464
rect 234062 231344 234068 231396
rect 234120 231384 234126 231396
rect 234430 231384 234436 231396
rect 234120 231356 234436 231384
rect 234120 231344 234126 231356
rect 234430 231344 234436 231356
rect 234488 231344 234494 231396
rect 246850 231344 246856 231396
rect 246908 231384 246914 231396
rect 277578 231384 277584 231396
rect 246908 231356 277584 231384
rect 246908 231344 246914 231356
rect 277578 231344 277584 231356
rect 277636 231384 277642 231396
rect 277854 231384 277860 231396
rect 277636 231356 277860 231384
rect 277636 231344 277642 231356
rect 277854 231344 277860 231356
rect 277912 231344 277918 231396
rect 199838 231276 199844 231328
rect 199896 231316 199902 231328
rect 259086 231316 259092 231328
rect 199896 231288 259092 231316
rect 199896 231276 199902 231288
rect 259086 231276 259092 231288
rect 259144 231316 259150 231328
rect 262490 231316 262496 231328
rect 259144 231288 262496 231316
rect 259144 231276 259150 231288
rect 262490 231276 262496 231288
rect 262548 231276 262554 231328
rect 267182 231276 267188 231328
rect 267240 231316 267246 231328
rect 291194 231316 291200 231328
rect 267240 231288 291200 231316
rect 267240 231276 267246 231288
rect 291194 231276 291200 231288
rect 291252 231276 291258 231328
rect 164142 231208 164148 231260
rect 164200 231248 164206 231260
rect 223114 231248 223120 231260
rect 164200 231220 223120 231248
rect 164200 231208 164206 231220
rect 223114 231208 223120 231220
rect 223172 231208 223178 231260
rect 227346 231208 227352 231260
rect 227404 231248 227410 231260
rect 266170 231248 266176 231260
rect 227404 231220 266176 231248
rect 227404 231208 227410 231220
rect 266170 231208 266176 231220
rect 266228 231208 266234 231260
rect 266446 231208 266452 231260
rect 266504 231248 266510 231260
rect 291286 231248 291292 231260
rect 266504 231220 291292 231248
rect 266504 231208 266510 231220
rect 291286 231208 291292 231220
rect 291344 231208 291350 231260
rect 199930 231140 199936 231192
rect 199988 231180 199994 231192
rect 259638 231180 259644 231192
rect 199988 231152 259644 231180
rect 199988 231140 199994 231152
rect 259638 231140 259644 231152
rect 259696 231140 259702 231192
rect 262306 231140 262312 231192
rect 262364 231180 262370 231192
rect 263226 231180 263232 231192
rect 262364 231152 263232 231180
rect 262364 231140 262370 231152
rect 263226 231140 263232 231152
rect 263284 231140 263290 231192
rect 264514 231140 264520 231192
rect 264572 231180 264578 231192
rect 278958 231180 278964 231192
rect 264572 231152 278964 231180
rect 264572 231140 264578 231152
rect 278958 231140 278964 231152
rect 279016 231180 279022 231192
rect 279510 231180 279516 231192
rect 279016 231152 279516 231180
rect 279016 231140 279022 231152
rect 279510 231140 279516 231152
rect 279568 231140 279574 231192
rect 198642 231072 198648 231124
rect 198700 231112 198706 231124
rect 258534 231112 258540 231124
rect 198700 231084 258540 231112
rect 198700 231072 198706 231084
rect 258534 231072 258540 231084
rect 258592 231072 258598 231124
rect 258810 231072 258816 231124
rect 258868 231112 258874 231124
rect 280154 231112 280160 231124
rect 258868 231084 280160 231112
rect 258868 231072 258874 231084
rect 280154 231072 280160 231084
rect 280212 231112 280218 231124
rect 332686 231112 332692 231124
rect 280212 231084 332692 231112
rect 280212 231072 280218 231084
rect 332686 231072 332692 231084
rect 332744 231072 332750 231124
rect 248138 231004 248144 231056
rect 248196 231044 248202 231056
rect 276198 231044 276204 231056
rect 248196 231016 276204 231044
rect 248196 231004 248202 231016
rect 276198 231004 276204 231016
rect 276256 231004 276262 231056
rect 226610 230936 226616 230988
rect 226668 230976 226674 230988
rect 227530 230976 227536 230988
rect 226668 230948 227536 230976
rect 226668 230936 226674 230948
rect 227530 230936 227536 230948
rect 227588 230936 227594 230988
rect 232590 230936 232596 230988
rect 232648 230976 232654 230988
rect 233602 230976 233608 230988
rect 232648 230948 233608 230976
rect 232648 230936 232654 230948
rect 233602 230936 233608 230948
rect 233660 230936 233666 230988
rect 250898 230936 250904 230988
rect 250956 230976 250962 230988
rect 329834 230976 329840 230988
rect 250956 230948 329840 230976
rect 250956 230936 250962 230948
rect 329834 230936 329840 230948
rect 329892 230936 329898 230988
rect 251726 230868 251732 230920
rect 251784 230908 251790 230920
rect 252278 230908 252284 230920
rect 251784 230880 252284 230908
rect 251784 230868 251790 230880
rect 252278 230868 252284 230880
rect 252336 230868 252342 230920
rect 256786 230868 256792 230920
rect 256844 230908 256850 230920
rect 257062 230908 257068 230920
rect 256844 230880 257068 230908
rect 256844 230868 256850 230880
rect 257062 230868 257068 230880
rect 257120 230868 257126 230920
rect 258258 230704 258264 230716
rect 238726 230676 258264 230704
rect 199746 230528 199752 230580
rect 199804 230568 199810 230580
rect 238726 230568 238754 230676
rect 258258 230664 258264 230676
rect 258316 230664 258322 230716
rect 265434 230596 265440 230648
rect 265492 230636 265498 230648
rect 265894 230636 265900 230648
rect 265492 230608 265900 230636
rect 265492 230596 265498 230608
rect 265894 230596 265900 230608
rect 265952 230596 265958 230648
rect 199804 230540 238754 230568
rect 199804 230528 199810 230540
rect 239306 230528 239312 230580
rect 239364 230568 239370 230580
rect 239582 230568 239588 230580
rect 239364 230540 239588 230568
rect 239364 230528 239370 230540
rect 239582 230528 239588 230540
rect 239640 230528 239646 230580
rect 254486 230568 254492 230580
rect 244246 230540 254492 230568
rect 198458 230460 198464 230512
rect 198516 230500 198522 230512
rect 244246 230500 244274 230540
rect 254486 230528 254492 230540
rect 254544 230528 254550 230580
rect 249242 230500 249248 230512
rect 198516 230472 244274 230500
rect 248984 230472 249248 230500
rect 198516 230460 198522 230472
rect 228910 230392 228916 230444
rect 228968 230432 228974 230444
rect 235994 230432 236000 230444
rect 228968 230404 236000 230432
rect 228968 230392 228974 230404
rect 235994 230392 236000 230404
rect 236052 230392 236058 230444
rect 244090 230392 244096 230444
rect 244148 230432 244154 230444
rect 244826 230432 244832 230444
rect 244148 230404 244832 230432
rect 244148 230392 244154 230404
rect 244826 230392 244832 230404
rect 244884 230392 244890 230444
rect 245286 230392 245292 230444
rect 245344 230432 245350 230444
rect 248984 230432 249012 230472
rect 249242 230460 249248 230472
rect 249300 230460 249306 230512
rect 245344 230404 249012 230432
rect 245344 230392 245350 230404
rect 249058 230392 249064 230444
rect 249116 230432 249122 230444
rect 301498 230432 301504 230444
rect 249116 230404 301504 230432
rect 249116 230392 249122 230404
rect 301498 230392 301504 230404
rect 301556 230392 301562 230444
rect 305638 230392 305644 230444
rect 305696 230432 305702 230444
rect 306006 230432 306012 230444
rect 305696 230404 306012 230432
rect 305696 230392 305702 230404
rect 306006 230392 306012 230404
rect 306064 230392 306070 230444
rect 230014 230324 230020 230376
rect 230072 230364 230078 230376
rect 240962 230364 240968 230376
rect 230072 230336 240968 230364
rect 230072 230324 230078 230336
rect 240962 230324 240968 230336
rect 241020 230324 241026 230376
rect 243998 230324 244004 230376
rect 244056 230364 244062 230376
rect 304442 230364 304448 230376
rect 244056 230336 304448 230364
rect 244056 230324 244062 230336
rect 304442 230324 304448 230336
rect 304500 230324 304506 230376
rect 217778 230256 217784 230308
rect 217836 230296 217842 230308
rect 237098 230296 237104 230308
rect 217836 230268 237104 230296
rect 217836 230256 217842 230268
rect 237098 230256 237104 230268
rect 237156 230256 237162 230308
rect 241330 230256 241336 230308
rect 241388 230296 241394 230308
rect 300210 230296 300216 230308
rect 241388 230268 300216 230296
rect 241388 230256 241394 230268
rect 300210 230256 300216 230268
rect 300268 230256 300274 230308
rect 223206 230188 223212 230240
rect 223264 230228 223270 230240
rect 239122 230228 239128 230240
rect 223264 230200 239128 230228
rect 223264 230188 223270 230200
rect 239122 230188 239128 230200
rect 239180 230188 239186 230240
rect 239398 230188 239404 230240
rect 239456 230228 239462 230240
rect 240042 230228 240048 230240
rect 239456 230200 240048 230228
rect 239456 230188 239462 230200
rect 240042 230188 240048 230200
rect 240100 230228 240106 230240
rect 249058 230228 249064 230240
rect 240100 230200 249064 230228
rect 240100 230188 240106 230200
rect 249058 230188 249064 230200
rect 249116 230188 249122 230240
rect 305638 230228 305644 230240
rect 249168 230200 305644 230228
rect 212442 230120 212448 230172
rect 212500 230160 212506 230172
rect 239858 230160 239864 230172
rect 212500 230132 239864 230160
rect 212500 230120 212506 230132
rect 239858 230120 239864 230132
rect 239916 230120 239922 230172
rect 244734 230120 244740 230172
rect 244792 230160 244798 230172
rect 245286 230160 245292 230172
rect 244792 230132 245292 230160
rect 244792 230120 244798 230132
rect 245286 230120 245292 230132
rect 245344 230120 245350 230172
rect 247402 230120 247408 230172
rect 247460 230160 247466 230172
rect 249168 230160 249196 230200
rect 305638 230188 305644 230200
rect 305696 230188 305702 230240
rect 247460 230132 249196 230160
rect 247460 230120 247466 230132
rect 249242 230120 249248 230172
rect 249300 230160 249306 230172
rect 301682 230160 301688 230172
rect 249300 230132 301688 230160
rect 249300 230120 249306 230132
rect 301682 230120 301688 230132
rect 301740 230120 301746 230172
rect 235902 230092 235908 230104
rect 219406 230064 235908 230092
rect 162210 229780 162216 229832
rect 162268 229820 162274 229832
rect 219406 229820 219434 230064
rect 235902 230052 235908 230064
rect 235960 230092 235966 230104
rect 288250 230092 288256 230104
rect 235960 230064 288256 230092
rect 235960 230052 235966 230064
rect 288250 230052 288256 230064
rect 288308 230052 288314 230104
rect 235994 229984 236000 230036
rect 236052 230024 236058 230036
rect 237190 230024 237196 230036
rect 236052 229996 237196 230024
rect 236052 229984 236058 229996
rect 237190 229984 237196 229996
rect 237248 230024 237254 230036
rect 287974 230024 287980 230036
rect 237248 229996 287980 230024
rect 237248 229984 237254 229996
rect 287974 229984 287980 229996
rect 288032 229984 288038 230036
rect 239122 229916 239128 229968
rect 239180 229956 239186 229968
rect 247402 229956 247408 229968
rect 239180 229928 247408 229956
rect 239180 229916 239186 229928
rect 247402 229916 247408 229928
rect 247460 229916 247466 229968
rect 247586 229916 247592 229968
rect 247644 229956 247650 229968
rect 287790 229956 287796 229968
rect 247644 229928 287796 229956
rect 247644 229916 247650 229928
rect 287790 229916 287796 229928
rect 287848 229916 287854 229968
rect 225414 229848 225420 229900
rect 225472 229888 225478 229900
rect 225782 229888 225788 229900
rect 225472 229860 225788 229888
rect 225472 229848 225478 229860
rect 225782 229848 225788 229860
rect 225840 229848 225846 229900
rect 225966 229848 225972 229900
rect 226024 229888 226030 229900
rect 226024 229860 229094 229888
rect 226024 229848 226030 229860
rect 162268 229792 219434 229820
rect 162268 229780 162274 229792
rect 228358 229780 228364 229832
rect 228416 229820 228422 229832
rect 228726 229820 228732 229832
rect 228416 229792 228732 229820
rect 228416 229780 228422 229792
rect 228726 229780 228732 229792
rect 228784 229780 228790 229832
rect 229066 229820 229094 229860
rect 232958 229848 232964 229900
rect 233016 229888 233022 229900
rect 276658 229888 276664 229900
rect 233016 229860 276664 229888
rect 233016 229848 233022 229860
rect 276658 229848 276664 229860
rect 276716 229848 276722 229900
rect 229066 229792 236224 229820
rect 160922 229712 160928 229764
rect 160980 229752 160986 229764
rect 236086 229752 236092 229764
rect 160980 229724 236092 229752
rect 160980 229712 160986 229724
rect 236086 229712 236092 229724
rect 236144 229712 236150 229764
rect 236196 229752 236224 229792
rect 240870 229780 240876 229832
rect 240928 229820 240934 229832
rect 247586 229820 247592 229832
rect 240928 229792 247592 229820
rect 240928 229780 240934 229792
rect 247586 229780 247592 229792
rect 247644 229780 247650 229832
rect 249242 229780 249248 229832
rect 249300 229820 249306 229832
rect 279602 229820 279608 229832
rect 249300 229792 279608 229820
rect 249300 229780 249306 229792
rect 279602 229780 279608 229792
rect 279660 229780 279666 229832
rect 236546 229752 236552 229764
rect 236196 229724 236552 229752
rect 236546 229712 236552 229724
rect 236604 229752 236610 229764
rect 269850 229752 269856 229764
rect 236604 229724 246804 229752
rect 236604 229712 236610 229724
rect 235258 229644 235264 229696
rect 235316 229684 235322 229696
rect 240870 229684 240876 229696
rect 235316 229656 240876 229684
rect 235316 229644 235322 229656
rect 240870 229644 240876 229656
rect 240928 229644 240934 229696
rect 245286 229644 245292 229696
rect 245344 229684 245350 229696
rect 245562 229684 245568 229696
rect 245344 229656 245568 229684
rect 245344 229644 245350 229656
rect 245562 229644 245568 229656
rect 245620 229644 245626 229696
rect 245746 229644 245752 229696
rect 245804 229684 245810 229696
rect 246666 229684 246672 229696
rect 245804 229656 246672 229684
rect 245804 229644 245810 229656
rect 246666 229644 246672 229656
rect 246724 229644 246730 229696
rect 246776 229684 246804 229724
rect 251146 229724 269856 229752
rect 251146 229684 251174 229724
rect 269850 229712 269856 229724
rect 269908 229712 269914 229764
rect 274726 229712 274732 229764
rect 274784 229752 274790 229764
rect 275370 229752 275376 229764
rect 274784 229724 275376 229752
rect 274784 229712 274790 229724
rect 275370 229712 275376 229724
rect 275428 229712 275434 229764
rect 275922 229712 275928 229764
rect 275980 229752 275986 229764
rect 277026 229752 277032 229764
rect 275980 229724 277032 229752
rect 275980 229712 275986 229724
rect 277026 229712 277032 229724
rect 277084 229712 277090 229764
rect 273990 229684 273996 229696
rect 246776 229656 251174 229684
rect 253768 229656 273996 229684
rect 251266 229576 251272 229628
rect 251324 229616 251330 229628
rect 252462 229616 252468 229628
rect 251324 229588 252468 229616
rect 251324 229576 251330 229588
rect 252462 229576 252468 229588
rect 252520 229576 252526 229628
rect 253768 229616 253796 229656
rect 273990 229644 273996 229656
rect 274048 229644 274054 229696
rect 274726 229616 274732 229628
rect 253584 229588 253796 229616
rect 253860 229588 274732 229616
rect 212350 229508 212356 229560
rect 212408 229548 212414 229560
rect 236730 229548 236736 229560
rect 212408 229520 236736 229548
rect 212408 229508 212414 229520
rect 236730 229508 236736 229520
rect 236788 229508 236794 229560
rect 239858 229508 239864 229560
rect 239916 229548 239922 229560
rect 249242 229548 249248 229560
rect 239916 229520 249248 229548
rect 239916 229508 239922 229520
rect 249242 229508 249248 229520
rect 249300 229508 249306 229560
rect 247494 229440 247500 229492
rect 247552 229480 247558 229492
rect 248322 229480 248328 229492
rect 247552 229452 248328 229480
rect 247552 229440 247558 229452
rect 248322 229440 248328 229452
rect 248380 229440 248386 229492
rect 245010 229372 245016 229424
rect 245068 229412 245074 229424
rect 253584 229412 253612 229588
rect 245068 229384 253612 229412
rect 245068 229372 245074 229384
rect 248598 229304 248604 229356
rect 248656 229344 248662 229356
rect 249242 229344 249248 229356
rect 248656 229316 249248 229344
rect 248656 229304 248662 229316
rect 249242 229304 249248 229316
rect 249300 229304 249306 229356
rect 249518 229304 249524 229356
rect 249576 229344 249582 229356
rect 253860 229344 253888 229588
rect 274726 229576 274732 229588
rect 274784 229576 274790 229628
rect 262858 229508 262864 229560
rect 262916 229548 262922 229560
rect 280246 229548 280252 229560
rect 262916 229520 280252 229548
rect 262916 229508 262922 229520
rect 280246 229508 280252 229520
rect 280304 229508 280310 229560
rect 249576 229316 253888 229344
rect 249576 229304 249582 229316
rect 252738 229236 252744 229288
rect 252796 229276 252802 229288
rect 253750 229276 253756 229288
rect 252796 229248 253756 229276
rect 252796 229236 252802 229248
rect 253750 229236 253756 229248
rect 253808 229236 253814 229288
rect 222930 229168 222936 229220
rect 222988 229208 222994 229220
rect 236454 229208 236460 229220
rect 222988 229180 236460 229208
rect 222988 229168 222994 229180
rect 236454 229168 236460 229180
rect 236512 229168 236518 229220
rect 227530 229100 227536 229152
rect 227588 229140 227594 229152
rect 244090 229140 244096 229152
rect 227588 229112 244096 229140
rect 227588 229100 227594 229112
rect 244090 229100 244096 229112
rect 244148 229100 244154 229152
rect 271138 229100 271144 229152
rect 271196 229140 271202 229152
rect 277394 229140 277400 229152
rect 271196 229112 277400 229140
rect 271196 229100 271202 229112
rect 277394 229100 277400 229112
rect 277452 229100 277458 229152
rect 208302 229032 208308 229084
rect 208360 229072 208366 229084
rect 230290 229072 230296 229084
rect 208360 229044 230296 229072
rect 208360 229032 208366 229044
rect 230290 229032 230296 229044
rect 230348 229032 230354 229084
rect 258442 229032 258448 229084
rect 258500 229072 258506 229084
rect 338206 229072 338212 229084
rect 258500 229044 338212 229072
rect 258500 229032 258506 229044
rect 338206 229032 338212 229044
rect 338264 229032 338270 229084
rect 230566 228964 230572 229016
rect 230624 229004 230630 229016
rect 231302 229004 231308 229016
rect 230624 228976 231308 229004
rect 230624 228964 230630 228976
rect 231302 228964 231308 228976
rect 231360 228964 231366 229016
rect 233326 228964 233332 229016
rect 233384 229004 233390 229016
rect 233786 229004 233792 229016
rect 233384 228976 233792 229004
rect 233384 228964 233390 228976
rect 233786 228964 233792 228976
rect 233844 228964 233850 229016
rect 260098 228964 260104 229016
rect 260156 229004 260162 229016
rect 335354 229004 335360 229016
rect 260156 228976 335360 229004
rect 260156 228964 260162 228976
rect 335354 228964 335360 228976
rect 335412 228964 335418 229016
rect 161566 228896 161572 228948
rect 161624 228936 161630 228948
rect 215202 228936 215208 228948
rect 161624 228908 215208 228936
rect 161624 228896 161630 228908
rect 215202 228896 215208 228908
rect 215260 228896 215266 228948
rect 231118 228896 231124 228948
rect 231176 228936 231182 228948
rect 236822 228936 236828 228948
rect 231176 228908 236828 228936
rect 231176 228896 231182 228908
rect 236822 228896 236828 228908
rect 236880 228896 236886 228948
rect 263502 228896 263508 228948
rect 263560 228936 263566 228948
rect 327258 228936 327264 228948
rect 263560 228908 327264 228936
rect 263560 228896 263566 228908
rect 327258 228896 327264 228908
rect 327316 228896 327322 228948
rect 154022 228828 154028 228880
rect 154080 228868 154086 228880
rect 208302 228868 208308 228880
rect 154080 228840 208308 228868
rect 154080 228828 154086 228840
rect 208302 228828 208308 228840
rect 208360 228828 208366 228880
rect 299014 228868 299020 228880
rect 244246 228840 299020 228868
rect 152734 228760 152740 228812
rect 152792 228800 152798 228812
rect 209498 228800 209504 228812
rect 152792 228772 209504 228800
rect 152792 228760 152798 228772
rect 209498 228760 209504 228772
rect 209556 228760 209562 228812
rect 213730 228760 213736 228812
rect 213788 228800 213794 228812
rect 239030 228800 239036 228812
rect 213788 228772 239036 228800
rect 213788 228760 213794 228772
rect 239030 228760 239036 228772
rect 239088 228800 239094 228812
rect 244246 228800 244274 228840
rect 299014 228828 299020 228840
rect 299072 228828 299078 228880
rect 239088 228772 244274 228800
rect 239088 228760 239094 228772
rect 249150 228760 249156 228812
rect 249208 228800 249214 228812
rect 258442 228800 258448 228812
rect 249208 228772 258448 228800
rect 249208 228760 249214 228772
rect 258442 228760 258448 228772
rect 258500 228760 258506 228812
rect 265618 228760 265624 228812
rect 265676 228800 265682 228812
rect 268194 228800 268200 228812
rect 265676 228772 268200 228800
rect 265676 228760 265682 228772
rect 268194 228760 268200 228772
rect 268252 228800 268258 228812
rect 327902 228800 327908 228812
rect 268252 228772 327908 228800
rect 268252 228760 268258 228772
rect 327902 228760 327908 228772
rect 327960 228760 327966 228812
rect 259914 228732 259920 228744
rect 258046 228704 259920 228732
rect 155586 228624 155592 228676
rect 155644 228664 155650 228676
rect 225598 228664 225604 228676
rect 155644 228636 225604 228664
rect 155644 228624 155650 228636
rect 225598 228624 225604 228636
rect 225656 228624 225662 228676
rect 239674 228624 239680 228676
rect 239732 228664 239738 228676
rect 258046 228664 258074 228704
rect 259914 228692 259920 228704
rect 259972 228732 259978 228744
rect 301866 228732 301872 228744
rect 259972 228704 301872 228732
rect 259972 228692 259978 228704
rect 301866 228692 301872 228704
rect 301924 228692 301930 228744
rect 239732 228636 258074 228664
rect 239732 228624 239738 228636
rect 264698 228624 264704 228676
rect 264756 228664 264762 228676
rect 325142 228664 325148 228676
rect 264756 228636 325148 228664
rect 264756 228624 264762 228636
rect 325142 228624 325148 228636
rect 325200 228624 325206 228676
rect 201218 228556 201224 228608
rect 201276 228596 201282 228608
rect 271874 228596 271880 228608
rect 201276 228568 271880 228596
rect 201276 228556 201282 228568
rect 271874 228556 271880 228568
rect 271932 228556 271938 228608
rect 152826 228488 152832 228540
rect 152884 228528 152890 228540
rect 225230 228528 225236 228540
rect 152884 228500 225236 228528
rect 152884 228488 152890 228500
rect 225230 228488 225236 228500
rect 225288 228488 225294 228540
rect 234430 228488 234436 228540
rect 234488 228528 234494 228540
rect 295242 228528 295248 228540
rect 234488 228500 295248 228528
rect 234488 228488 234494 228500
rect 295242 228488 295248 228500
rect 295300 228488 295306 228540
rect 197906 228420 197912 228472
rect 197964 228460 197970 228472
rect 271966 228460 271972 228472
rect 197964 228432 271972 228460
rect 197964 228420 197970 228432
rect 271966 228420 271972 228432
rect 272024 228420 272030 228472
rect 160830 228352 160836 228404
rect 160888 228392 160894 228404
rect 237834 228392 237840 228404
rect 160888 228364 237840 228392
rect 160888 228352 160894 228364
rect 237834 228352 237840 228364
rect 237892 228352 237898 228404
rect 239766 228352 239772 228404
rect 239824 228392 239830 228404
rect 260098 228392 260104 228404
rect 239824 228364 260104 228392
rect 239824 228352 239830 228364
rect 260098 228352 260104 228364
rect 260156 228352 260162 228404
rect 266538 228352 266544 228404
rect 266596 228392 266602 228404
rect 267182 228392 267188 228404
rect 266596 228364 267188 228392
rect 266596 228352 266602 228364
rect 267182 228352 267188 228364
rect 267240 228352 267246 228404
rect 232682 228284 232688 228336
rect 232740 228324 232746 228336
rect 288158 228324 288164 228336
rect 232740 228296 288164 228324
rect 232740 228284 232746 228296
rect 288158 228284 288164 228296
rect 288216 228284 288222 228336
rect 233694 228216 233700 228268
rect 233752 228256 233758 228268
rect 234154 228256 234160 228268
rect 233752 228228 234160 228256
rect 233752 228216 233758 228228
rect 234154 228216 234160 228228
rect 234212 228216 234218 228268
rect 235534 228216 235540 228268
rect 235592 228256 235598 228268
rect 286502 228256 286508 228268
rect 235592 228228 286508 228256
rect 235592 228216 235598 228228
rect 286502 228216 286508 228228
rect 286560 228216 286566 228268
rect 236454 228148 236460 228200
rect 236512 228188 236518 228200
rect 273622 228188 273628 228200
rect 236512 228160 273628 228188
rect 236512 228148 236518 228160
rect 273622 228148 273628 228160
rect 273680 228148 273686 228200
rect 202598 228080 202604 228132
rect 202656 228120 202662 228132
rect 272426 228120 272432 228132
rect 202656 228092 272432 228120
rect 202656 228080 202662 228092
rect 272426 228080 272432 228092
rect 272484 228080 272490 228132
rect 234798 227740 234804 227792
rect 234856 227780 234862 227792
rect 235534 227780 235540 227792
rect 234856 227752 235540 227780
rect 234856 227740 234862 227752
rect 235534 227740 235540 227752
rect 235592 227740 235598 227792
rect 262858 227740 262864 227792
rect 262916 227780 262922 227792
rect 263502 227780 263508 227792
rect 262916 227752 263508 227780
rect 262916 227740 262922 227752
rect 263502 227740 263508 227752
rect 263560 227740 263566 227792
rect 260558 227712 260564 227724
rect 258046 227684 260564 227712
rect 215110 227536 215116 227588
rect 215168 227576 215174 227588
rect 258046 227576 258074 227684
rect 260558 227672 260564 227684
rect 260616 227712 260622 227724
rect 321002 227712 321008 227724
rect 260616 227684 321008 227712
rect 260616 227672 260622 227684
rect 321002 227672 321008 227684
rect 321060 227672 321066 227724
rect 262950 227604 262956 227656
rect 263008 227644 263014 227656
rect 323854 227644 323860 227656
rect 263008 227616 323860 227644
rect 263008 227604 263014 227616
rect 323854 227604 323860 227616
rect 323912 227604 323918 227656
rect 215168 227548 258074 227576
rect 215168 227536 215174 227548
rect 263226 227536 263232 227588
rect 263284 227576 263290 227588
rect 323762 227576 323768 227588
rect 263284 227548 323768 227576
rect 263284 227536 263290 227548
rect 323762 227536 323768 227548
rect 323820 227536 323826 227588
rect 228174 227468 228180 227520
rect 228232 227508 228238 227520
rect 228634 227508 228640 227520
rect 228232 227480 228640 227508
rect 228232 227468 228238 227480
rect 228634 227468 228640 227480
rect 228692 227468 228698 227520
rect 260926 227468 260932 227520
rect 260984 227508 260990 227520
rect 321646 227508 321652 227520
rect 260984 227480 321652 227508
rect 260984 227468 260990 227480
rect 321646 227468 321652 227480
rect 321704 227468 321710 227520
rect 234706 227400 234712 227452
rect 234764 227440 234770 227452
rect 294598 227440 294604 227452
rect 234764 227412 294604 227440
rect 234764 227400 234770 227412
rect 294598 227400 294604 227412
rect 294656 227400 294662 227452
rect 239306 227372 239312 227384
rect 238726 227344 239312 227372
rect 223022 227264 223028 227316
rect 223080 227304 223086 227316
rect 238726 227304 238754 227344
rect 239306 227332 239312 227344
rect 239364 227372 239370 227384
rect 289170 227372 289176 227384
rect 239364 227344 289176 227372
rect 239364 227332 239370 227344
rect 289170 227332 289176 227344
rect 289228 227332 289234 227384
rect 223080 227276 238754 227304
rect 223080 227264 223086 227276
rect 251082 227264 251088 227316
rect 251140 227304 251146 227316
rect 278222 227304 278228 227316
rect 251140 227276 278228 227304
rect 251140 227264 251146 227276
rect 278222 227264 278228 227276
rect 278280 227264 278286 227316
rect 287514 227264 287520 227316
rect 287572 227304 287578 227316
rect 336826 227304 336832 227316
rect 287572 227276 336832 227304
rect 287572 227264 287578 227276
rect 336826 227264 336832 227276
rect 336884 227264 336890 227316
rect 226978 227196 226984 227248
rect 227036 227236 227042 227248
rect 257062 227236 257068 227248
rect 227036 227208 257068 227236
rect 227036 227196 227042 227208
rect 257062 227196 257068 227208
rect 257120 227196 257126 227248
rect 258350 227196 258356 227248
rect 258408 227236 258414 227248
rect 292666 227236 292672 227248
rect 258408 227208 292672 227236
rect 258408 227196 258414 227208
rect 292666 227196 292672 227208
rect 292724 227196 292730 227248
rect 256602 227128 256608 227180
rect 256660 227168 256666 227180
rect 282362 227168 282368 227180
rect 256660 227140 282368 227168
rect 256660 227128 256666 227140
rect 282362 227128 282368 227140
rect 282420 227128 282426 227180
rect 234338 227060 234344 227112
rect 234396 227100 234402 227112
rect 235994 227100 236000 227112
rect 234396 227072 236000 227100
rect 234396 227060 234402 227072
rect 235994 227060 236000 227072
rect 236052 227100 236058 227112
rect 280890 227100 280896 227112
rect 236052 227072 280896 227100
rect 236052 227060 236058 227072
rect 280890 227060 280896 227072
rect 280948 227060 280954 227112
rect 333054 227100 333060 227112
rect 291028 227072 333060 227100
rect 155402 226992 155408 227044
rect 155460 227032 155466 227044
rect 210970 227032 210976 227044
rect 155460 227004 210976 227032
rect 155460 226992 155466 227004
rect 210970 226992 210976 227004
rect 211028 226992 211034 227044
rect 211706 226992 211712 227044
rect 211764 227032 211770 227044
rect 269390 227032 269396 227044
rect 211764 227004 269396 227032
rect 211764 226992 211770 227004
rect 269390 226992 269396 227004
rect 269448 226992 269454 227044
rect 255774 226924 255780 226976
rect 255832 226964 255838 226976
rect 289262 226964 289268 226976
rect 255832 226936 289268 226964
rect 255832 226924 255838 226936
rect 289262 226924 289268 226936
rect 289320 226964 289326 226976
rect 291028 226964 291056 227072
rect 333054 227060 333060 227072
rect 333112 227060 333118 227112
rect 292666 226992 292672 227044
rect 292724 227032 292730 227044
rect 293218 227032 293224 227044
rect 292724 227004 293224 227032
rect 292724 226992 292730 227004
rect 293218 226992 293224 227004
rect 293276 227032 293282 227044
rect 336918 227032 336924 227044
rect 293276 227004 336924 227032
rect 293276 226992 293282 227004
rect 336918 226992 336924 227004
rect 336976 226992 336982 227044
rect 289320 226936 291056 226964
rect 289320 226924 289326 226936
rect 239858 226856 239864 226908
rect 239916 226896 239922 226908
rect 265526 226896 265532 226908
rect 239916 226868 265532 226896
rect 239916 226856 239922 226868
rect 265526 226856 265532 226868
rect 265584 226856 265590 226908
rect 265802 226856 265808 226908
rect 265860 226896 265866 226908
rect 285766 226896 285772 226908
rect 265860 226868 285772 226896
rect 265860 226856 265866 226868
rect 285766 226856 285772 226868
rect 285824 226856 285830 226908
rect 262030 226788 262036 226840
rect 262088 226828 262094 226840
rect 281994 226828 282000 226840
rect 262088 226800 282000 226828
rect 262088 226788 262094 226800
rect 281994 226788 282000 226800
rect 282052 226788 282058 226840
rect 250622 226720 250628 226772
rect 250680 226760 250686 226772
rect 251082 226760 251088 226772
rect 250680 226732 251088 226760
rect 250680 226720 250686 226732
rect 251082 226720 251088 226732
rect 251140 226720 251146 226772
rect 265710 226652 265716 226704
rect 265768 226692 265774 226704
rect 266262 226692 266268 226704
rect 265768 226664 266268 226692
rect 265768 226652 265774 226664
rect 266262 226652 266268 226664
rect 266320 226652 266326 226704
rect 285766 226652 285772 226704
rect 285824 226692 285830 226704
rect 286962 226692 286968 226704
rect 285824 226664 286968 226692
rect 285824 226652 285830 226664
rect 286962 226652 286968 226664
rect 287020 226652 287026 226704
rect 250806 226584 250812 226636
rect 250864 226624 250870 226636
rect 251082 226624 251088 226636
rect 250864 226596 251088 226624
rect 250864 226584 250870 226596
rect 251082 226584 251088 226596
rect 251140 226584 251146 226636
rect 234706 226516 234712 226568
rect 234764 226556 234770 226568
rect 235442 226556 235448 226568
rect 234764 226528 235448 226556
rect 234764 226516 234770 226528
rect 235442 226516 235448 226528
rect 235500 226516 235506 226568
rect 260098 226312 260104 226364
rect 260156 226352 260162 226364
rect 260926 226352 260932 226364
rect 260156 226324 260932 226352
rect 260156 226312 260162 226324
rect 260926 226312 260932 226324
rect 260984 226312 260990 226364
rect 281534 226312 281540 226364
rect 281592 226352 281598 226364
rect 281994 226352 282000 226364
rect 281592 226324 282000 226352
rect 281592 226312 281598 226324
rect 281994 226312 282000 226324
rect 282052 226312 282058 226364
rect 287514 226312 287520 226364
rect 287572 226352 287578 226364
rect 287790 226352 287796 226364
rect 287572 226324 287796 226352
rect 287572 226312 287578 226324
rect 287790 226312 287796 226324
rect 287848 226312 287854 226364
rect 202690 226244 202696 226296
rect 202748 226284 202754 226296
rect 227070 226284 227076 226296
rect 202748 226256 227076 226284
rect 202748 226244 202754 226256
rect 227070 226244 227076 226256
rect 227128 226244 227134 226296
rect 249886 226244 249892 226296
rect 249944 226284 249950 226296
rect 250530 226284 250536 226296
rect 249944 226256 250536 226284
rect 249944 226244 249950 226256
rect 250530 226244 250536 226256
rect 250588 226244 250594 226296
rect 258258 226244 258264 226296
rect 258316 226284 258322 226296
rect 345014 226284 345020 226296
rect 258316 226256 345020 226284
rect 258316 226244 258322 226256
rect 345014 226244 345020 226256
rect 345072 226244 345078 226296
rect 266262 226176 266268 226228
rect 266320 226216 266326 226228
rect 342254 226216 342260 226228
rect 266320 226188 342260 226216
rect 266320 226176 266326 226188
rect 342254 226176 342260 226188
rect 342312 226176 342318 226228
rect 241146 226108 241152 226160
rect 241204 226148 241210 226160
rect 301774 226148 301780 226160
rect 241204 226120 301780 226148
rect 241204 226108 241210 226120
rect 301774 226108 301780 226120
rect 301832 226108 301838 226160
rect 246298 226040 246304 226092
rect 246356 226080 246362 226092
rect 307018 226080 307024 226092
rect 246356 226052 307024 226080
rect 246356 226040 246362 226052
rect 307018 226040 307024 226052
rect 307076 226040 307082 226092
rect 245470 225972 245476 226024
rect 245528 226012 245534 226024
rect 305730 226012 305736 226024
rect 245528 225984 305736 226012
rect 245528 225972 245534 225984
rect 305730 225972 305736 225984
rect 305788 225972 305794 226024
rect 250438 225904 250444 225956
rect 250496 225944 250502 225956
rect 309962 225944 309968 225956
rect 250496 225916 309968 225944
rect 250496 225904 250502 225916
rect 309962 225904 309968 225916
rect 310020 225904 310026 225956
rect 245194 225836 245200 225888
rect 245252 225876 245258 225888
rect 245470 225876 245476 225888
rect 245252 225848 245476 225876
rect 245252 225836 245258 225848
rect 245470 225836 245476 225848
rect 245528 225836 245534 225888
rect 250530 225836 250536 225888
rect 250588 225876 250594 225888
rect 310054 225876 310060 225888
rect 250588 225848 310060 225876
rect 250588 225836 250594 225848
rect 310054 225836 310060 225848
rect 310112 225836 310118 225888
rect 255590 225768 255596 225820
rect 255648 225808 255654 225820
rect 255958 225808 255964 225820
rect 255648 225780 255964 225808
rect 255648 225768 255654 225780
rect 255958 225768 255964 225780
rect 256016 225808 256022 225820
rect 315666 225808 315672 225820
rect 256016 225780 315672 225808
rect 256016 225768 256022 225780
rect 315666 225768 315672 225780
rect 315724 225768 315730 225820
rect 243906 225700 243912 225752
rect 243964 225740 243970 225752
rect 302970 225740 302976 225752
rect 243964 225712 302976 225740
rect 243964 225700 243970 225712
rect 302970 225700 302976 225712
rect 303028 225700 303034 225752
rect 234246 225632 234252 225684
rect 234304 225672 234310 225684
rect 240502 225672 240508 225684
rect 234304 225644 240508 225672
rect 234304 225632 234310 225644
rect 240502 225632 240508 225644
rect 240560 225672 240566 225684
rect 295978 225672 295984 225684
rect 240560 225644 295984 225672
rect 240560 225632 240566 225644
rect 295978 225632 295984 225644
rect 296036 225632 296042 225684
rect 156782 225564 156788 225616
rect 156840 225604 156846 225616
rect 202690 225604 202696 225616
rect 156840 225576 202696 225604
rect 156840 225564 156846 225576
rect 202690 225564 202696 225576
rect 202748 225564 202754 225616
rect 244090 225564 244096 225616
rect 244148 225604 244154 225616
rect 296714 225604 296720 225616
rect 244148 225576 296720 225604
rect 244148 225564 244154 225576
rect 296714 225564 296720 225576
rect 296772 225604 296778 225616
rect 297358 225604 297364 225616
rect 296772 225576 297364 225604
rect 296772 225564 296778 225576
rect 297358 225564 297364 225576
rect 297416 225564 297422 225616
rect 241698 225496 241704 225548
rect 241756 225536 241762 225548
rect 242710 225536 242716 225548
rect 241756 225508 242716 225536
rect 241756 225496 241762 225508
rect 242710 225496 242716 225508
rect 242768 225536 242774 225548
rect 285030 225536 285036 225548
rect 242768 225508 285036 225536
rect 242768 225496 242774 225508
rect 285030 225496 285036 225508
rect 285088 225496 285094 225548
rect 242526 225428 242532 225480
rect 242584 225468 242590 225480
rect 284110 225468 284116 225480
rect 242584 225440 284116 225468
rect 242584 225428 242590 225440
rect 284110 225428 284116 225440
rect 284168 225428 284174 225480
rect 243814 225360 243820 225412
rect 243872 225400 243878 225412
rect 282638 225400 282644 225412
rect 243872 225372 282644 225400
rect 243872 225360 243878 225372
rect 282638 225360 282644 225372
rect 282696 225360 282702 225412
rect 243538 225020 243544 225072
rect 243596 225060 243602 225072
rect 243814 225060 243820 225072
rect 243596 225032 243820 225060
rect 243596 225020 243602 225032
rect 243814 225020 243820 225032
rect 243872 225020 243878 225072
rect 240870 224952 240876 225004
rect 240928 224992 240934 225004
rect 241146 224992 241152 225004
rect 240928 224964 241152 224992
rect 240928 224952 240934 224964
rect 241146 224952 241152 224964
rect 241204 224952 241210 225004
rect 242158 224952 242164 225004
rect 242216 224992 242222 225004
rect 242526 224992 242532 225004
rect 242216 224964 242532 224992
rect 242216 224952 242222 224964
rect 242526 224952 242532 224964
rect 242584 224952 242590 225004
rect 243630 224952 243636 225004
rect 243688 224992 243694 225004
rect 243906 224992 243912 225004
rect 243688 224964 243912 224992
rect 243688 224952 243694 224964
rect 243906 224952 243912 224964
rect 243964 224952 243970 225004
rect 248966 224952 248972 225004
rect 249024 224992 249030 225004
rect 249334 224992 249340 225004
rect 249024 224964 249340 224992
rect 249024 224952 249030 224964
rect 249334 224952 249340 224964
rect 249392 224952 249398 225004
rect 222010 224884 222016 224936
rect 222068 224924 222074 224936
rect 298002 224924 298008 224936
rect 222068 224896 298008 224924
rect 222068 224884 222074 224896
rect 298002 224884 298008 224896
rect 298060 224884 298066 224936
rect 236730 224816 236736 224868
rect 236788 224856 236794 224868
rect 237282 224856 237288 224868
rect 236788 224828 237288 224856
rect 236788 224816 236794 224828
rect 237282 224816 237288 224828
rect 237340 224856 237346 224868
rect 301590 224856 301596 224868
rect 237340 224828 301596 224856
rect 237340 224816 237346 224828
rect 301590 224816 301596 224828
rect 301648 224816 301654 224868
rect 234154 224748 234160 224800
rect 234212 224788 234218 224800
rect 298278 224788 298284 224800
rect 234212 224760 298284 224788
rect 234212 224748 234218 224760
rect 298278 224748 298284 224760
rect 298336 224748 298342 224800
rect 225874 224680 225880 224732
rect 225932 224720 225938 224732
rect 245102 224720 245108 224732
rect 225932 224692 245108 224720
rect 225932 224680 225938 224692
rect 245102 224680 245108 224692
rect 245160 224680 245166 224732
rect 252002 224680 252008 224732
rect 252060 224720 252066 224732
rect 312814 224720 312820 224732
rect 252060 224692 312820 224720
rect 252060 224680 252066 224692
rect 312814 224680 312820 224692
rect 312872 224680 312878 224732
rect 238570 224652 238576 224664
rect 219406 224624 238576 224652
rect 209406 224272 209412 224324
rect 209464 224312 209470 224324
rect 219406 224312 219434 224624
rect 238570 224612 238576 224624
rect 238628 224652 238634 224664
rect 298738 224652 298744 224664
rect 238628 224624 298744 224652
rect 238628 224612 238634 224624
rect 298738 224612 298744 224624
rect 298796 224612 298802 224664
rect 239582 224544 239588 224596
rect 239640 224584 239646 224596
rect 299566 224584 299572 224596
rect 239640 224556 299572 224584
rect 239640 224544 239646 224556
rect 299566 224544 299572 224556
rect 299624 224544 299630 224596
rect 240962 224476 240968 224528
rect 241020 224516 241026 224528
rect 300118 224516 300124 224528
rect 241020 224488 300124 224516
rect 241020 224476 241026 224488
rect 300118 224476 300124 224488
rect 300176 224476 300182 224528
rect 232866 224408 232872 224460
rect 232924 224448 232930 224460
rect 285214 224448 285220 224460
rect 232924 224420 285220 224448
rect 232924 224408 232930 224420
rect 285214 224408 285220 224420
rect 285272 224408 285278 224460
rect 243722 224340 243728 224392
rect 243780 224380 243786 224392
rect 293310 224380 293316 224392
rect 243780 224352 293316 224380
rect 243780 224340 243786 224352
rect 293310 224340 293316 224352
rect 293368 224340 293374 224392
rect 209464 224284 219434 224312
rect 209464 224272 209470 224284
rect 240686 224272 240692 224324
rect 240744 224312 240750 224324
rect 242894 224312 242900 224324
rect 240744 224284 242900 224312
rect 240744 224272 240750 224284
rect 242894 224272 242900 224284
rect 242952 224312 242958 224324
rect 297450 224312 297456 224324
rect 242952 224284 297456 224312
rect 242952 224272 242958 224284
rect 297450 224272 297456 224284
rect 297508 224272 297514 224324
rect 160738 224204 160744 224256
rect 160796 224244 160802 224256
rect 237650 224244 237656 224256
rect 160796 224216 237656 224244
rect 160796 224204 160802 224216
rect 237650 224204 237656 224216
rect 237708 224204 237714 224256
rect 240778 224204 240784 224256
rect 240836 224244 240842 224256
rect 241238 224244 241244 224256
rect 240836 224216 241244 224244
rect 240836 224204 240842 224216
rect 241238 224204 241244 224216
rect 241296 224204 241302 224256
rect 242066 224204 242072 224256
rect 242124 224244 242130 224256
rect 244274 224244 244280 224256
rect 242124 224216 244280 224244
rect 242124 224204 242130 224216
rect 244274 224204 244280 224216
rect 244332 224244 244338 224256
rect 302878 224244 302884 224256
rect 244332 224216 302884 224244
rect 244332 224204 244338 224216
rect 302878 224204 302884 224216
rect 302936 224204 302942 224256
rect 230198 224136 230204 224188
rect 230256 224176 230262 224188
rect 230658 224176 230664 224188
rect 230256 224148 230664 224176
rect 230256 224136 230262 224148
rect 230658 224136 230664 224148
rect 230716 224136 230722 224188
rect 238202 224136 238208 224188
rect 238260 224176 238266 224188
rect 283742 224176 283748 224188
rect 238260 224148 283748 224176
rect 238260 224136 238266 224148
rect 283742 224136 283748 224148
rect 283800 224136 283806 224188
rect 241238 224068 241244 224120
rect 241296 224108 241302 224120
rect 286686 224108 286692 224120
rect 241296 224080 286692 224108
rect 241296 224068 241302 224080
rect 286686 224068 286692 224080
rect 286744 224068 286750 224120
rect 238018 224000 238024 224052
rect 238076 224040 238082 224052
rect 247218 224040 247224 224052
rect 238076 224012 247224 224040
rect 238076 224000 238082 224012
rect 247218 224000 247224 224012
rect 247276 224000 247282 224052
rect 252830 224000 252836 224052
rect 252888 224040 252894 224052
rect 253290 224040 253296 224052
rect 252888 224012 253296 224040
rect 252888 224000 252894 224012
rect 253290 224000 253296 224012
rect 253348 224040 253354 224052
rect 272610 224040 272616 224052
rect 253348 224012 272616 224040
rect 253348 224000 253354 224012
rect 272610 224000 272616 224012
rect 272668 224000 272674 224052
rect 264330 223932 264336 223984
rect 264388 223972 264394 223984
rect 264606 223972 264612 223984
rect 264388 223944 264612 223972
rect 264388 223932 264394 223944
rect 264606 223932 264612 223944
rect 264664 223932 264670 223984
rect 264146 223864 264152 223916
rect 264204 223904 264210 223916
rect 264422 223904 264428 223916
rect 264204 223876 264428 223904
rect 264204 223864 264210 223876
rect 264422 223864 264428 223876
rect 264480 223864 264486 223916
rect 251450 223524 251456 223576
rect 251508 223564 251514 223576
rect 252186 223564 252192 223576
rect 251508 223536 252192 223564
rect 251508 223524 251514 223536
rect 252186 223524 252192 223536
rect 252244 223524 252250 223576
rect 258994 223524 259000 223576
rect 259052 223564 259058 223576
rect 319714 223564 319720 223576
rect 259052 223536 319720 223564
rect 259052 223524 259058 223536
rect 319714 223524 319720 223536
rect 319772 223524 319778 223576
rect 251358 223456 251364 223508
rect 251416 223496 251422 223508
rect 251910 223496 251916 223508
rect 251416 223468 251916 223496
rect 251416 223456 251422 223468
rect 251910 223456 251916 223468
rect 251968 223456 251974 223508
rect 256878 223456 256884 223508
rect 256936 223496 256942 223508
rect 257338 223496 257344 223508
rect 256936 223468 257344 223496
rect 256936 223456 256942 223468
rect 257338 223456 257344 223468
rect 257396 223496 257402 223508
rect 318334 223496 318340 223508
rect 257396 223468 318340 223496
rect 257396 223456 257402 223468
rect 318334 223456 318340 223468
rect 318392 223456 318398 223508
rect 256694 223388 256700 223440
rect 256752 223428 256758 223440
rect 257430 223428 257436 223440
rect 256752 223400 257436 223428
rect 256752 223388 256758 223400
rect 257430 223388 257436 223400
rect 257488 223428 257494 223440
rect 318242 223428 318248 223440
rect 257488 223400 318248 223428
rect 257488 223388 257494 223400
rect 318242 223388 318248 223400
rect 318300 223388 318306 223440
rect 256050 223320 256056 223372
rect 256108 223360 256114 223372
rect 256418 223360 256424 223372
rect 256108 223332 256424 223360
rect 256108 223320 256114 223332
rect 256418 223320 256424 223332
rect 256476 223360 256482 223372
rect 316678 223360 316684 223372
rect 256476 223332 316684 223360
rect 256476 223320 256482 223332
rect 316678 223320 316684 223332
rect 316736 223320 316742 223372
rect 260466 223252 260472 223304
rect 260524 223292 260530 223304
rect 319438 223292 319444 223304
rect 260524 223264 319444 223292
rect 260524 223252 260530 223264
rect 319438 223252 319444 223264
rect 319496 223252 319502 223304
rect 258902 223184 258908 223236
rect 258960 223224 258966 223236
rect 318150 223224 318156 223236
rect 258960 223196 318156 223224
rect 258960 223184 258966 223196
rect 318150 223184 318156 223196
rect 318208 223184 318214 223236
rect 251910 223116 251916 223168
rect 251968 223156 251974 223168
rect 311250 223156 311256 223168
rect 251968 223128 311256 223156
rect 251968 223116 251974 223128
rect 311250 223116 311256 223128
rect 311308 223116 311314 223168
rect 252186 223048 252192 223100
rect 252244 223088 252250 223100
rect 311158 223088 311164 223100
rect 252244 223060 311164 223088
rect 252244 223048 252250 223060
rect 311158 223048 311164 223060
rect 311216 223048 311222 223100
rect 226610 223020 226616 223032
rect 224926 222992 226616 223020
rect 155494 222844 155500 222896
rect 155552 222884 155558 222896
rect 224926 222884 224954 222992
rect 226610 222980 226616 222992
rect 226668 223020 226674 223032
rect 280798 223020 280804 223032
rect 226668 222992 280804 223020
rect 226668 222980 226674 222992
rect 280798 222980 280804 222992
rect 280856 222980 280862 223032
rect 303614 222980 303620 223032
rect 303672 223020 303678 223032
rect 304350 223020 304356 223032
rect 303672 222992 304356 223020
rect 303672 222980 303678 222992
rect 304350 222980 304356 222992
rect 304408 222980 304414 223032
rect 155552 222856 224954 222884
rect 155552 222844 155558 222856
rect 245838 222844 245844 222896
rect 245896 222884 245902 222896
rect 246298 222884 246304 222896
rect 245896 222856 246304 222884
rect 245896 222844 245902 222856
rect 246298 222844 246304 222856
rect 246356 222884 246362 222896
rect 303614 222884 303620 222896
rect 246356 222856 303620 222884
rect 246356 222844 246362 222856
rect 303614 222844 303620 222856
rect 303672 222844 303678 222896
rect 254320 222176 254900 222204
rect 251266 222096 251272 222148
rect 251324 222136 251330 222148
rect 252094 222136 252100 222148
rect 251324 222108 252100 222136
rect 251324 222096 251330 222108
rect 252094 222096 252100 222108
rect 252152 222096 252158 222148
rect 252738 222096 252744 222148
rect 252796 222136 252802 222148
rect 253382 222136 253388 222148
rect 252796 222108 253388 222136
rect 252796 222096 252802 222108
rect 253382 222096 253388 222108
rect 253440 222096 253446 222148
rect 252646 222028 252652 222080
rect 252704 222068 252710 222080
rect 253566 222068 253572 222080
rect 252704 222040 253572 222068
rect 252704 222028 252710 222040
rect 253566 222028 253572 222040
rect 253624 222068 253630 222080
rect 254320 222068 254348 222176
rect 254394 222096 254400 222148
rect 254452 222136 254458 222148
rect 254762 222136 254768 222148
rect 254452 222108 254768 222136
rect 254452 222096 254458 222108
rect 254762 222096 254768 222108
rect 254820 222096 254826 222148
rect 254872 222136 254900 222176
rect 340966 222136 340972 222148
rect 254872 222108 340972 222136
rect 340966 222096 340972 222108
rect 341024 222096 341030 222148
rect 253624 222040 254348 222068
rect 254780 222068 254808 222096
rect 336734 222068 336740 222080
rect 254780 222040 336740 222068
rect 253624 222028 253630 222040
rect 336734 222028 336740 222040
rect 336792 222028 336798 222080
rect 254302 221960 254308 222012
rect 254360 222000 254366 222012
rect 254854 222000 254860 222012
rect 254360 221972 254860 222000
rect 254360 221960 254366 221972
rect 254854 221960 254860 221972
rect 254912 221960 254918 222012
rect 254946 221960 254952 222012
rect 255004 222000 255010 222012
rect 312906 222000 312912 222012
rect 255004 221972 312912 222000
rect 255004 221960 255010 221972
rect 312906 221960 312912 221972
rect 312964 221960 312970 222012
rect 254872 221932 254900 221960
rect 314286 221932 314292 221944
rect 254872 221904 314292 221932
rect 314286 221892 314292 221904
rect 314344 221892 314350 221944
rect 227070 221824 227076 221876
rect 227128 221864 227134 221876
rect 248506 221864 248512 221876
rect 227128 221836 248512 221864
rect 227128 221824 227134 221836
rect 248506 221824 248512 221836
rect 248564 221824 248570 221876
rect 252094 221824 252100 221876
rect 252152 221864 252158 221876
rect 254946 221864 254952 221876
rect 252152 221836 254952 221864
rect 252152 221824 252158 221836
rect 254946 221824 254952 221836
rect 255004 221824 255010 221876
rect 255038 221824 255044 221876
rect 255096 221864 255102 221876
rect 314102 221864 314108 221876
rect 255096 221836 314108 221864
rect 255096 221824 255102 221836
rect 314102 221824 314108 221836
rect 314160 221824 314166 221876
rect 230106 221756 230112 221808
rect 230164 221796 230170 221808
rect 254026 221796 254032 221808
rect 230164 221768 254032 221796
rect 230164 221756 230170 221768
rect 254026 221756 254032 221768
rect 254084 221796 254090 221808
rect 254210 221796 254216 221808
rect 254084 221768 254216 221796
rect 254084 221756 254090 221768
rect 254210 221756 254216 221768
rect 254268 221756 254274 221808
rect 254670 221756 254676 221808
rect 254728 221796 254734 221808
rect 314194 221796 314200 221808
rect 254728 221768 314200 221796
rect 254728 221756 254734 221768
rect 314194 221756 314200 221768
rect 314252 221756 314258 221808
rect 223114 221688 223120 221740
rect 223172 221728 223178 221740
rect 250254 221728 250260 221740
rect 223172 221700 250260 221728
rect 223172 221688 223178 221700
rect 250254 221688 250260 221700
rect 250312 221688 250318 221740
rect 253382 221688 253388 221740
rect 253440 221728 253446 221740
rect 307202 221728 307208 221740
rect 253440 221700 307208 221728
rect 253440 221688 253446 221700
rect 307202 221688 307208 221700
rect 307260 221688 307266 221740
rect 233694 221660 233700 221672
rect 219406 221632 233700 221660
rect 158254 221484 158260 221536
rect 158312 221524 158318 221536
rect 219406 221524 219434 221632
rect 233694 221620 233700 221632
rect 233752 221660 233758 221672
rect 283834 221660 283840 221672
rect 233752 221632 283840 221660
rect 233752 221620 233758 221632
rect 283834 221620 283840 221632
rect 283892 221620 283898 221672
rect 234982 221552 234988 221604
rect 235040 221592 235046 221604
rect 276382 221592 276388 221604
rect 235040 221564 276388 221592
rect 235040 221552 235046 221564
rect 276382 221552 276388 221564
rect 276440 221552 276446 221604
rect 158312 221496 219434 221524
rect 158312 221484 158318 221496
rect 242618 221484 242624 221536
rect 242676 221524 242682 221536
rect 272426 221524 272432 221536
rect 242676 221496 272432 221524
rect 242676 221484 242682 221496
rect 272426 221484 272432 221496
rect 272484 221524 272490 221536
rect 286318 221524 286324 221536
rect 272484 221496 286324 221524
rect 272484 221484 272490 221496
rect 286318 221484 286324 221496
rect 286376 221484 286382 221536
rect 160646 221416 160652 221468
rect 160704 221456 160710 221468
rect 238294 221456 238300 221468
rect 160704 221428 238300 221456
rect 160704 221416 160710 221428
rect 238294 221416 238300 221428
rect 238352 221416 238358 221468
rect 254026 221416 254032 221468
rect 254084 221456 254090 221468
rect 255038 221456 255044 221468
rect 254084 221428 255044 221456
rect 254084 221416 254090 221428
rect 255038 221416 255044 221428
rect 255096 221416 255102 221468
rect 260834 221416 260840 221468
rect 260892 221456 260898 221468
rect 294598 221456 294604 221468
rect 260892 221428 294604 221456
rect 260892 221416 260898 221428
rect 294598 221416 294604 221428
rect 294656 221456 294662 221468
rect 320818 221456 320824 221468
rect 294656 221428 320824 221456
rect 294656 221416 294662 221428
rect 320818 221416 320824 221428
rect 320876 221416 320882 221468
rect 248966 220736 248972 220788
rect 249024 220776 249030 220788
rect 249334 220776 249340 220788
rect 249024 220748 249340 220776
rect 249024 220736 249030 220748
rect 249334 220736 249340 220748
rect 249392 220736 249398 220788
rect 258718 220736 258724 220788
rect 258776 220776 258782 220788
rect 338114 220776 338120 220788
rect 258776 220748 338120 220776
rect 258776 220736 258782 220748
rect 338114 220736 338120 220748
rect 338172 220736 338178 220788
rect 247034 220668 247040 220720
rect 247092 220708 247098 220720
rect 247678 220708 247684 220720
rect 247092 220680 247684 220708
rect 247092 220668 247098 220680
rect 247678 220668 247684 220680
rect 247736 220708 247742 220720
rect 307110 220708 307116 220720
rect 247736 220680 307116 220708
rect 247736 220668 247742 220680
rect 307110 220668 307116 220680
rect 307168 220668 307174 220720
rect 226058 220600 226064 220652
rect 226116 220640 226122 220652
rect 279418 220640 279424 220652
rect 226116 220612 279424 220640
rect 226116 220600 226122 220612
rect 279418 220600 279424 220612
rect 279476 220600 279482 220652
rect 246666 220532 246672 220584
rect 246724 220572 246730 220584
rect 281166 220572 281172 220584
rect 246724 220544 281172 220572
rect 246724 220532 246730 220544
rect 281166 220532 281172 220544
rect 281224 220532 281230 220584
rect 225506 220260 225512 220312
rect 225564 220300 225570 220312
rect 226058 220300 226064 220312
rect 225564 220272 226064 220300
rect 225564 220260 225570 220272
rect 226058 220260 226064 220272
rect 226116 220260 226122 220312
rect 257614 220124 257620 220176
rect 257672 220164 257678 220176
rect 283742 220164 283748 220176
rect 257672 220136 283748 220164
rect 257672 220124 257678 220136
rect 283742 220124 283748 220136
rect 283800 220164 283806 220176
rect 318058 220164 318064 220176
rect 283800 220136 318064 220164
rect 283800 220124 283806 220136
rect 318058 220124 318064 220136
rect 318116 220124 318122 220176
rect 232774 220056 232780 220108
rect 232832 220096 232838 220108
rect 247034 220096 247040 220108
rect 232832 220068 247040 220096
rect 232832 220056 232838 220068
rect 247034 220056 247040 220068
rect 247092 220056 247098 220108
rect 249334 220056 249340 220108
rect 249392 220096 249398 220108
rect 309778 220096 309784 220108
rect 249392 220068 309784 220096
rect 249392 220056 249398 220068
rect 309778 220056 309784 220068
rect 309836 220056 309842 220108
rect 231854 219376 231860 219428
rect 231912 219416 231918 219428
rect 232314 219416 232320 219428
rect 231912 219388 232320 219416
rect 231912 219376 231918 219388
rect 232314 219376 232320 219388
rect 232372 219416 232378 219428
rect 292574 219416 292580 219428
rect 232372 219388 292580 219416
rect 232372 219376 232378 219388
rect 292574 219376 292580 219388
rect 292632 219376 292638 219428
rect 256418 219308 256424 219360
rect 256476 219348 256482 219360
rect 315298 219348 315304 219360
rect 256476 219320 315304 219348
rect 256476 219308 256482 219320
rect 315298 219308 315304 219320
rect 315356 219308 315362 219360
rect 246574 219240 246580 219292
rect 246632 219280 246638 219292
rect 304258 219280 304264 219292
rect 246632 219252 304264 219280
rect 246632 219240 246638 219252
rect 304258 219240 304264 219252
rect 304316 219240 304322 219292
rect 238386 219172 238392 219224
rect 238444 219212 238450 219224
rect 290458 219212 290464 219224
rect 238444 219184 290464 219212
rect 238444 219172 238450 219184
rect 290458 219172 290464 219184
rect 290516 219172 290522 219224
rect 255130 219104 255136 219156
rect 255188 219144 255194 219156
rect 294690 219144 294696 219156
rect 255188 219116 294696 219144
rect 255188 219104 255194 219116
rect 294690 219104 294696 219116
rect 294748 219104 294754 219156
rect 253750 219036 253756 219088
rect 253808 219076 253814 219088
rect 288066 219076 288072 219088
rect 253808 219048 288072 219076
rect 253808 219036 253814 219048
rect 288066 219036 288072 219048
rect 288124 219036 288130 219088
rect 253934 218900 253940 218952
rect 253992 218940 253998 218952
rect 254946 218940 254952 218952
rect 253992 218912 254952 218940
rect 253992 218900 253998 218912
rect 254946 218900 254952 218912
rect 255004 218900 255010 218952
rect 158162 218696 158168 218748
rect 158220 218736 158226 218748
rect 231854 218736 231860 218748
rect 158220 218708 231860 218736
rect 158220 218696 158226 218708
rect 231854 218696 231860 218708
rect 231912 218696 231918 218748
rect 254946 218696 254952 218748
rect 255004 218736 255010 218748
rect 313918 218736 313924 218748
rect 255004 218708 313924 218736
rect 255004 218696 255010 218708
rect 313918 218696 313924 218708
rect 313976 218696 313982 218748
rect 238110 218084 238116 218136
rect 238168 218124 238174 218136
rect 238386 218124 238392 218136
rect 238168 218096 238392 218124
rect 238168 218084 238174 218096
rect 238386 218084 238392 218096
rect 238444 218084 238450 218136
rect 246574 218084 246580 218136
rect 246632 218124 246638 218136
rect 246850 218124 246856 218136
rect 246632 218096 246856 218124
rect 246632 218084 246638 218096
rect 246850 218084 246856 218096
rect 246908 218084 246914 218136
rect 158070 218016 158076 218068
rect 158128 218056 158134 218068
rect 230566 218056 230572 218068
rect 158128 218028 230572 218056
rect 158128 218016 158134 218028
rect 230566 218016 230572 218028
rect 230624 218056 230630 218068
rect 231486 218056 231492 218068
rect 230624 218028 231492 218056
rect 230624 218016 230630 218028
rect 231486 218016 231492 218028
rect 231544 218016 231550 218068
rect 236914 218016 236920 218068
rect 236972 218056 236978 218068
rect 240962 218056 240968 218068
rect 236972 218028 240968 218056
rect 236972 218016 236978 218028
rect 240962 218016 240968 218028
rect 241020 218016 241026 218068
rect 204070 217948 204076 218000
rect 204128 217988 204134 218000
rect 223574 217988 223580 218000
rect 204128 217960 223580 217988
rect 204128 217948 204134 217960
rect 223574 217948 223580 217960
rect 223632 217948 223638 218000
rect 227162 217948 227168 218000
rect 227220 217988 227226 218000
rect 227714 217988 227720 218000
rect 227220 217960 227720 217988
rect 227220 217948 227226 217960
rect 227714 217948 227720 217960
rect 227772 217948 227778 218000
rect 187510 217336 187516 217388
rect 187568 217376 187574 217388
rect 215018 217376 215024 217388
rect 187568 217348 215024 217376
rect 187568 217336 187574 217348
rect 215018 217336 215024 217348
rect 215076 217336 215082 217388
rect 227714 217336 227720 217388
rect 227772 217376 227778 217388
rect 287882 217376 287888 217388
rect 227772 217348 287888 217376
rect 227772 217336 227778 217348
rect 287882 217336 287888 217348
rect 287940 217336 287946 217388
rect 151538 217268 151544 217320
rect 151596 217308 151602 217320
rect 204070 217308 204076 217320
rect 151596 217280 204076 217308
rect 151596 217268 151602 217280
rect 204070 217268 204076 217280
rect 204128 217268 204134 217320
rect 247126 217268 247132 217320
rect 247184 217308 247190 217320
rect 247678 217308 247684 217320
rect 247184 217280 247684 217308
rect 247184 217268 247190 217280
rect 247678 217268 247684 217280
rect 247736 217308 247742 217320
rect 308398 217308 308404 217320
rect 247736 217280 308404 217308
rect 247736 217268 247742 217280
rect 308398 217268 308404 217280
rect 308456 217268 308462 217320
rect 226794 216588 226800 216640
rect 226852 216628 226858 216640
rect 227162 216628 227168 216640
rect 226852 216600 227168 216628
rect 226852 216588 226858 216600
rect 227162 216588 227168 216600
rect 227220 216588 227226 216640
rect 228450 216588 228456 216640
rect 228508 216628 228514 216640
rect 228634 216628 228640 216640
rect 228508 216600 228640 216628
rect 228508 216588 228514 216600
rect 228634 216588 228640 216600
rect 228692 216588 228698 216640
rect 228726 216588 228732 216640
rect 228784 216628 228790 216640
rect 292850 216628 292856 216640
rect 228784 216600 292856 216628
rect 228784 216588 228790 216600
rect 292850 216588 292856 216600
rect 292908 216588 292914 216640
rect 227180 216560 227208 216588
rect 227180 216532 234614 216560
rect 227990 216452 227996 216504
rect 228048 216492 228054 216504
rect 228634 216492 228640 216504
rect 228048 216464 228640 216492
rect 228048 216452 228054 216464
rect 228634 216452 228640 216464
rect 228692 216452 228698 216504
rect 234586 216492 234614 216532
rect 246482 216520 246488 216572
rect 246540 216560 246546 216572
rect 247862 216560 247868 216572
rect 246540 216532 247868 216560
rect 246540 216520 246546 216532
rect 247862 216520 247868 216532
rect 247920 216560 247926 216572
rect 307110 216560 307116 216572
rect 247920 216532 307116 216560
rect 247920 216520 247926 216532
rect 307110 216520 307116 216532
rect 307168 216560 307174 216572
rect 307478 216560 307484 216572
rect 307168 216532 307484 216560
rect 307168 216520 307174 216532
rect 307478 216520 307484 216532
rect 307536 216520 307542 216572
rect 286410 216492 286416 216504
rect 234586 216464 286416 216492
rect 286410 216452 286416 216464
rect 286468 216452 286474 216504
rect 228450 216384 228456 216436
rect 228508 216424 228514 216436
rect 283650 216424 283656 216436
rect 228508 216396 283656 216424
rect 228508 216384 228514 216396
rect 283650 216384 283656 216396
rect 283708 216384 283714 216436
rect 228634 216316 228640 216368
rect 228692 216356 228698 216368
rect 283926 216356 283932 216368
rect 228692 216328 283932 216356
rect 228692 216316 228698 216328
rect 283926 216316 283932 216328
rect 283984 216316 283990 216368
rect 225322 216248 225328 216300
rect 225380 216288 225386 216300
rect 228726 216288 228732 216300
rect 225380 216260 228732 216288
rect 225380 216248 225386 216260
rect 228726 216248 228732 216260
rect 228784 216248 228790 216300
rect 230566 216248 230572 216300
rect 230624 216288 230630 216300
rect 282178 216288 282184 216300
rect 230624 216260 282184 216288
rect 230624 216248 230630 216260
rect 282178 216248 282184 216260
rect 282236 216248 282242 216300
rect 193398 216044 193404 216096
rect 193456 216084 193462 216096
rect 209038 216084 209044 216096
rect 193456 216056 209044 216084
rect 193456 216044 193462 216056
rect 209038 216044 209044 216056
rect 209096 216044 209102 216096
rect 180886 215976 180892 216028
rect 180944 216016 180950 216028
rect 217226 216016 217232 216028
rect 180944 215988 217232 216016
rect 180944 215976 180950 215988
rect 217226 215976 217232 215988
rect 217284 215976 217290 216028
rect 161658 215908 161664 215960
rect 161716 215948 161722 215960
rect 222286 215948 222292 215960
rect 161716 215920 222292 215948
rect 161716 215908 161722 215920
rect 222286 215908 222292 215920
rect 222344 215908 222350 215960
rect 205726 215228 205732 215280
rect 205784 215268 205790 215280
rect 206830 215268 206836 215280
rect 205784 215240 206836 215268
rect 205784 215228 205790 215240
rect 206830 215228 206836 215240
rect 206888 215268 206894 215280
rect 228174 215268 228180 215280
rect 206888 215240 228180 215268
rect 206888 215228 206894 215240
rect 228174 215228 228180 215240
rect 228232 215228 228238 215280
rect 205634 215160 205640 215212
rect 205692 215200 205698 215212
rect 206922 215200 206928 215212
rect 205692 215172 206928 215200
rect 205692 215160 205698 215172
rect 206922 215160 206928 215172
rect 206980 215200 206986 215212
rect 226886 215200 226892 215212
rect 206980 215172 226892 215200
rect 206980 215160 206986 215172
rect 226886 215160 226892 215172
rect 226944 215160 226950 215212
rect 183094 214752 183100 214804
rect 183152 214792 183158 214804
rect 214742 214792 214748 214804
rect 183152 214764 214748 214792
rect 183152 214752 183158 214764
rect 214742 214752 214748 214764
rect 214800 214752 214806 214804
rect 157978 214684 157984 214736
rect 158036 214724 158042 214736
rect 205634 214724 205640 214736
rect 158036 214696 205640 214724
rect 158036 214684 158042 214696
rect 205634 214684 205640 214696
rect 205692 214684 205698 214736
rect 156690 214616 156696 214668
rect 156748 214656 156754 214668
rect 205726 214656 205732 214668
rect 156748 214628 205732 214656
rect 156748 214616 156754 214628
rect 205726 214616 205732 214628
rect 205784 214616 205790 214668
rect 166994 214548 167000 214600
rect 167052 214588 167058 214600
rect 167730 214588 167736 214600
rect 167052 214560 167736 214588
rect 167052 214548 167058 214560
rect 167730 214548 167736 214560
rect 167788 214548 167794 214600
rect 168374 214548 168380 214600
rect 168432 214588 168438 214600
rect 168834 214588 168840 214600
rect 168432 214560 168840 214588
rect 168432 214548 168438 214560
rect 168834 214548 168840 214560
rect 168892 214548 168898 214600
rect 222194 214588 222200 214600
rect 169312 214560 222200 214588
rect 168466 214480 168472 214532
rect 168524 214520 168530 214532
rect 169202 214520 169208 214532
rect 168524 214492 169208 214520
rect 168524 214480 168530 214492
rect 169202 214480 169208 214492
rect 169260 214480 169266 214532
rect 161750 214412 161756 214464
rect 161808 214452 161814 214464
rect 169312 214452 169340 214560
rect 222194 214548 222200 214560
rect 222252 214548 222258 214600
rect 171134 214480 171140 214532
rect 171192 214520 171198 214532
rect 172146 214520 172152 214532
rect 171192 214492 172152 214520
rect 171192 214480 171198 214492
rect 172146 214480 172152 214492
rect 172204 214480 172210 214532
rect 172514 214480 172520 214532
rect 172572 214520 172578 214532
rect 173250 214520 173256 214532
rect 172572 214492 173256 214520
rect 172572 214480 172578 214492
rect 173250 214480 173256 214492
rect 173308 214480 173314 214532
rect 178034 214480 178040 214532
rect 178092 214520 178098 214532
rect 178770 214520 178776 214532
rect 178092 214492 178776 214520
rect 178092 214480 178098 214492
rect 178770 214480 178776 214492
rect 178828 214480 178834 214532
rect 180794 214480 180800 214532
rect 180852 214520 180858 214532
rect 181346 214520 181352 214532
rect 180852 214492 181352 214520
rect 180852 214480 180858 214492
rect 181346 214480 181352 214492
rect 181404 214480 181410 214532
rect 182266 214480 182272 214532
rect 182324 214520 182330 214532
rect 183186 214520 183192 214532
rect 182324 214492 183192 214520
rect 182324 214480 182330 214492
rect 183186 214480 183192 214492
rect 183244 214480 183250 214532
rect 183554 214480 183560 214532
rect 183612 214520 183618 214532
rect 184290 214520 184296 214532
rect 183612 214492 184296 214520
rect 183612 214480 183618 214492
rect 184290 214480 184296 214492
rect 184348 214480 184354 214532
rect 185026 214480 185032 214532
rect 185084 214520 185090 214532
rect 185394 214520 185400 214532
rect 185084 214492 185400 214520
rect 185084 214480 185090 214492
rect 185394 214480 185400 214492
rect 185452 214480 185458 214532
rect 186314 214480 186320 214532
rect 186372 214520 186378 214532
rect 186498 214520 186504 214532
rect 186372 214492 186504 214520
rect 186372 214480 186378 214492
rect 186498 214480 186504 214492
rect 186556 214480 186562 214532
rect 187694 214480 187700 214532
rect 187752 214520 187758 214532
rect 188338 214520 188344 214532
rect 187752 214492 188344 214520
rect 187752 214480 187758 214492
rect 188338 214480 188344 214492
rect 188396 214480 188402 214532
rect 189074 214480 189080 214532
rect 189132 214520 189138 214532
rect 189810 214520 189816 214532
rect 189132 214492 189816 214520
rect 189132 214480 189138 214492
rect 189810 214480 189816 214492
rect 189868 214480 189874 214532
rect 190454 214480 190460 214532
rect 190512 214520 190518 214532
rect 190914 214520 190920 214532
rect 190512 214492 190920 214520
rect 190512 214480 190518 214492
rect 190914 214480 190920 214492
rect 190972 214480 190978 214532
rect 191926 214480 191932 214532
rect 191984 214520 191990 214532
rect 192386 214520 192392 214532
rect 191984 214492 192392 214520
rect 191984 214480 191990 214492
rect 192386 214480 192392 214492
rect 192444 214480 192450 214532
rect 193306 214480 193312 214532
rect 193364 214520 193370 214532
rect 193858 214520 193864 214532
rect 193364 214492 193864 214520
rect 193364 214480 193370 214492
rect 193858 214480 193864 214492
rect 193916 214480 193922 214532
rect 194594 214480 194600 214532
rect 194652 214520 194658 214532
rect 195330 214520 195336 214532
rect 194652 214492 195336 214520
rect 194652 214480 194658 214492
rect 195330 214480 195336 214492
rect 195388 214480 195394 214532
rect 161808 214424 169340 214452
rect 161808 214412 161814 214424
rect 183646 214412 183652 214464
rect 183704 214452 183710 214464
rect 183922 214452 183928 214464
rect 183704 214424 183928 214452
rect 183704 214412 183710 214424
rect 183922 214412 183928 214424
rect 183980 214412 183986 214464
rect 184934 214412 184940 214464
rect 184992 214452 184998 214464
rect 185210 214452 185216 214464
rect 184992 214424 185216 214452
rect 184992 214412 184998 214424
rect 185210 214412 185216 214424
rect 185268 214412 185274 214464
rect 187786 214412 187792 214464
rect 187844 214452 187850 214464
rect 188706 214452 188712 214464
rect 187844 214424 188712 214452
rect 187844 214412 187850 214424
rect 188706 214412 188712 214424
rect 188764 214412 188770 214464
rect 186038 214208 186044 214260
rect 186096 214248 186102 214260
rect 189902 214248 189908 214260
rect 186096 214220 189908 214248
rect 186096 214208 186102 214220
rect 189902 214208 189908 214220
rect 189960 214208 189966 214260
rect 202874 214004 202880 214056
rect 202932 214044 202938 214056
rect 203150 214044 203156 214056
rect 202932 214016 203156 214044
rect 202932 214004 202938 214016
rect 203150 214004 203156 214016
rect 203208 214004 203214 214056
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 3200 213948 195284 213976
rect 3200 213936 3206 213948
rect 195256 213908 195284 213948
rect 200666 213908 200672 213920
rect 195256 213880 200672 213908
rect 200666 213868 200672 213880
rect 200724 213868 200730 213920
rect 202874 213868 202880 213920
rect 202932 213908 202938 213920
rect 204162 213908 204168 213920
rect 202932 213880 204168 213908
rect 202932 213868 202938 213880
rect 204162 213868 204168 213880
rect 204220 213908 204226 213920
rect 224402 213908 224408 213920
rect 204220 213880 224408 213908
rect 204220 213868 204226 213880
rect 224402 213868 224408 213880
rect 224460 213868 224466 213920
rect 177206 213392 177212 213444
rect 177264 213432 177270 213444
rect 209130 213432 209136 213444
rect 177264 213404 209136 213432
rect 177264 213392 177270 213404
rect 209130 213392 209136 213404
rect 209188 213392 209194 213444
rect 181990 213324 181996 213376
rect 182048 213364 182054 213376
rect 214650 213364 214656 213376
rect 182048 213336 214656 213364
rect 182048 213324 182054 213336
rect 214650 213324 214656 213336
rect 214708 213324 214714 213376
rect 153930 213256 153936 213308
rect 153988 213296 153994 213308
rect 202874 213296 202880 213308
rect 153988 213268 202880 213296
rect 153988 213256 153994 213268
rect 202874 213256 202880 213268
rect 202932 213256 202938 213308
rect 184842 213188 184848 213240
rect 184900 213228 184906 213240
rect 243998 213228 244004 213240
rect 184900 213200 244004 213228
rect 184900 213188 184906 213200
rect 243998 213188 244004 213200
rect 244056 213188 244062 213240
rect 249242 213188 249248 213240
rect 249300 213228 249306 213240
rect 335354 213228 335360 213240
rect 249300 213200 335360 213228
rect 249300 213188 249306 213200
rect 335354 213188 335360 213200
rect 335412 213228 335418 213240
rect 335998 213228 336004 213240
rect 335412 213200 336004 213228
rect 335412 213188 335418 213200
rect 335998 213188 336004 213200
rect 336056 213188 336062 213240
rect 194686 212712 194692 212764
rect 194744 212752 194750 212764
rect 194962 212752 194968 212764
rect 194744 212724 194968 212752
rect 194744 212712 194750 212724
rect 194962 212712 194968 212724
rect 195020 212712 195026 212764
rect 159266 212508 159272 212560
rect 159324 212548 159330 212560
rect 163498 212548 163504 212560
rect 159324 212520 163504 212548
rect 159324 212508 159330 212520
rect 163498 212508 163504 212520
rect 163556 212508 163562 212560
rect 165614 212440 165620 212492
rect 165672 212480 165678 212492
rect 170398 212480 170404 212492
rect 165672 212452 170404 212480
rect 165672 212440 165678 212452
rect 170398 212440 170404 212452
rect 170456 212440 170462 212492
rect 177574 212440 177580 212492
rect 177632 212480 177638 212492
rect 178678 212480 178684 212492
rect 177632 212452 178684 212480
rect 177632 212440 177638 212452
rect 178678 212440 178684 212452
rect 178736 212440 178742 212492
rect 187878 212440 187884 212492
rect 187936 212480 187942 212492
rect 189718 212480 189724 212492
rect 187936 212452 189724 212480
rect 187936 212440 187942 212452
rect 189718 212440 189724 212452
rect 189776 212440 189782 212492
rect 200574 212480 200580 212492
rect 195946 212452 200580 212480
rect 186314 212372 186320 212424
rect 186372 212412 186378 212424
rect 195946 212412 195974 212452
rect 200574 212440 200580 212452
rect 200632 212440 200638 212492
rect 200666 212440 200672 212492
rect 200724 212480 200730 212492
rect 219894 212480 219900 212492
rect 200724 212452 219900 212480
rect 200724 212440 200730 212452
rect 219894 212440 219900 212452
rect 219952 212440 219958 212492
rect 186372 212384 195974 212412
rect 186372 212372 186378 212384
rect 196342 212372 196348 212424
rect 196400 212412 196406 212424
rect 196400 212384 205634 212412
rect 196400 212372 196406 212384
rect 162026 212304 162032 212356
rect 162084 212344 162090 212356
rect 162762 212344 162768 212356
rect 162084 212316 162768 212344
rect 162084 212304 162090 212316
rect 162762 212304 162768 212316
rect 162820 212304 162826 212356
rect 200758 212344 200764 212356
rect 195946 212316 200764 212344
rect 179782 212236 179788 212288
rect 179840 212276 179846 212288
rect 189626 212276 189632 212288
rect 179840 212248 189632 212276
rect 179840 212236 179846 212248
rect 189626 212236 189632 212248
rect 189684 212236 189690 212288
rect 176470 212168 176476 212220
rect 176528 212208 176534 212220
rect 195946 212208 195974 212316
rect 200758 212304 200764 212316
rect 200816 212304 200822 212356
rect 202690 212344 202696 212356
rect 200868 212316 202696 212344
rect 197446 212236 197452 212288
rect 197504 212276 197510 212288
rect 198550 212276 198556 212288
rect 197504 212248 198556 212276
rect 197504 212236 197510 212248
rect 198550 212236 198556 212248
rect 198608 212236 198614 212288
rect 198918 212236 198924 212288
rect 198976 212276 198982 212288
rect 200022 212276 200028 212288
rect 198976 212248 200028 212276
rect 198976 212236 198982 212248
rect 200022 212236 200028 212248
rect 200080 212236 200086 212288
rect 200574 212236 200580 212288
rect 200632 212276 200638 212288
rect 200868 212276 200896 212316
rect 202690 212304 202696 212316
rect 202748 212344 202754 212356
rect 203702 212344 203708 212356
rect 202748 212316 203708 212344
rect 202748 212304 202754 212316
rect 203702 212304 203708 212316
rect 203760 212304 203766 212356
rect 205606 212344 205634 212384
rect 211798 212344 211804 212356
rect 205606 212316 211804 212344
rect 211798 212304 211804 212316
rect 211856 212304 211862 212356
rect 200632 212248 200896 212276
rect 200632 212236 200638 212248
rect 201218 212236 201224 212288
rect 201276 212276 201282 212288
rect 202598 212276 202604 212288
rect 201276 212248 202604 212276
rect 201276 212236 201282 212248
rect 202598 212236 202604 212248
rect 202656 212236 202662 212288
rect 202782 212236 202788 212288
rect 202840 212276 202846 212288
rect 203334 212276 203340 212288
rect 202840 212248 203340 212276
rect 202840 212236 202846 212248
rect 203334 212236 203340 212248
rect 203392 212236 203398 212288
rect 221918 212276 221924 212288
rect 205606 212248 221924 212276
rect 176528 212180 195974 212208
rect 176528 212168 176534 212180
rect 199286 212168 199292 212220
rect 199344 212208 199350 212220
rect 205606 212208 205634 212248
rect 221918 212236 221924 212248
rect 221976 212236 221982 212288
rect 199344 212180 205634 212208
rect 199344 212168 199350 212180
rect 175734 212100 175740 212152
rect 175792 212140 175798 212152
rect 180058 212140 180064 212152
rect 175792 212112 180064 212140
rect 175792 212100 175798 212112
rect 180058 212100 180064 212112
rect 180116 212100 180122 212152
rect 186958 212140 186964 212152
rect 180168 212112 186964 212140
rect 174630 212032 174636 212084
rect 174688 212072 174694 212084
rect 180168 212072 180196 212112
rect 186958 212100 186964 212112
rect 187016 212100 187022 212152
rect 189718 212100 189724 212152
rect 189776 212140 189782 212152
rect 221826 212140 221832 212152
rect 189776 212112 221832 212140
rect 189776 212100 189782 212112
rect 221826 212100 221832 212112
rect 221884 212100 221890 212152
rect 212258 212072 212264 212084
rect 174688 212044 180196 212072
rect 180260 212044 212264 212072
rect 174688 212032 174694 212044
rect 172054 211964 172060 212016
rect 172112 212004 172118 212016
rect 180260 212004 180288 212044
rect 212258 212032 212264 212044
rect 212316 212032 212322 212084
rect 172112 211976 180288 212004
rect 172112 211964 172118 211976
rect 180518 211964 180524 212016
rect 180576 212004 180582 212016
rect 221734 212004 221740 212016
rect 180576 211976 221740 212004
rect 180576 211964 180582 211976
rect 221734 211964 221740 211976
rect 221792 211964 221798 212016
rect 161934 211896 161940 211948
rect 161992 211936 161998 211948
rect 162670 211936 162676 211948
rect 161992 211908 162676 211936
rect 161992 211896 161998 211908
rect 162670 211896 162676 211908
rect 162728 211936 162734 211948
rect 166534 211936 166540 211948
rect 162728 211908 166540 211936
rect 162728 211896 162734 211908
rect 166534 211896 166540 211908
rect 166592 211896 166598 211948
rect 167638 211896 167644 211948
rect 167696 211936 167702 211948
rect 168282 211936 168288 211948
rect 167696 211908 168288 211936
rect 167696 211896 167702 211908
rect 168282 211896 168288 211908
rect 168340 211896 168346 211948
rect 175366 211896 175372 211948
rect 175424 211936 175430 211948
rect 217686 211936 217692 211948
rect 175424 211908 217692 211936
rect 175424 211896 175430 211908
rect 217686 211896 217692 211908
rect 217744 211896 217750 211948
rect 156598 211828 156604 211880
rect 156656 211868 156662 211880
rect 201494 211868 201500 211880
rect 156656 211840 201500 211868
rect 156656 211828 156662 211840
rect 201494 211828 201500 211840
rect 201552 211828 201558 211880
rect 11698 211760 11704 211812
rect 11756 211800 11762 211812
rect 201218 211800 201224 211812
rect 11756 211772 201224 211800
rect 11756 211760 11762 211772
rect 201218 211760 201224 211772
rect 201276 211760 201282 211812
rect 272242 211800 272248 211812
rect 205606 211772 272248 211800
rect 189074 211692 189080 211744
rect 189132 211732 189138 211744
rect 202782 211732 202788 211744
rect 189132 211704 202788 211732
rect 189132 211692 189138 211704
rect 202782 211692 202788 211704
rect 202840 211692 202846 211744
rect 95878 211488 95884 211540
rect 95936 211528 95942 211540
rect 204806 211528 204812 211540
rect 95936 211500 204812 211528
rect 95936 211488 95942 211500
rect 204806 211488 204812 211500
rect 204864 211528 204870 211540
rect 205606 211528 205634 211772
rect 272242 211760 272248 211772
rect 272300 211760 272306 211812
rect 204864 211500 205634 211528
rect 204864 211488 204870 211500
rect 170122 211420 170128 211472
rect 170180 211460 170186 211472
rect 187602 211460 187608 211472
rect 170180 211432 187608 211460
rect 170180 211420 170186 211432
rect 187602 211420 187608 211432
rect 187660 211420 187666 211472
rect 168742 211352 168748 211404
rect 168800 211392 168806 211404
rect 182542 211392 182548 211404
rect 168800 211364 182548 211392
rect 168800 211352 168806 211364
rect 182542 211352 182548 211364
rect 182600 211352 182606 211404
rect 168282 211284 168288 211336
rect 168340 211324 168346 211336
rect 189534 211324 189540 211336
rect 168340 211296 189540 211324
rect 168340 211284 168346 211296
rect 189534 211284 189540 211296
rect 189592 211284 189598 211336
rect 191742 211284 191748 211336
rect 191800 211324 191806 211336
rect 202138 211324 202144 211336
rect 191800 211296 202144 211324
rect 191800 211284 191806 211296
rect 202138 211284 202144 211296
rect 202196 211284 202202 211336
rect 183462 211216 183468 211268
rect 183520 211256 183526 211268
rect 206278 211256 206284 211268
rect 183520 211228 206284 211256
rect 183520 211216 183526 211228
rect 206278 211216 206284 211228
rect 206336 211216 206342 211268
rect 162026 211148 162032 211200
rect 162084 211188 162090 211200
rect 165430 211188 165436 211200
rect 162084 211160 165436 211188
rect 162084 211148 162090 211160
rect 165430 211148 165436 211160
rect 165488 211148 165494 211200
rect 195974 211012 195980 211064
rect 196032 211052 196038 211064
rect 196434 211052 196440 211064
rect 196032 211024 196440 211052
rect 196032 211012 196038 211024
rect 196434 211012 196440 211024
rect 196492 211012 196498 211064
rect 200114 210740 200120 210792
rect 200172 210780 200178 210792
rect 201126 210780 201132 210792
rect 200172 210752 201132 210780
rect 200172 210740 200178 210752
rect 201126 210740 201132 210752
rect 201184 210740 201190 210792
rect 174262 210672 174268 210724
rect 174320 210712 174326 210724
rect 212074 210712 212080 210724
rect 174320 210684 212080 210712
rect 174320 210672 174326 210684
rect 212074 210672 212080 210684
rect 212132 210672 212138 210724
rect 3418 210604 3424 210656
rect 3476 210644 3482 210656
rect 183462 210644 183468 210656
rect 3476 210616 183468 210644
rect 3476 210604 3482 210616
rect 183462 210604 183468 210616
rect 183520 210604 183526 210656
rect 3602 210536 3608 210588
rect 3660 210576 3666 210588
rect 186314 210576 186320 210588
rect 3660 210548 186320 210576
rect 3660 210536 3666 210548
rect 186314 210536 186320 210548
rect 186372 210536 186378 210588
rect 197354 210536 197360 210588
rect 197412 210576 197418 210588
rect 197630 210576 197636 210588
rect 197412 210548 197636 210576
rect 197412 210536 197418 210548
rect 197630 210536 197636 210548
rect 197688 210536 197694 210588
rect 3510 210468 3516 210520
rect 3568 210508 3574 210520
rect 189074 210508 189080 210520
rect 3568 210480 189080 210508
rect 3568 210468 3574 210480
rect 189074 210468 189080 210480
rect 189132 210468 189138 210520
rect 3694 210400 3700 210452
rect 3752 210440 3758 210452
rect 191742 210440 191748 210452
rect 3752 210412 191748 210440
rect 3752 210400 3758 210412
rect 191742 210400 191748 210412
rect 191800 210400 191806 210452
rect 193214 210264 193220 210316
rect 193272 210304 193278 210316
rect 194502 210304 194508 210316
rect 193272 210276 194508 210304
rect 193272 210264 193278 210276
rect 194502 210264 194508 210276
rect 194560 210264 194566 210316
rect 160554 209924 160560 209976
rect 160612 209964 160618 209976
rect 200942 209964 200948 209976
rect 160612 209936 200948 209964
rect 160612 209924 160618 209936
rect 200942 209924 200948 209936
rect 201000 209924 201006 209976
rect 202414 209964 202420 209976
rect 201972 209936 202420 209964
rect 159358 209856 159364 209908
rect 159416 209896 159422 209908
rect 201678 209896 201684 209908
rect 159416 209868 201684 209896
rect 159416 209856 159422 209868
rect 201678 209856 201684 209868
rect 201736 209896 201742 209908
rect 201972 209896 202000 209936
rect 202414 209924 202420 209936
rect 202472 209924 202478 209976
rect 201736 209868 202000 209896
rect 201736 209856 201742 209868
rect 155218 209788 155224 209840
rect 155276 209828 155282 209840
rect 204622 209828 204628 209840
rect 155276 209800 204628 209828
rect 155276 209788 155282 209800
rect 204622 209788 204628 209800
rect 204680 209788 204686 209840
rect 187694 209720 187700 209772
rect 187752 209760 187758 209772
rect 219250 209760 219256 209772
rect 187752 209732 219256 209760
rect 187752 209720 187758 209732
rect 219250 209720 219256 209732
rect 219308 209720 219314 209772
rect 199194 209584 199200 209636
rect 199252 209624 199258 209636
rect 199838 209624 199844 209636
rect 199252 209596 199844 209624
rect 199252 209584 199258 209596
rect 199838 209584 199844 209596
rect 199896 209584 199902 209636
rect 202874 209420 202880 209432
rect 195946 209392 202880 209420
rect 142798 209176 142804 209228
rect 142856 209216 142862 209228
rect 195946 209216 195974 209392
rect 202874 209380 202880 209392
rect 202932 209380 202938 209432
rect 203150 209380 203156 209432
rect 203208 209380 203214 209432
rect 203886 209380 203892 209432
rect 203944 209380 203950 209432
rect 204346 209420 204352 209432
rect 203996 209392 204352 209420
rect 203168 209352 203196 209380
rect 203904 209352 203932 209380
rect 142856 209188 195974 209216
rect 200960 209324 203932 209352
rect 142856 209176 142862 209188
rect 120718 209108 120724 209160
rect 120776 209148 120782 209160
rect 200960 209148 200988 209324
rect 203996 209284 204024 209392
rect 204346 209380 204352 209392
rect 204404 209420 204410 209432
rect 204990 209420 204996 209432
rect 204404 209392 204996 209420
rect 204404 209380 204410 209392
rect 204990 209380 204996 209392
rect 205048 209380 205054 209432
rect 120776 209120 200988 209148
rect 201880 209256 204024 209284
rect 120776 209108 120782 209120
rect 43438 209040 43444 209092
rect 43496 209080 43502 209092
rect 201880 209080 201908 209256
rect 43496 209052 201908 209080
rect 43496 209040 43502 209052
rect 219250 209040 219256 209092
rect 219308 209080 219314 209092
rect 579982 209080 579988 209092
rect 219308 209052 579988 209080
rect 219308 209040 219314 209052
rect 579982 209040 579988 209052
rect 580040 209040 580046 209092
rect 209130 207748 209136 207800
rect 209188 207788 209194 207800
rect 263226 207788 263232 207800
rect 209188 207760 263232 207788
rect 209188 207748 209194 207760
rect 263226 207748 263232 207760
rect 263284 207748 263290 207800
rect 209498 207680 209504 207732
rect 209556 207720 209562 207732
rect 264330 207720 264336 207732
rect 209556 207692 264336 207720
rect 209556 207680 209562 207692
rect 264330 207680 264336 207692
rect 264388 207680 264394 207732
rect 209038 207612 209044 207664
rect 209096 207652 209102 207664
rect 265802 207652 265808 207664
rect 209096 207624 265808 207652
rect 209096 207612 209102 207624
rect 265802 207612 265808 207624
rect 265860 207612 265866 207664
rect 210786 206252 210792 206304
rect 210844 206292 210850 206304
rect 263318 206292 263324 206304
rect 210844 206264 263324 206292
rect 210844 206252 210850 206264
rect 263318 206252 263324 206264
rect 263376 206252 263382 206304
rect 245654 204212 245660 204264
rect 245712 204252 245718 204264
rect 246758 204252 246764 204264
rect 245712 204224 246764 204252
rect 245712 204212 245718 204224
rect 246758 204212 246764 204224
rect 246816 204252 246822 204264
rect 327718 204252 327724 204264
rect 246816 204224 327724 204252
rect 246816 204212 246822 204224
rect 327718 204212 327724 204224
rect 327776 204212 327782 204264
rect 237006 203532 237012 203584
rect 237064 203572 237070 203584
rect 245654 203572 245660 203584
rect 237064 203544 245660 203572
rect 237064 203532 237070 203544
rect 245654 203532 245660 203544
rect 245712 203532 245718 203584
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 156598 202824 156604 202836
rect 3384 202796 156604 202824
rect 3384 202784 3390 202796
rect 156598 202784 156604 202796
rect 156656 202784 156662 202836
rect 209590 202104 209596 202156
rect 209648 202144 209654 202156
rect 259086 202144 259092 202156
rect 209648 202116 259092 202144
rect 209648 202104 209654 202116
rect 259086 202104 259092 202116
rect 259144 202104 259150 202156
rect 247034 200064 247040 200116
rect 247092 200104 247098 200116
rect 248138 200104 248144 200116
rect 247092 200076 248144 200104
rect 247092 200064 247098 200076
rect 248138 200064 248144 200076
rect 248196 200104 248202 200116
rect 342254 200104 342260 200116
rect 248196 200076 342260 200104
rect 248196 200064 248202 200076
rect 342254 200064 342260 200076
rect 342312 200064 342318 200116
rect 342254 199452 342260 199504
rect 342312 199492 342318 199504
rect 342898 199492 342904 199504
rect 342312 199464 342904 199492
rect 342312 199452 342318 199464
rect 342898 199452 342904 199464
rect 342956 199452 342962 199504
rect 235810 199384 235816 199436
rect 235868 199424 235874 199436
rect 247034 199424 247040 199436
rect 235868 199396 247040 199424
rect 235868 199384 235874 199396
rect 247034 199384 247040 199396
rect 247092 199384 247098 199436
rect 210878 196596 210884 196648
rect 210936 196636 210942 196648
rect 224126 196636 224132 196648
rect 210936 196608 224132 196636
rect 210936 196596 210942 196608
rect 224126 196596 224132 196608
rect 224184 196596 224190 196648
rect 338758 193128 338764 193180
rect 338816 193168 338822 193180
rect 580166 193168 580172 193180
rect 338816 193140 580172 193168
rect 338816 193128 338822 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 210970 192448 210976 192500
rect 211028 192488 211034 192500
rect 223390 192488 223396 192500
rect 211028 192460 223396 192488
rect 211028 192448 211034 192460
rect 223390 192448 223396 192460
rect 223448 192448 223454 192500
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 160554 189020 160560 189032
rect 3384 188992 160560 189020
rect 3384 188980 3390 188992
rect 160554 188980 160560 188992
rect 160612 188980 160618 189032
rect 211062 186940 211068 186992
rect 211120 186980 211126 186992
rect 224034 186980 224040 186992
rect 211120 186952 224040 186980
rect 211120 186940 211126 186952
rect 224034 186940 224040 186952
rect 224092 186940 224098 186992
rect 242710 186940 242716 186992
rect 242768 186980 242774 186992
rect 259454 186980 259460 186992
rect 242768 186952 259460 186980
rect 242768 186940 242774 186952
rect 259454 186940 259460 186952
rect 259512 186940 259518 186992
rect 257522 186328 257528 186380
rect 257580 186368 257586 186380
rect 257798 186368 257804 186380
rect 257580 186340 257804 186368
rect 257580 186328 257586 186340
rect 257798 186328 257804 186340
rect 257856 186368 257862 186380
rect 442994 186368 443000 186380
rect 257856 186340 443000 186368
rect 257856 186328 257862 186340
rect 442994 186328 443000 186340
rect 443052 186328 443058 186380
rect 230198 184152 230204 184204
rect 230256 184192 230262 184204
rect 250714 184192 250720 184204
rect 230256 184164 250720 184192
rect 230256 184152 230262 184164
rect 250714 184152 250720 184164
rect 250772 184192 250778 184204
rect 361574 184192 361580 184204
rect 250772 184164 361580 184192
rect 250772 184152 250778 184164
rect 361574 184152 361580 184164
rect 361632 184152 361638 184204
rect 209682 177284 209688 177336
rect 209740 177324 209746 177336
rect 266354 177324 266360 177336
rect 209740 177296 266360 177324
rect 209740 177284 209746 177296
rect 266354 177284 266360 177296
rect 266412 177284 266418 177336
rect 246574 176672 246580 176724
rect 246632 176712 246638 176724
rect 246850 176712 246856 176724
rect 246632 176684 246856 176712
rect 246632 176672 246638 176684
rect 246850 176672 246856 176684
rect 246908 176712 246914 176724
rect 304994 176712 305000 176724
rect 246908 176684 305000 176712
rect 246908 176672 246914 176684
rect 304994 176672 305000 176684
rect 305052 176672 305058 176724
rect 259362 175244 259368 175296
rect 259420 175284 259426 175296
rect 467834 175284 467840 175296
rect 259420 175256 467840 175284
rect 259420 175244 259426 175256
rect 467834 175244 467840 175256
rect 467892 175244 467898 175296
rect 256234 173952 256240 174004
rect 256292 173992 256298 174004
rect 256510 173992 256516 174004
rect 256292 173964 256516 173992
rect 256292 173952 256298 173964
rect 256510 173952 256516 173964
rect 256568 173992 256574 174004
rect 425054 173992 425060 174004
rect 256568 173964 425060 173992
rect 256568 173952 256574 173964
rect 425054 173952 425060 173964
rect 425112 173952 425118 174004
rect 256142 173884 256148 173936
rect 256200 173924 256206 173936
rect 432046 173924 432052 173936
rect 256200 173896 432052 173924
rect 256200 173884 256206 173896
rect 432046 173884 432052 173896
rect 432104 173884 432110 173936
rect 208946 173136 208952 173188
rect 209004 173176 209010 173188
rect 262306 173176 262312 173188
rect 209004 173148 262312 173176
rect 209004 173136 209010 173148
rect 262306 173136 262312 173148
rect 262364 173136 262370 173188
rect 245286 171096 245292 171148
rect 245344 171136 245350 171148
rect 298094 171136 298100 171148
rect 245344 171108 298100 171136
rect 245344 171096 245350 171108
rect 298094 171096 298100 171108
rect 298152 171096 298158 171148
rect 260374 169736 260380 169788
rect 260432 169776 260438 169788
rect 481726 169776 481732 169788
rect 260432 169748 481732 169776
rect 260432 169736 260438 169748
rect 481726 169736 481732 169748
rect 481784 169736 481790 169788
rect 245378 168376 245384 168428
rect 245436 168416 245442 168428
rect 287054 168416 287060 168428
rect 245436 168388 287060 168416
rect 245436 168376 245442 168388
rect 287054 168376 287060 168388
rect 287112 168376 287118 168428
rect 257614 167016 257620 167068
rect 257672 167056 257678 167068
rect 257982 167056 257988 167068
rect 257672 167028 257988 167056
rect 257672 167016 257678 167028
rect 257982 167016 257988 167028
rect 258040 167056 258046 167068
rect 447134 167056 447140 167068
rect 258040 167028 447140 167056
rect 258040 167016 258046 167028
rect 447134 167016 447140 167028
rect 447192 167016 447198 167068
rect 156966 166336 156972 166388
rect 157024 166336 157030 166388
rect 156874 166132 156880 166184
rect 156932 166172 156938 166184
rect 156984 166172 157012 166336
rect 156932 166144 157012 166172
rect 156932 166132 156938 166144
rect 253750 165588 253756 165640
rect 253808 165628 253814 165640
rect 397454 165628 397460 165640
rect 253808 165600 397460 165628
rect 253808 165588 253814 165600
rect 397454 165588 397460 165600
rect 397512 165588 397518 165640
rect 209774 164840 209780 164892
rect 209832 164880 209838 164892
rect 226058 164880 226064 164892
rect 209832 164852 226064 164880
rect 209832 164840 209838 164852
rect 226058 164840 226064 164852
rect 226116 164840 226122 164892
rect 161566 161508 161572 161560
rect 161624 161548 161630 161560
rect 162394 161548 162400 161560
rect 161624 161520 162400 161548
rect 161624 161508 161630 161520
rect 162394 161508 162400 161520
rect 162452 161508 162458 161560
rect 189046 161384 207612 161412
rect 189046 161344 189074 161384
rect 185228 161316 189074 161344
rect 185228 161072 185256 161316
rect 207474 161276 207480 161288
rect 179386 161044 185256 161072
rect 186976 161248 207480 161276
rect 179386 161004 179414 161044
rect 169772 160976 179414 161004
rect 158622 160624 158628 160676
rect 158680 160664 158686 160676
rect 161842 160664 161848 160676
rect 158680 160636 161848 160664
rect 158680 160624 158686 160636
rect 161842 160624 161848 160636
rect 161900 160624 161906 160676
rect 160002 160488 160008 160540
rect 160060 160528 160066 160540
rect 160060 160500 161474 160528
rect 160060 160488 160066 160500
rect 161446 160460 161474 160500
rect 162302 160460 162308 160472
rect 161446 160432 162308 160460
rect 162302 160420 162308 160432
rect 162360 160420 162366 160472
rect 156966 160352 156972 160404
rect 157024 160392 157030 160404
rect 157024 160364 163912 160392
rect 157024 160352 157030 160364
rect 159174 160284 159180 160336
rect 159232 160324 159238 160336
rect 159232 160296 161474 160324
rect 159232 160284 159238 160296
rect 161446 160120 161474 160296
rect 163884 160256 163912 160364
rect 163884 160228 167776 160256
rect 161446 160092 165844 160120
rect 161446 160024 165476 160052
rect 158070 159944 158076 159996
rect 158128 159984 158134 159996
rect 161446 159984 161474 160024
rect 158128 159956 161474 159984
rect 158128 159944 158134 159956
rect 152458 159876 152464 159928
rect 152516 159916 152522 159928
rect 152826 159916 152832 159928
rect 152516 159888 152832 159916
rect 152516 159876 152522 159888
rect 152826 159876 152832 159888
rect 152884 159876 152890 159928
rect 161750 159876 161756 159928
rect 161808 159916 161814 159928
rect 162578 159916 162584 159928
rect 161808 159888 162584 159916
rect 161808 159876 161814 159888
rect 162578 159876 162584 159888
rect 162636 159876 162642 159928
rect 162872 159888 163544 159916
rect 152844 159848 152872 159876
rect 159174 159848 159180 159860
rect 152844 159820 159180 159848
rect 159174 159808 159180 159820
rect 159232 159808 159238 159860
rect 161658 159808 161664 159860
rect 161716 159848 161722 159860
rect 162670 159848 162676 159860
rect 161716 159820 162676 159848
rect 161716 159808 161722 159820
rect 162670 159808 162676 159820
rect 162728 159808 162734 159860
rect 162486 159740 162492 159792
rect 162544 159780 162550 159792
rect 162872 159780 162900 159888
rect 163406 159848 163412 159860
rect 162544 159752 162900 159780
rect 163240 159820 163412 159848
rect 162544 159740 162550 159752
rect 161198 159672 161204 159724
rect 161256 159712 161262 159724
rect 161256 159684 162808 159712
rect 161256 159672 161262 159684
rect 156506 159604 156512 159656
rect 156564 159644 156570 159656
rect 156966 159644 156972 159656
rect 156564 159616 156972 159644
rect 156564 159604 156570 159616
rect 156966 159604 156972 159616
rect 157024 159604 157030 159656
rect 158346 159604 158352 159656
rect 158404 159644 158410 159656
rect 162670 159644 162676 159656
rect 158404 159616 162676 159644
rect 158404 159604 158410 159616
rect 162670 159604 162676 159616
rect 162728 159604 162734 159656
rect 162780 159644 162808 159684
rect 162946 159672 162952 159724
rect 163004 159712 163010 159724
rect 163240 159712 163268 159820
rect 163406 159808 163412 159820
rect 163464 159808 163470 159860
rect 163516 159780 163544 159888
rect 164786 159876 164792 159928
rect 164844 159876 164850 159928
rect 164804 159792 164832 159876
rect 165448 159792 165476 160024
rect 165816 159928 165844 160092
rect 167748 159928 167776 160228
rect 165798 159876 165804 159928
rect 165856 159876 165862 159928
rect 167730 159876 167736 159928
rect 167788 159876 167794 159928
rect 167822 159876 167828 159928
rect 167880 159916 167886 159928
rect 169772 159916 169800 160976
rect 186976 160936 187004 161248
rect 207474 161236 207480 161248
rect 207532 161236 207538 161288
rect 207584 161072 207612 161384
rect 207658 161100 207664 161152
rect 207716 161140 207722 161152
rect 249334 161140 249340 161152
rect 207716 161112 249340 161140
rect 207716 161100 207722 161112
rect 249334 161100 249340 161112
rect 249392 161100 249398 161152
rect 225598 161072 225604 161084
rect 207584 161044 225604 161072
rect 225598 161032 225604 161044
rect 225656 161032 225662 161084
rect 208394 160964 208400 161016
rect 208452 161004 208458 161016
rect 250622 161004 250628 161016
rect 208452 160976 250628 161004
rect 208452 160964 208458 160976
rect 250622 160964 250628 160976
rect 250680 160964 250686 161016
rect 173866 160908 187004 160936
rect 173866 160120 173894 160908
rect 207474 160896 207480 160948
rect 207532 160936 207538 160948
rect 229738 160936 229744 160948
rect 207532 160908 229744 160936
rect 207532 160896 207538 160908
rect 229738 160896 229744 160908
rect 229796 160896 229802 160948
rect 230750 160868 230756 160880
rect 190426 160840 230756 160868
rect 190426 160256 190454 160840
rect 230750 160828 230756 160840
rect 230808 160828 230814 160880
rect 249058 160800 249064 160812
rect 197740 160772 249064 160800
rect 197740 160392 197768 160772
rect 249058 160760 249064 160772
rect 249116 160760 249122 160812
rect 253198 160732 253204 160744
rect 205606 160704 253204 160732
rect 205606 160596 205634 160704
rect 253198 160692 253204 160704
rect 253256 160692 253262 160744
rect 170416 160092 173894 160120
rect 182146 160228 190454 160256
rect 193048 160364 197768 160392
rect 204226 160568 205634 160596
rect 170416 159928 170444 160092
rect 170600 160024 178448 160052
rect 167880 159888 169800 159916
rect 167880 159876 167886 159888
rect 170398 159876 170404 159928
rect 170456 159876 170462 159928
rect 170490 159848 170496 159860
rect 165632 159820 170496 159848
rect 165632 159792 165660 159820
rect 170490 159808 170496 159820
rect 170548 159808 170554 159860
rect 163682 159780 163688 159792
rect 163516 159752 163688 159780
rect 163682 159740 163688 159752
rect 163740 159740 163746 159792
rect 164786 159740 164792 159792
rect 164844 159740 164850 159792
rect 165430 159740 165436 159792
rect 165488 159740 165494 159792
rect 165614 159740 165620 159792
rect 165672 159740 165678 159792
rect 170600 159712 170628 160024
rect 170876 159956 175044 159984
rect 170876 159928 170904 159956
rect 170858 159876 170864 159928
rect 170916 159876 170922 159928
rect 170950 159876 170956 159928
rect 171008 159916 171014 159928
rect 171410 159916 171416 159928
rect 171008 159888 171088 159916
rect 171008 159876 171014 159888
rect 171060 159724 171088 159888
rect 171336 159888 171416 159916
rect 171336 159848 171364 159888
rect 171410 159876 171416 159888
rect 171468 159876 171474 159928
rect 171870 159876 171876 159928
rect 171928 159876 171934 159928
rect 174354 159876 174360 159928
rect 174412 159876 174418 159928
rect 174446 159876 174452 159928
rect 174504 159876 174510 159928
rect 174722 159916 174728 159928
rect 174648 159888 174728 159916
rect 171336 159820 171640 159848
rect 163004 159684 163268 159712
rect 163332 159684 170628 159712
rect 163004 159672 163010 159684
rect 163332 159644 163360 159684
rect 171042 159672 171048 159724
rect 171100 159672 171106 159724
rect 162780 159616 163360 159644
rect 165430 159604 165436 159656
rect 165488 159644 165494 159656
rect 165488 159616 170076 159644
rect 165488 159604 165494 159616
rect 153010 159536 153016 159588
rect 153068 159576 153074 159588
rect 169938 159576 169944 159588
rect 153068 159548 169944 159576
rect 153068 159536 153074 159548
rect 169938 159536 169944 159548
rect 169996 159536 170002 159588
rect 170048 159576 170076 159616
rect 170214 159604 170220 159656
rect 170272 159644 170278 159656
rect 171226 159644 171232 159656
rect 170272 159616 171232 159644
rect 170272 159604 170278 159616
rect 171226 159604 171232 159616
rect 171284 159604 171290 159656
rect 171318 159576 171324 159588
rect 170048 159548 171324 159576
rect 171318 159536 171324 159548
rect 171376 159536 171382 159588
rect 171612 159520 171640 159820
rect 171888 159780 171916 159876
rect 172698 159848 172704 159860
rect 172624 159820 172704 159848
rect 171962 159780 171968 159792
rect 171888 159752 171968 159780
rect 171962 159740 171968 159752
rect 172020 159740 172026 159792
rect 172624 159724 172652 159820
rect 172698 159808 172704 159820
rect 172756 159808 172762 159860
rect 173342 159808 173348 159860
rect 173400 159808 173406 159860
rect 172882 159740 172888 159792
rect 172940 159780 172946 159792
rect 173360 159780 173388 159808
rect 172940 159752 173388 159780
rect 172940 159740 172946 159752
rect 172606 159672 172612 159724
rect 172664 159672 172670 159724
rect 173342 159672 173348 159724
rect 173400 159712 173406 159724
rect 174372 159712 174400 159876
rect 174464 159724 174492 159876
rect 173400 159684 174400 159712
rect 173400 159672 173406 159684
rect 174446 159672 174452 159724
rect 174504 159672 174510 159724
rect 171870 159604 171876 159656
rect 171928 159644 171934 159656
rect 171928 159616 174308 159644
rect 171928 159604 171934 159616
rect 171778 159536 171784 159588
rect 171836 159576 171842 159588
rect 174280 159576 174308 159616
rect 174354 159604 174360 159656
rect 174412 159644 174418 159656
rect 174648 159644 174676 159888
rect 174722 159876 174728 159888
rect 174780 159876 174786 159928
rect 174814 159876 174820 159928
rect 174872 159876 174878 159928
rect 175016 159916 175044 159956
rect 178420 159916 178448 160024
rect 178494 159916 178500 159928
rect 175016 159888 175136 159916
rect 178420 159888 178500 159916
rect 174412 159616 174676 159644
rect 174832 159644 174860 159876
rect 175108 159848 175136 159888
rect 178494 159876 178500 159888
rect 178552 159876 178558 159928
rect 182146 159848 182174 160228
rect 193048 159984 193076 160364
rect 204226 160324 204254 160568
rect 191116 159956 193076 159984
rect 193600 160296 204254 160324
rect 175108 159820 182174 159848
rect 183094 159808 183100 159860
rect 183152 159808 183158 159860
rect 188982 159808 188988 159860
rect 189040 159848 189046 159860
rect 191116 159848 191144 159956
rect 191742 159876 191748 159928
rect 191800 159876 191806 159928
rect 193122 159876 193128 159928
rect 193180 159916 193186 159928
rect 193600 159916 193628 160296
rect 209130 160256 209136 160268
rect 203536 160228 209136 160256
rect 193180 159888 193628 159916
rect 193180 159876 193186 159888
rect 199286 159876 199292 159928
rect 199344 159876 199350 159928
rect 203426 159876 203432 159928
rect 203484 159916 203490 159928
rect 203536 159916 203564 160228
rect 209130 160216 209136 160228
rect 209188 160216 209194 160268
rect 208394 160188 208400 160200
rect 203484 159888 203564 159916
rect 203628 160160 208400 160188
rect 203484 159876 203490 159888
rect 189040 159820 191144 159848
rect 189040 159808 189046 159820
rect 182542 159740 182548 159792
rect 182600 159780 182606 159792
rect 183112 159780 183140 159808
rect 182600 159752 183140 159780
rect 182600 159740 182606 159752
rect 191098 159740 191104 159792
rect 191156 159780 191162 159792
rect 191760 159780 191788 159876
rect 199304 159848 199332 159876
rect 203628 159848 203656 160160
rect 208394 160148 208400 160160
rect 208452 160148 208458 160200
rect 208118 160120 208124 160132
rect 199304 159820 199424 159848
rect 199396 159792 199424 159820
rect 200224 159820 203656 159848
rect 205468 160092 208124 160120
rect 200224 159792 200252 159820
rect 191156 159752 191788 159780
rect 191156 159740 191162 159752
rect 199010 159740 199016 159792
rect 199068 159780 199074 159792
rect 199286 159780 199292 159792
rect 199068 159752 199292 159780
rect 199068 159740 199074 159752
rect 199286 159740 199292 159752
rect 199344 159740 199350 159792
rect 199378 159740 199384 159792
rect 199436 159740 199442 159792
rect 200206 159740 200212 159792
rect 200264 159740 200270 159792
rect 203242 159740 203248 159792
rect 203300 159780 203306 159792
rect 205468 159780 205496 160092
rect 208118 160080 208124 160092
rect 208176 160080 208182 160132
rect 280798 160080 280804 160132
rect 280856 160120 280862 160132
rect 300854 160120 300860 160132
rect 280856 160092 300860 160120
rect 280856 160080 280862 160092
rect 300854 160080 300860 160092
rect 300912 160080 300918 160132
rect 207842 160052 207848 160064
rect 203300 159752 205496 159780
rect 205606 160024 207848 160052
rect 203300 159740 203306 159752
rect 205606 159712 205634 160024
rect 207842 160012 207848 160024
rect 207900 160012 207906 160064
rect 207750 159984 207756 159996
rect 206204 159956 207756 159984
rect 206204 159928 206232 159956
rect 207750 159944 207756 159956
rect 207808 159944 207814 159996
rect 206186 159876 206192 159928
rect 206244 159876 206250 159928
rect 207014 159876 207020 159928
rect 207072 159916 207078 159928
rect 209682 159916 209688 159928
rect 207072 159888 209688 159916
rect 207072 159876 207078 159888
rect 209682 159876 209688 159888
rect 209740 159876 209746 159928
rect 207106 159808 207112 159860
rect 207164 159848 207170 159860
rect 207566 159848 207572 159860
rect 207164 159820 207572 159848
rect 207164 159808 207170 159820
rect 207566 159808 207572 159820
rect 207624 159808 207630 159860
rect 206278 159740 206284 159792
rect 206336 159780 206342 159792
rect 208302 159780 208308 159792
rect 206336 159752 208308 159780
rect 206336 159740 206342 159752
rect 208302 159740 208308 159752
rect 208360 159740 208366 159792
rect 175108 159684 205634 159712
rect 174906 159644 174912 159656
rect 174832 159616 174912 159644
rect 174412 159604 174418 159616
rect 174906 159604 174912 159616
rect 174964 159604 174970 159656
rect 175108 159576 175136 159684
rect 180058 159604 180064 159656
rect 180116 159644 180122 159656
rect 209314 159644 209320 159656
rect 180116 159616 209320 159644
rect 180116 159604 180122 159616
rect 209314 159604 209320 159616
rect 209372 159604 209378 159656
rect 171836 159548 174124 159576
rect 174280 159548 175136 159576
rect 171836 159536 171842 159548
rect 132494 159468 132500 159520
rect 132552 159508 132558 159520
rect 158622 159508 158628 159520
rect 132552 159480 158628 159508
rect 132552 159468 132558 159480
rect 158622 159468 158628 159480
rect 158680 159468 158686 159520
rect 161290 159468 161296 159520
rect 161348 159508 161354 159520
rect 170766 159508 170772 159520
rect 161348 159480 170772 159508
rect 161348 159468 161354 159480
rect 170766 159468 170772 159480
rect 170824 159468 170830 159520
rect 171594 159468 171600 159520
rect 171652 159468 171658 159520
rect 128354 159400 128360 159452
rect 128412 159440 128418 159452
rect 159266 159440 159272 159452
rect 128412 159412 159272 159440
rect 128412 159400 128418 159412
rect 159266 159400 159272 159412
rect 159324 159440 159330 159452
rect 171410 159440 171416 159452
rect 159324 159412 171416 159440
rect 159324 159400 159330 159412
rect 171410 159400 171416 159412
rect 171468 159400 171474 159452
rect 171686 159400 171692 159452
rect 171744 159440 171750 159452
rect 173986 159440 173992 159452
rect 171744 159412 173992 159440
rect 171744 159400 171750 159412
rect 173986 159400 173992 159412
rect 174044 159400 174050 159452
rect 174096 159440 174124 159548
rect 191006 159536 191012 159588
rect 191064 159576 191070 159588
rect 200206 159576 200212 159588
rect 191064 159548 200212 159576
rect 191064 159536 191070 159548
rect 200206 159536 200212 159548
rect 200264 159536 200270 159588
rect 204070 159536 204076 159588
rect 204128 159576 204134 159588
rect 207014 159576 207020 159588
rect 204128 159548 207020 159576
rect 204128 159536 204134 159548
rect 207014 159536 207020 159548
rect 207072 159536 207078 159588
rect 207474 159536 207480 159588
rect 207532 159576 207538 159588
rect 208210 159576 208216 159588
rect 207532 159548 208216 159576
rect 207532 159536 207538 159548
rect 208210 159536 208216 159548
rect 208268 159536 208274 159588
rect 174372 159480 182174 159508
rect 174372 159440 174400 159480
rect 174096 159412 174400 159440
rect 176102 159400 176108 159452
rect 176160 159440 176166 159452
rect 176286 159440 176292 159452
rect 176160 159412 176292 159440
rect 176160 159400 176166 159412
rect 176286 159400 176292 159412
rect 176344 159400 176350 159452
rect 182146 159440 182174 159480
rect 183738 159468 183744 159520
rect 183796 159508 183802 159520
rect 202690 159508 202696 159520
rect 183796 159480 202696 159508
rect 183796 159468 183802 159480
rect 202690 159468 202696 159480
rect 202748 159468 202754 159520
rect 205174 159468 205180 159520
rect 205232 159508 205238 159520
rect 205358 159508 205364 159520
rect 205232 159480 205364 159508
rect 205232 159468 205238 159480
rect 205358 159468 205364 159480
rect 205416 159468 205422 159520
rect 206186 159468 206192 159520
rect 206244 159508 206250 159520
rect 235626 159508 235632 159520
rect 206244 159480 235632 159508
rect 206244 159468 206250 159480
rect 235626 159468 235632 159480
rect 235684 159468 235690 159520
rect 207934 159440 207940 159452
rect 182146 159412 207940 159440
rect 207934 159400 207940 159412
rect 207992 159400 207998 159452
rect 96614 159332 96620 159384
rect 96672 159372 96678 159384
rect 152734 159372 152740 159384
rect 96672 159344 152740 159372
rect 96672 159332 96678 159344
rect 152734 159332 152740 159344
rect 152792 159372 152798 159384
rect 153010 159372 153016 159384
rect 152792 159344 153016 159372
rect 152792 159332 152798 159344
rect 153010 159332 153016 159344
rect 153068 159332 153074 159384
rect 162762 159332 162768 159384
rect 162820 159372 162826 159384
rect 163498 159372 163504 159384
rect 162820 159344 163504 159372
rect 162820 159332 162826 159344
rect 163498 159332 163504 159344
rect 163556 159372 163562 159384
rect 171870 159372 171876 159384
rect 163556 159344 171876 159372
rect 163556 159332 163562 159344
rect 171870 159332 171876 159344
rect 171928 159332 171934 159384
rect 174722 159332 174728 159384
rect 174780 159372 174786 159384
rect 175090 159372 175096 159384
rect 174780 159344 175096 159372
rect 174780 159332 174786 159344
rect 175090 159332 175096 159344
rect 175148 159332 175154 159384
rect 187694 159332 187700 159384
rect 187752 159372 187758 159384
rect 228358 159372 228364 159384
rect 187752 159344 228364 159372
rect 187752 159332 187758 159344
rect 228358 159332 228364 159344
rect 228416 159332 228422 159384
rect 153930 159264 153936 159316
rect 153988 159304 153994 159316
rect 164234 159304 164240 159316
rect 153988 159276 164240 159304
rect 153988 159264 153994 159276
rect 164234 159264 164240 159276
rect 164292 159304 164298 159316
rect 164786 159304 164792 159316
rect 164292 159276 164792 159304
rect 164292 159264 164298 159276
rect 164786 159264 164792 159276
rect 164844 159264 164850 159316
rect 165798 159264 165804 159316
rect 165856 159304 165862 159316
rect 166074 159304 166080 159316
rect 165856 159276 166080 159304
rect 165856 159264 165862 159276
rect 166074 159264 166080 159276
rect 166132 159264 166138 159316
rect 166810 159264 166816 159316
rect 166868 159304 166874 159316
rect 170398 159304 170404 159316
rect 166868 159276 170404 159304
rect 166868 159264 166874 159276
rect 170398 159264 170404 159276
rect 170456 159264 170462 159316
rect 170582 159264 170588 159316
rect 170640 159304 170646 159316
rect 170950 159304 170956 159316
rect 170640 159276 170956 159304
rect 170640 159264 170646 159276
rect 170950 159264 170956 159276
rect 171008 159264 171014 159316
rect 171226 159264 171232 159316
rect 171284 159304 171290 159316
rect 175274 159304 175280 159316
rect 171284 159276 175280 159304
rect 171284 159264 171290 159276
rect 175274 159264 175280 159276
rect 175332 159264 175338 159316
rect 176102 159264 176108 159316
rect 176160 159304 176166 159316
rect 210142 159304 210148 159316
rect 176160 159276 210148 159304
rect 176160 159264 176166 159276
rect 210142 159264 210148 159276
rect 210200 159264 210206 159316
rect 154114 159196 154120 159248
rect 154172 159236 154178 159248
rect 164142 159236 164148 159248
rect 154172 159208 164148 159236
rect 154172 159196 154178 159208
rect 164142 159196 164148 159208
rect 164200 159196 164206 159248
rect 166166 159196 166172 159248
rect 166224 159236 166230 159248
rect 222378 159236 222384 159248
rect 166224 159208 222384 159236
rect 166224 159196 166230 159208
rect 222378 159196 222384 159208
rect 222436 159196 222442 159248
rect 162670 159128 162676 159180
rect 162728 159168 162734 159180
rect 164786 159168 164792 159180
rect 162728 159140 164792 159168
rect 162728 159128 162734 159140
rect 164786 159128 164792 159140
rect 164844 159128 164850 159180
rect 165890 159128 165896 159180
rect 165948 159168 165954 159180
rect 166074 159168 166080 159180
rect 165948 159140 166080 159168
rect 165948 159128 165954 159140
rect 166074 159128 166080 159140
rect 166132 159128 166138 159180
rect 223298 159168 223304 159180
rect 166966 159140 223304 159168
rect 161842 159060 161848 159112
rect 161900 159100 161906 159112
rect 162946 159100 162952 159112
rect 161900 159072 162952 159100
rect 161900 159060 161906 159072
rect 162946 159060 162952 159072
rect 163004 159060 163010 159112
rect 163130 159060 163136 159112
rect 163188 159100 163194 159112
rect 163682 159100 163688 159112
rect 163188 159072 163688 159100
rect 163188 159060 163194 159072
rect 163682 159060 163688 159072
rect 163740 159060 163746 159112
rect 164418 159060 164424 159112
rect 164476 159100 164482 159112
rect 164694 159100 164700 159112
rect 164476 159072 164700 159100
rect 164476 159060 164482 159072
rect 164694 159060 164700 159072
rect 164752 159100 164758 159112
rect 166966 159100 166994 159140
rect 223298 159128 223304 159140
rect 223356 159128 223362 159180
rect 164752 159072 166994 159100
rect 164752 159060 164758 159072
rect 169754 159060 169760 159112
rect 169812 159100 169818 159112
rect 170582 159100 170588 159112
rect 169812 159072 170588 159100
rect 169812 159060 169818 159072
rect 170582 159060 170588 159072
rect 170640 159100 170646 159112
rect 170640 159072 176654 159100
rect 170640 159060 170646 159072
rect 155586 158992 155592 159044
rect 155644 159032 155650 159044
rect 155644 159004 157334 159032
rect 155644 158992 155650 159004
rect 157306 158964 157334 159004
rect 162210 158992 162216 159044
rect 162268 159032 162274 159044
rect 171318 159032 171324 159044
rect 162268 159004 171324 159032
rect 162268 158992 162274 159004
rect 171318 158992 171324 159004
rect 171376 158992 171382 159044
rect 171410 158992 171416 159044
rect 171468 159032 171474 159044
rect 172422 159032 172428 159044
rect 171468 159004 172428 159032
rect 171468 158992 171474 159004
rect 172422 158992 172428 159004
rect 172480 158992 172486 159044
rect 174722 158992 174728 159044
rect 174780 159032 174786 159044
rect 174780 159004 174952 159032
rect 174780 158992 174786 159004
rect 165338 158964 165344 158976
rect 157306 158936 165344 158964
rect 165338 158924 165344 158936
rect 165396 158924 165402 158976
rect 172606 158964 172612 158976
rect 168484 158936 172612 158964
rect 162854 158856 162860 158908
rect 162912 158896 162918 158908
rect 163130 158896 163136 158908
rect 162912 158868 163136 158896
rect 162912 158856 162918 158868
rect 163130 158856 163136 158868
rect 163188 158856 163194 158908
rect 163222 158856 163228 158908
rect 163280 158896 163286 158908
rect 163406 158896 163412 158908
rect 163280 158868 163412 158896
rect 163280 158856 163286 158868
rect 163406 158856 163412 158868
rect 163464 158856 163470 158908
rect 168484 158896 168512 158936
rect 172606 158924 172612 158936
rect 172664 158924 172670 158976
rect 174924 158964 174952 159004
rect 175274 158992 175280 159044
rect 175332 159032 175338 159044
rect 175642 159032 175648 159044
rect 175332 159004 175648 159032
rect 175332 158992 175338 159004
rect 175642 158992 175648 159004
rect 175700 158992 175706 159044
rect 176626 159032 176654 159072
rect 185118 159060 185124 159112
rect 185176 159100 185182 159112
rect 245010 159100 245016 159112
rect 185176 159072 245016 159100
rect 185176 159060 185182 159072
rect 245010 159060 245016 159072
rect 245068 159060 245074 159112
rect 229186 159032 229192 159044
rect 176626 159004 229192 159032
rect 229186 158992 229192 159004
rect 229244 158992 229250 159044
rect 180058 158964 180064 158976
rect 174924 158936 180064 158964
rect 180058 158924 180064 158936
rect 180116 158924 180122 158976
rect 190914 158924 190920 158976
rect 190972 158964 190978 158976
rect 200206 158964 200212 158976
rect 190972 158936 200212 158964
rect 190972 158924 190978 158936
rect 200206 158924 200212 158936
rect 200264 158924 200270 158976
rect 253658 158964 253664 158976
rect 200776 158936 253664 158964
rect 163516 158868 168512 158896
rect 158622 158788 158628 158840
rect 158680 158828 158686 158840
rect 163516 158828 163544 158868
rect 170766 158856 170772 158908
rect 170824 158896 170830 158908
rect 176654 158896 176660 158908
rect 170824 158868 176660 158896
rect 170824 158856 170830 158868
rect 176654 158856 176660 158868
rect 176712 158856 176718 158908
rect 192938 158856 192944 158908
rect 192996 158896 193002 158908
rect 192996 158868 193168 158896
rect 192996 158856 193002 158868
rect 193140 158840 193168 158868
rect 193306 158856 193312 158908
rect 193364 158896 193370 158908
rect 200776 158896 200804 158936
rect 253658 158924 253664 158936
rect 253716 158924 253722 158976
rect 193364 158868 200804 158896
rect 193364 158856 193370 158868
rect 200850 158856 200856 158908
rect 200908 158896 200914 158908
rect 269114 158896 269120 158908
rect 200908 158868 269120 158896
rect 200908 158856 200914 158868
rect 269114 158856 269120 158868
rect 269172 158896 269178 158908
rect 270218 158896 270224 158908
rect 269172 158868 270224 158896
rect 269172 158856 269178 158868
rect 270218 158856 270224 158868
rect 270276 158856 270282 158908
rect 158680 158800 163544 158828
rect 158680 158788 158686 158800
rect 164786 158788 164792 158840
rect 164844 158828 164850 158840
rect 171226 158828 171232 158840
rect 164844 158800 171232 158828
rect 164844 158788 164850 158800
rect 171226 158788 171232 158800
rect 171284 158788 171290 158840
rect 171318 158788 171324 158840
rect 171376 158828 171382 158840
rect 176378 158828 176384 158840
rect 171376 158800 176384 158828
rect 171376 158788 171382 158800
rect 162854 158720 162860 158772
rect 162912 158760 162918 158772
rect 164050 158760 164056 158772
rect 162912 158732 164056 158760
rect 162912 158720 162918 158732
rect 164050 158720 164056 158732
rect 164108 158720 164114 158772
rect 167362 158720 167368 158772
rect 167420 158760 167426 158772
rect 167822 158760 167828 158772
rect 167420 158732 167828 158760
rect 167420 158720 167426 158732
rect 167822 158720 167828 158732
rect 167880 158720 167886 158772
rect 168742 158720 168748 158772
rect 168800 158760 168806 158772
rect 174722 158760 174728 158772
rect 168800 158732 174728 158760
rect 168800 158720 168806 158732
rect 174722 158720 174728 158732
rect 174780 158720 174786 158772
rect 158346 158652 158352 158704
rect 158404 158692 158410 158704
rect 164694 158692 164700 158704
rect 158404 158664 164700 158692
rect 158404 158652 158410 158664
rect 164694 158652 164700 158664
rect 164752 158652 164758 158704
rect 167086 158652 167092 158704
rect 167144 158692 167150 158704
rect 171686 158692 171692 158704
rect 167144 158664 171692 158692
rect 167144 158652 167150 158664
rect 171686 158652 171692 158664
rect 171744 158652 171750 158704
rect 168558 158624 168564 158636
rect 162964 158596 168564 158624
rect 156690 158516 156696 158568
rect 156748 158556 156754 158568
rect 162964 158556 162992 158596
rect 168558 158584 168564 158596
rect 168616 158584 168622 158636
rect 171318 158584 171324 158636
rect 171376 158624 171382 158636
rect 171594 158624 171600 158636
rect 171376 158596 171600 158624
rect 171376 158584 171382 158596
rect 171594 158584 171600 158596
rect 171652 158584 171658 158636
rect 171962 158584 171968 158636
rect 172020 158624 172026 158636
rect 172422 158624 172428 158636
rect 172020 158596 172428 158624
rect 172020 158584 172026 158596
rect 172422 158584 172428 158596
rect 172480 158584 172486 158636
rect 174078 158584 174084 158636
rect 174136 158624 174142 158636
rect 174814 158624 174820 158636
rect 174136 158596 174820 158624
rect 174136 158584 174142 158596
rect 174814 158584 174820 158596
rect 174872 158584 174878 158636
rect 174998 158584 175004 158636
rect 175056 158584 175062 158636
rect 156748 158528 162992 158556
rect 156748 158516 156754 158528
rect 163130 158516 163136 158568
rect 163188 158556 163194 158568
rect 163590 158556 163596 158568
rect 163188 158528 163596 158556
rect 163188 158516 163194 158528
rect 163590 158516 163596 158528
rect 163648 158516 163654 158568
rect 165154 158556 165160 158568
rect 164436 158528 165160 158556
rect 161014 158448 161020 158500
rect 161072 158488 161078 158500
rect 163682 158488 163688 158500
rect 161072 158460 163688 158488
rect 161072 158448 161078 158460
rect 163682 158448 163688 158460
rect 163740 158448 163746 158500
rect 156598 158380 156604 158432
rect 156656 158420 156662 158432
rect 163866 158420 163872 158432
rect 156656 158392 163872 158420
rect 156656 158380 156662 158392
rect 163866 158380 163872 158392
rect 163924 158380 163930 158432
rect 151078 158312 151084 158364
rect 151136 158352 151142 158364
rect 164436 158352 164464 158528
rect 165154 158516 165160 158528
rect 165212 158516 165218 158568
rect 166074 158516 166080 158568
rect 166132 158556 166138 158568
rect 175016 158556 175044 158584
rect 166132 158528 175044 158556
rect 175384 158556 175412 158800
rect 176378 158788 176384 158800
rect 176436 158788 176442 158840
rect 193122 158788 193128 158840
rect 193180 158788 193186 158840
rect 199378 158788 199384 158840
rect 199436 158828 199442 158840
rect 272334 158828 272340 158840
rect 199436 158800 272340 158828
rect 199436 158788 199442 158800
rect 272334 158788 272340 158800
rect 272392 158788 272398 158840
rect 175734 158720 175740 158772
rect 175792 158760 175798 158772
rect 176010 158760 176016 158772
rect 175792 158732 176016 158760
rect 175792 158720 175798 158732
rect 176010 158720 176016 158732
rect 176068 158720 176074 158772
rect 185854 158720 185860 158772
rect 185912 158760 185918 158772
rect 280798 158760 280804 158772
rect 185912 158732 192892 158760
rect 185912 158720 185918 158732
rect 175458 158652 175464 158704
rect 175516 158692 175522 158704
rect 176378 158692 176384 158704
rect 175516 158664 176384 158692
rect 175516 158652 175522 158664
rect 176378 158652 176384 158664
rect 176436 158652 176442 158704
rect 182726 158652 182732 158704
rect 182784 158692 182790 158704
rect 187418 158692 187424 158704
rect 182784 158664 187424 158692
rect 182784 158652 182790 158664
rect 187418 158652 187424 158664
rect 187476 158652 187482 158704
rect 190454 158652 190460 158704
rect 190512 158692 190518 158704
rect 190914 158692 190920 158704
rect 190512 158664 190920 158692
rect 190512 158652 190518 158664
rect 190914 158652 190920 158664
rect 190972 158652 190978 158704
rect 191006 158652 191012 158704
rect 191064 158692 191070 158704
rect 191558 158692 191564 158704
rect 191064 158664 191564 158692
rect 191064 158652 191070 158664
rect 191558 158652 191564 158664
rect 191616 158652 191622 158704
rect 192386 158652 192392 158704
rect 192444 158692 192450 158704
rect 192662 158692 192668 158704
rect 192444 158664 192668 158692
rect 192444 158652 192450 158664
rect 192662 158652 192668 158664
rect 192720 158652 192726 158704
rect 192864 158692 192892 158732
rect 193048 158732 203380 158760
rect 193048 158692 193076 158732
rect 192864 158664 193076 158692
rect 194594 158652 194600 158704
rect 194652 158692 194658 158704
rect 194652 158664 200620 158692
rect 194652 158652 194658 158664
rect 187142 158584 187148 158636
rect 187200 158624 187206 158636
rect 187200 158596 191604 158624
rect 187200 158584 187206 158596
rect 175458 158556 175464 158568
rect 175384 158528 175464 158556
rect 166132 158516 166138 158528
rect 175458 158516 175464 158528
rect 175516 158516 175522 158568
rect 178494 158516 178500 158568
rect 178552 158556 178558 158568
rect 182726 158556 182732 158568
rect 178552 158528 182732 158556
rect 178552 158516 178558 158528
rect 182726 158516 182732 158528
rect 182784 158516 182790 158568
rect 186866 158516 186872 158568
rect 186924 158556 186930 158568
rect 188522 158556 188528 158568
rect 186924 158528 188528 158556
rect 186924 158516 186930 158528
rect 188522 158516 188528 158528
rect 188580 158516 188586 158568
rect 168006 158448 168012 158500
rect 168064 158488 168070 158500
rect 168282 158488 168288 158500
rect 168064 158460 168288 158488
rect 168064 158448 168070 158460
rect 168282 158448 168288 158460
rect 168340 158448 168346 158500
rect 168558 158448 168564 158500
rect 168616 158488 168622 158500
rect 170214 158488 170220 158500
rect 168616 158460 170220 158488
rect 168616 158448 168622 158460
rect 170214 158448 170220 158460
rect 170272 158448 170278 158500
rect 182450 158448 182456 158500
rect 182508 158488 182514 158500
rect 189718 158488 189724 158500
rect 182508 158460 189724 158488
rect 182508 158448 182514 158460
rect 189718 158448 189724 158460
rect 189776 158448 189782 158500
rect 191576 158488 191604 158596
rect 192018 158584 192024 158636
rect 192076 158624 192082 158636
rect 193674 158624 193680 158636
rect 192076 158596 193680 158624
rect 192076 158584 192082 158596
rect 193674 158584 193680 158596
rect 193732 158584 193738 158636
rect 194870 158584 194876 158636
rect 194928 158624 194934 158636
rect 195698 158624 195704 158636
rect 194928 158596 195704 158624
rect 194928 158584 194934 158596
rect 195698 158584 195704 158596
rect 195756 158584 195762 158636
rect 198918 158584 198924 158636
rect 198976 158624 198982 158636
rect 200022 158624 200028 158636
rect 198976 158596 200028 158624
rect 198976 158584 198982 158596
rect 200022 158584 200028 158596
rect 200080 158584 200086 158636
rect 200592 158624 200620 158664
rect 200666 158652 200672 158704
rect 200724 158692 200730 158704
rect 201218 158692 201224 158704
rect 200724 158664 201224 158692
rect 200724 158652 200730 158664
rect 201218 158652 201224 158664
rect 201276 158652 201282 158704
rect 203352 158692 203380 158732
rect 203536 158732 280804 158760
rect 203536 158692 203564 158732
rect 280798 158720 280804 158732
rect 280856 158720 280862 158772
rect 203352 158664 203564 158692
rect 204254 158652 204260 158704
rect 204312 158692 204318 158704
rect 207658 158692 207664 158704
rect 204312 158664 207664 158692
rect 204312 158652 204318 158664
rect 207658 158652 207664 158664
rect 207716 158652 207722 158704
rect 204070 158624 204076 158636
rect 200592 158596 204076 158624
rect 204070 158584 204076 158596
rect 204128 158584 204134 158636
rect 234522 158624 234528 158636
rect 205376 158596 234528 158624
rect 193766 158516 193772 158568
rect 193824 158556 193830 158568
rect 195238 158556 195244 158568
rect 193824 158528 195244 158556
rect 193824 158516 193830 158528
rect 195238 158516 195244 158528
rect 195296 158516 195302 158568
rect 197354 158516 197360 158568
rect 197412 158556 197418 158568
rect 200850 158556 200856 158568
rect 197412 158528 200856 158556
rect 197412 158516 197418 158528
rect 200850 158516 200856 158528
rect 200908 158516 200914 158568
rect 202138 158516 202144 158568
rect 202196 158556 202202 158568
rect 202598 158556 202604 158568
rect 202196 158528 202604 158556
rect 202196 158516 202202 158528
rect 202598 158516 202604 158528
rect 202656 158516 202662 158568
rect 202690 158516 202696 158568
rect 202748 158556 202754 158568
rect 203334 158556 203340 158568
rect 202748 158528 203340 158556
rect 202748 158516 202754 158528
rect 203334 158516 203340 158528
rect 203392 158516 203398 158568
rect 205376 158556 205404 158596
rect 234522 158584 234528 158596
rect 234580 158584 234586 158636
rect 205284 158528 205404 158556
rect 199654 158488 199660 158500
rect 191576 158460 199660 158488
rect 199654 158448 199660 158460
rect 199712 158448 199718 158500
rect 201770 158448 201776 158500
rect 201828 158488 201834 158500
rect 205284 158488 205312 158528
rect 207382 158516 207388 158568
rect 207440 158556 207446 158568
rect 208302 158556 208308 158568
rect 207440 158528 208308 158556
rect 207440 158516 207446 158528
rect 208302 158516 208308 158528
rect 208360 158516 208366 158568
rect 201828 158460 205312 158488
rect 201828 158448 201834 158460
rect 165982 158380 165988 158432
rect 166040 158420 166046 158432
rect 208854 158420 208860 158432
rect 166040 158392 205312 158420
rect 166040 158380 166046 158392
rect 151136 158324 164464 158352
rect 151136 158312 151142 158324
rect 164878 158312 164884 158364
rect 164936 158352 164942 158364
rect 165062 158352 165068 158364
rect 164936 158324 165068 158352
rect 164936 158312 164942 158324
rect 165062 158312 165068 158324
rect 165120 158312 165126 158364
rect 168742 158312 168748 158364
rect 168800 158352 168806 158364
rect 169294 158352 169300 158364
rect 168800 158324 169300 158352
rect 168800 158312 168806 158324
rect 169294 158312 169300 158324
rect 169352 158312 169358 158364
rect 171042 158312 171048 158364
rect 171100 158352 171106 158364
rect 205284 158352 205312 158392
rect 205468 158392 208860 158420
rect 205468 158352 205496 158392
rect 208854 158380 208860 158392
rect 208912 158380 208918 158432
rect 171100 158324 205220 158352
rect 205284 158324 205496 158352
rect 171100 158312 171106 158324
rect 162118 158244 162124 158296
rect 162176 158284 162182 158296
rect 169386 158284 169392 158296
rect 162176 158256 169392 158284
rect 162176 158244 162182 158256
rect 169386 158244 169392 158256
rect 169444 158244 169450 158296
rect 188798 158244 188804 158296
rect 188856 158284 188862 158296
rect 192662 158284 192668 158296
rect 188856 158256 192668 158284
rect 188856 158244 188862 158256
rect 192662 158244 192668 158256
rect 192720 158244 192726 158296
rect 194042 158244 194048 158296
rect 194100 158284 194106 158296
rect 194502 158284 194508 158296
rect 194100 158256 194508 158284
rect 194100 158244 194106 158256
rect 194502 158244 194508 158256
rect 194560 158244 194566 158296
rect 194704 158256 202874 158284
rect 160830 158176 160836 158228
rect 160888 158216 160894 158228
rect 177942 158216 177948 158228
rect 160888 158188 177948 158216
rect 160888 158176 160894 158188
rect 177942 158176 177948 158188
rect 178000 158176 178006 158228
rect 189166 158216 189172 158228
rect 186516 158188 189172 158216
rect 78674 158108 78680 158160
rect 78732 158148 78738 158160
rect 156690 158148 156696 158160
rect 78732 158120 156696 158148
rect 78732 158108 78738 158120
rect 156690 158108 156696 158120
rect 156748 158108 156754 158160
rect 160646 158108 160652 158160
rect 160704 158148 160710 158160
rect 171778 158148 171784 158160
rect 160704 158120 171784 158148
rect 160704 158108 160710 158120
rect 171778 158108 171784 158120
rect 171836 158108 171842 158160
rect 180518 158108 180524 158160
rect 180576 158148 180582 158160
rect 186314 158148 186320 158160
rect 180576 158120 186320 158148
rect 180576 158108 180582 158120
rect 186314 158108 186320 158120
rect 186372 158108 186378 158160
rect 60734 158040 60740 158092
rect 60792 158080 60798 158092
rect 157978 158080 157984 158092
rect 60792 158052 157984 158080
rect 60792 158040 60798 158052
rect 157978 158040 157984 158052
rect 158036 158080 158042 158092
rect 158622 158080 158628 158092
rect 158036 158052 158628 158080
rect 158036 158040 158042 158052
rect 158622 158040 158628 158052
rect 158680 158040 158686 158092
rect 161382 158040 161388 158092
rect 161440 158080 161446 158092
rect 161440 158052 166994 158080
rect 161440 158040 161446 158052
rect 4154 157972 4160 158024
rect 4212 158012 4218 158024
rect 161474 158012 161480 158024
rect 4212 157984 161480 158012
rect 4212 157972 4218 157984
rect 161474 157972 161480 157984
rect 161532 158012 161538 158024
rect 162578 158012 162584 158024
rect 161532 157984 162584 158012
rect 161532 157972 161538 157984
rect 162578 157972 162584 157984
rect 162636 157972 162642 158024
rect 166966 158012 166994 158052
rect 169386 158040 169392 158092
rect 169444 158080 169450 158092
rect 176102 158080 176108 158092
rect 169444 158052 176108 158080
rect 169444 158040 169450 158052
rect 176102 158040 176108 158052
rect 176160 158080 176166 158092
rect 176286 158080 176292 158092
rect 176160 158052 176292 158080
rect 176160 158040 176166 158052
rect 176286 158040 176292 158052
rect 176344 158040 176350 158092
rect 177390 158080 177396 158092
rect 176626 158052 177396 158080
rect 176010 158012 176016 158024
rect 166966 157984 176016 158012
rect 176010 157972 176016 157984
rect 176068 157972 176074 158024
rect 160738 157904 160744 157956
rect 160796 157944 160802 157956
rect 176626 157944 176654 158052
rect 177390 158040 177396 158052
rect 177448 158040 177454 158092
rect 180794 158040 180800 158092
rect 180852 158080 180858 158092
rect 186516 158080 186544 158188
rect 189166 158176 189172 158188
rect 189224 158176 189230 158228
rect 189350 158176 189356 158228
rect 189408 158216 189414 158228
rect 189408 158188 194548 158216
rect 189408 158176 189414 158188
rect 194520 158148 194548 158188
rect 194704 158148 194732 158256
rect 197906 158176 197912 158228
rect 197964 158216 197970 158228
rect 202414 158216 202420 158228
rect 197964 158188 202420 158216
rect 197964 158176 197970 158188
rect 202414 158176 202420 158188
rect 202472 158176 202478 158228
rect 202846 158216 202874 158256
rect 203702 158244 203708 158296
rect 203760 158284 203766 158296
rect 204162 158284 204168 158296
rect 203760 158256 204168 158284
rect 203760 158244 203766 158256
rect 204162 158244 204168 158256
rect 204220 158244 204226 158296
rect 204254 158216 204260 158228
rect 202846 158188 204260 158216
rect 204254 158176 204260 158188
rect 204312 158176 204318 158228
rect 205192 158216 205220 158324
rect 207842 158244 207848 158296
rect 207900 158284 207906 158296
rect 227438 158284 227444 158296
rect 207900 158256 227444 158284
rect 207900 158244 207906 158256
rect 227438 158244 227444 158256
rect 227496 158244 227502 158296
rect 208026 158216 208032 158228
rect 205192 158188 208032 158216
rect 208026 158176 208032 158188
rect 208084 158176 208090 158228
rect 208394 158176 208400 158228
rect 208452 158216 208458 158228
rect 246482 158216 246488 158228
rect 208452 158188 246488 158216
rect 208452 158176 208458 158188
rect 246482 158176 246488 158188
rect 246540 158176 246546 158228
rect 180852 158052 186544 158080
rect 186976 158120 191834 158148
rect 194520 158120 194732 158148
rect 180852 158040 180858 158052
rect 181346 157972 181352 158024
rect 181404 158012 181410 158024
rect 186976 158012 187004 158120
rect 191806 158080 191834 158120
rect 198274 158108 198280 158160
rect 198332 158148 198338 158160
rect 203242 158148 203248 158160
rect 198332 158120 203248 158148
rect 198332 158108 198338 158120
rect 203242 158108 203248 158120
rect 203300 158108 203306 158160
rect 207934 158108 207940 158160
rect 207992 158148 207998 158160
rect 246298 158148 246304 158160
rect 207992 158120 246304 158148
rect 207992 158108 207998 158120
rect 246298 158108 246304 158120
rect 246356 158108 246362 158160
rect 197998 158080 198004 158092
rect 191806 158052 198004 158080
rect 197998 158040 198004 158052
rect 198056 158040 198062 158092
rect 202782 158040 202788 158092
rect 202840 158040 202846 158092
rect 204806 158040 204812 158092
rect 204864 158080 204870 158092
rect 205358 158080 205364 158092
rect 204864 158052 205364 158080
rect 204864 158040 204870 158052
rect 205358 158040 205364 158052
rect 205416 158040 205422 158092
rect 206278 158080 206284 158092
rect 205468 158052 206284 158080
rect 181404 157984 187004 158012
rect 181404 157972 181410 157984
rect 189166 157972 189172 158024
rect 189224 158012 189230 158024
rect 197078 158012 197084 158024
rect 189224 157984 197084 158012
rect 189224 157972 189230 157984
rect 197078 157972 197084 157984
rect 197136 157972 197142 158024
rect 202800 158012 202828 158040
rect 205468 158012 205496 158052
rect 206278 158040 206284 158052
rect 206336 158040 206342 158092
rect 208026 158040 208032 158092
rect 208084 158080 208090 158092
rect 250438 158080 250444 158092
rect 208084 158052 250444 158080
rect 208084 158040 208090 158052
rect 250438 158040 250444 158052
rect 250496 158040 250502 158092
rect 207474 158012 207480 158024
rect 202800 157984 205496 158012
rect 205606 157984 207480 158012
rect 160796 157916 176654 157944
rect 160796 157904 160802 157916
rect 180518 157904 180524 157956
rect 180576 157944 180582 157956
rect 180702 157944 180708 157956
rect 180576 157916 180708 157944
rect 180576 157904 180582 157916
rect 180702 157904 180708 157916
rect 180760 157904 180766 157956
rect 185210 157904 185216 157956
rect 185268 157944 185274 157956
rect 194870 157944 194876 157956
rect 185268 157916 194876 157944
rect 185268 157904 185274 157916
rect 194870 157904 194876 157916
rect 194928 157904 194934 157956
rect 196158 157904 196164 157956
rect 196216 157944 196222 157956
rect 198182 157944 198188 157956
rect 196216 157916 198188 157944
rect 196216 157904 196222 157916
rect 198182 157904 198188 157916
rect 198240 157904 198246 157956
rect 202598 157944 202604 157956
rect 199488 157916 202604 157944
rect 148318 157836 148324 157888
rect 148376 157876 148382 157888
rect 165614 157876 165620 157888
rect 148376 157848 165620 157876
rect 148376 157836 148382 157848
rect 165614 157836 165620 157848
rect 165672 157836 165678 157888
rect 167822 157836 167828 157888
rect 167880 157876 167886 157888
rect 168558 157876 168564 157888
rect 167880 157848 168564 157876
rect 167880 157836 167886 157848
rect 168558 157836 168564 157848
rect 168616 157836 168622 157888
rect 176010 157836 176016 157888
rect 176068 157876 176074 157888
rect 176286 157876 176292 157888
rect 176068 157848 176292 157876
rect 176068 157836 176074 157848
rect 176286 157836 176292 157848
rect 176344 157836 176350 157888
rect 185854 157836 185860 157888
rect 185912 157876 185918 157888
rect 186038 157876 186044 157888
rect 185912 157848 186044 157876
rect 185912 157836 185918 157848
rect 186038 157836 186044 157848
rect 186096 157836 186102 157888
rect 186314 157836 186320 157888
rect 186372 157876 186378 157888
rect 195514 157876 195520 157888
rect 186372 157848 195520 157876
rect 186372 157836 186378 157848
rect 195514 157836 195520 157848
rect 195572 157836 195578 157888
rect 171778 157768 171784 157820
rect 171836 157808 171842 157820
rect 177666 157808 177672 157820
rect 171836 157780 177672 157808
rect 171836 157768 171842 157780
rect 177666 157768 177672 157780
rect 177724 157768 177730 157820
rect 181990 157768 181996 157820
rect 182048 157808 182054 157820
rect 182048 157780 186314 157808
rect 182048 157768 182054 157780
rect 124858 157700 124864 157752
rect 124916 157740 124922 157752
rect 160738 157740 160744 157752
rect 124916 157712 160744 157740
rect 124916 157700 124922 157712
rect 160738 157700 160744 157712
rect 160796 157700 160802 157752
rect 163038 157700 163044 157752
rect 163096 157740 163102 157752
rect 165798 157740 165804 157752
rect 163096 157712 165804 157740
rect 163096 157700 163102 157712
rect 165798 157700 165804 157712
rect 165856 157700 165862 157752
rect 166074 157700 166080 157752
rect 166132 157740 166138 157752
rect 167178 157740 167184 157752
rect 166132 157712 167184 157740
rect 166132 157700 166138 157712
rect 167178 157700 167184 157712
rect 167236 157700 167242 157752
rect 184382 157700 184388 157752
rect 184440 157740 184446 157752
rect 186038 157740 186044 157752
rect 184440 157712 186044 157740
rect 184440 157700 184446 157712
rect 186038 157700 186044 157712
rect 186096 157700 186102 157752
rect 186286 157740 186314 157780
rect 192110 157768 192116 157820
rect 192168 157808 192174 157820
rect 194134 157808 194140 157820
rect 192168 157780 194140 157808
rect 192168 157768 192174 157780
rect 194134 157768 194140 157780
rect 194192 157768 194198 157820
rect 195146 157768 195152 157820
rect 195204 157808 195210 157820
rect 197722 157808 197728 157820
rect 195204 157780 197728 157808
rect 195204 157768 195210 157780
rect 197722 157768 197728 157780
rect 197780 157768 197786 157820
rect 192202 157740 192208 157752
rect 186286 157712 192208 157740
rect 192202 157700 192208 157712
rect 192260 157700 192266 157752
rect 194410 157700 194416 157752
rect 194468 157740 194474 157752
rect 196802 157740 196808 157752
rect 194468 157712 196808 157740
rect 194468 157700 194474 157712
rect 196802 157700 196808 157712
rect 196860 157700 196866 157752
rect 160922 157632 160928 157684
rect 160980 157672 160986 157684
rect 177114 157672 177120 157684
rect 160980 157644 177120 157672
rect 160980 157632 160986 157644
rect 177114 157632 177120 157644
rect 177172 157672 177178 157684
rect 181346 157672 181352 157684
rect 177172 157644 181352 157672
rect 177172 157632 177178 157644
rect 181346 157632 181352 157644
rect 181404 157632 181410 157684
rect 183278 157632 183284 157684
rect 183336 157672 183342 157684
rect 184474 157672 184480 157684
rect 183336 157644 184480 157672
rect 183336 157632 183342 157644
rect 184474 157632 184480 157644
rect 184532 157632 184538 157684
rect 185762 157632 185768 157684
rect 185820 157672 185826 157684
rect 187142 157672 187148 157684
rect 185820 157644 187148 157672
rect 185820 157632 185826 157644
rect 187142 157632 187148 157644
rect 187200 157632 187206 157684
rect 190454 157632 190460 157684
rect 190512 157672 190518 157684
rect 191098 157672 191104 157684
rect 190512 157644 191104 157672
rect 190512 157632 190518 157644
rect 191098 157632 191104 157644
rect 191156 157632 191162 157684
rect 195422 157632 195428 157684
rect 195480 157672 195486 157684
rect 199378 157672 199384 157684
rect 195480 157644 199384 157672
rect 195480 157632 195486 157644
rect 199378 157632 199384 157644
rect 199436 157632 199442 157684
rect 165062 157564 165068 157616
rect 165120 157604 165126 157616
rect 199488 157604 199516 157916
rect 202598 157904 202604 157916
rect 202656 157904 202662 157956
rect 202782 157904 202788 157956
rect 202840 157944 202846 157956
rect 205606 157944 205634 157984
rect 207474 157972 207480 157984
rect 207532 157972 207538 158024
rect 208486 157972 208492 158024
rect 208544 158012 208550 158024
rect 253566 158012 253572 158024
rect 208544 157984 253572 158012
rect 208544 157972 208550 157984
rect 253566 157972 253572 157984
rect 253624 157972 253630 158024
rect 202840 157916 205634 157944
rect 202840 157904 202846 157916
rect 207014 157904 207020 157956
rect 207072 157944 207078 157956
rect 221550 157944 221556 157956
rect 207072 157916 221556 157944
rect 207072 157904 207078 157916
rect 221550 157904 221556 157916
rect 221608 157904 221614 157956
rect 199562 157836 199568 157888
rect 199620 157876 199626 157888
rect 199620 157848 202460 157876
rect 199620 157836 199626 157848
rect 202432 157808 202460 157848
rect 207106 157836 207112 157888
rect 207164 157876 207170 157888
rect 208210 157876 208216 157888
rect 207164 157848 208216 157876
rect 207164 157836 207170 157848
rect 208210 157836 208216 157848
rect 208268 157836 208274 157888
rect 260282 157808 260288 157820
rect 202432 157780 260288 157808
rect 260282 157768 260288 157780
rect 260340 157768 260346 157820
rect 202138 157700 202144 157752
rect 202196 157740 202202 157752
rect 210786 157740 210792 157752
rect 202196 157712 210792 157740
rect 202196 157700 202202 157712
rect 210786 157700 210792 157712
rect 210844 157700 210850 157752
rect 200942 157632 200948 157684
rect 201000 157672 201006 157684
rect 209590 157672 209596 157684
rect 201000 157644 209596 157672
rect 201000 157632 201006 157644
rect 209590 157632 209596 157644
rect 209648 157632 209654 157684
rect 210878 157604 210884 157616
rect 165120 157576 199516 157604
rect 200408 157576 210884 157604
rect 165120 157564 165126 157576
rect 163406 157536 163412 157548
rect 154546 157508 163412 157536
rect 152918 157292 152924 157344
rect 152976 157332 152982 157344
rect 154546 157332 154574 157508
rect 163406 157496 163412 157508
rect 163464 157496 163470 157548
rect 164326 157496 164332 157548
rect 164384 157536 164390 157548
rect 164878 157536 164884 157548
rect 164384 157508 164884 157536
rect 164384 157496 164390 157508
rect 164878 157496 164884 157508
rect 164936 157496 164942 157548
rect 165614 157496 165620 157548
rect 165672 157536 165678 157548
rect 198274 157536 198280 157548
rect 165672 157508 198280 157536
rect 165672 157496 165678 157508
rect 198274 157496 198280 157508
rect 198332 157496 198338 157548
rect 158622 157428 158628 157480
rect 158680 157468 158686 157480
rect 166074 157468 166080 157480
rect 158680 157440 166080 157468
rect 158680 157428 158686 157440
rect 166074 157428 166080 157440
rect 166132 157428 166138 157480
rect 170398 157428 170404 157480
rect 170456 157468 170462 157480
rect 171042 157468 171048 157480
rect 170456 157440 171048 157468
rect 170456 157428 170462 157440
rect 171042 157428 171048 157440
rect 171100 157428 171106 157480
rect 200408 157468 200436 157576
rect 210878 157564 210884 157576
rect 210936 157564 210942 157616
rect 205634 157496 205640 157548
rect 205692 157536 205698 157548
rect 205818 157536 205824 157548
rect 205692 157508 205824 157536
rect 205692 157496 205698 157508
rect 205818 157496 205824 157508
rect 205876 157496 205882 157548
rect 207198 157496 207204 157548
rect 207256 157536 207262 157548
rect 214926 157536 214932 157548
rect 207256 157508 214932 157536
rect 207256 157496 207262 157508
rect 214926 157496 214932 157508
rect 214984 157496 214990 157548
rect 171796 157440 200436 157468
rect 161014 157360 161020 157412
rect 161072 157400 161078 157412
rect 164050 157400 164056 157412
rect 161072 157372 164056 157400
rect 161072 157360 161078 157372
rect 164050 157360 164056 157372
rect 164108 157400 164114 157412
rect 171796 157400 171824 157440
rect 211062 157400 211068 157412
rect 164108 157372 171824 157400
rect 173866 157372 211068 157400
rect 164108 157360 164114 157372
rect 152976 157304 154574 157332
rect 152976 157292 152982 157304
rect 162762 157292 162768 157344
rect 162820 157332 162826 157344
rect 163038 157332 163044 157344
rect 162820 157304 163044 157332
rect 162820 157292 162826 157304
rect 163038 157292 163044 157304
rect 163096 157292 163102 157344
rect 163498 157292 163504 157344
rect 163556 157332 163562 157344
rect 170122 157332 170128 157344
rect 163556 157304 170128 157332
rect 163556 157292 163562 157304
rect 170122 157292 170128 157304
rect 170180 157292 170186 157344
rect 154298 157224 154304 157276
rect 154356 157264 154362 157276
rect 154356 157236 162072 157264
rect 154356 157224 154362 157236
rect 159634 157156 159640 157208
rect 159692 157196 159698 157208
rect 161842 157196 161848 157208
rect 159692 157168 161848 157196
rect 159692 157156 159698 157168
rect 161842 157156 161848 157168
rect 161900 157156 161906 157208
rect 162044 157196 162072 157236
rect 162118 157224 162124 157276
rect 162176 157264 162182 157276
rect 166534 157264 166540 157276
rect 162176 157236 166540 157264
rect 162176 157224 162182 157236
rect 166534 157224 166540 157236
rect 166592 157224 166598 157276
rect 169938 157224 169944 157276
rect 169996 157264 170002 157276
rect 171042 157264 171048 157276
rect 169996 157236 171048 157264
rect 169996 157224 170002 157236
rect 171042 157224 171048 157236
rect 171100 157224 171106 157276
rect 163406 157196 163412 157208
rect 162044 157168 163412 157196
rect 163406 157156 163412 157168
rect 163464 157196 163470 157208
rect 163958 157196 163964 157208
rect 163464 157168 163964 157196
rect 163464 157156 163470 157168
rect 163958 157156 163964 157168
rect 164016 157156 164022 157208
rect 164878 157156 164884 157208
rect 164936 157196 164942 157208
rect 173866 157196 173894 157372
rect 211062 157360 211068 157372
rect 211120 157360 211126 157412
rect 187970 157292 187976 157344
rect 188028 157332 188034 157344
rect 208394 157332 208400 157344
rect 188028 157304 208400 157332
rect 188028 157292 188034 157304
rect 208394 157292 208400 157304
rect 208452 157292 208458 157344
rect 190730 157224 190736 157276
rect 190788 157264 190794 157276
rect 200942 157264 200948 157276
rect 190788 157236 200948 157264
rect 190788 157224 190794 157236
rect 200942 157224 200948 157236
rect 201000 157224 201006 157276
rect 202230 157224 202236 157276
rect 202288 157264 202294 157276
rect 202782 157264 202788 157276
rect 202288 157236 202788 157264
rect 202288 157224 202294 157236
rect 202782 157224 202788 157236
rect 202840 157224 202846 157276
rect 164936 157168 173894 157196
rect 164936 157156 164942 157168
rect 190178 157156 190184 157208
rect 190236 157196 190242 157208
rect 191650 157196 191656 157208
rect 190236 157168 191656 157196
rect 190236 157156 190242 157168
rect 191650 157156 191656 157168
rect 191708 157156 191714 157208
rect 192386 157156 192392 157208
rect 192444 157196 192450 157208
rect 206186 157196 206192 157208
rect 192444 157168 206192 157196
rect 192444 157156 192450 157168
rect 206186 157156 206192 157168
rect 206244 157156 206250 157208
rect 160738 157088 160744 157140
rect 160796 157128 160802 157140
rect 171594 157128 171600 157140
rect 160796 157100 171600 157128
rect 160796 157088 160802 157100
rect 171594 157088 171600 157100
rect 171652 157088 171658 157140
rect 183094 157088 183100 157140
rect 183152 157128 183158 157140
rect 242158 157128 242164 157140
rect 183152 157100 242164 157128
rect 183152 157088 183158 157100
rect 242158 157088 242164 157100
rect 242216 157088 242222 157140
rect 143534 157020 143540 157072
rect 143592 157060 143598 157072
rect 173526 157060 173532 157072
rect 143592 157032 173532 157060
rect 143592 157020 143598 157032
rect 173526 157020 173532 157032
rect 173584 157060 173590 157072
rect 213178 157060 213184 157072
rect 173584 157032 213184 157060
rect 173584 157020 173590 157032
rect 213178 157020 213184 157032
rect 213236 157020 213242 157072
rect 130378 156952 130384 157004
rect 130436 156992 130442 157004
rect 161474 156992 161480 157004
rect 130436 156964 161480 156992
rect 130436 156952 130442 156964
rect 161474 156952 161480 156964
rect 161532 156952 161538 157004
rect 163498 156992 163504 157004
rect 161768 156964 163504 156992
rect 99374 156884 99380 156936
rect 99432 156924 99438 156936
rect 161768 156924 161796 156964
rect 163498 156952 163504 156964
rect 163556 156952 163562 157004
rect 163590 156952 163596 157004
rect 163648 156992 163654 157004
rect 164142 156992 164148 157004
rect 163648 156964 164148 156992
rect 163648 156952 163654 156964
rect 164142 156952 164148 156964
rect 164200 156952 164206 157004
rect 165798 156952 165804 157004
rect 165856 156992 165862 157004
rect 166166 156992 166172 157004
rect 165856 156964 166172 156992
rect 165856 156952 165862 156964
rect 166166 156952 166172 156964
rect 166224 156952 166230 157004
rect 170490 156952 170496 157004
rect 170548 156992 170554 157004
rect 171042 156992 171048 157004
rect 170548 156964 171048 156992
rect 170548 156952 170554 156964
rect 171042 156952 171048 156964
rect 171100 156952 171106 157004
rect 179046 156952 179052 157004
rect 179104 156992 179110 157004
rect 213914 156992 213920 157004
rect 179104 156964 213920 156992
rect 179104 156952 179110 156964
rect 213914 156952 213920 156964
rect 213972 156952 213978 157004
rect 99432 156896 161796 156924
rect 99432 156884 99438 156896
rect 161842 156884 161848 156936
rect 161900 156924 161906 156936
rect 165614 156924 165620 156936
rect 161900 156896 165620 156924
rect 161900 156884 161906 156896
rect 165614 156884 165620 156896
rect 165672 156924 165678 156936
rect 166626 156924 166632 156936
rect 165672 156896 166632 156924
rect 165672 156884 165678 156896
rect 166626 156884 166632 156896
rect 166684 156884 166690 156936
rect 196250 156884 196256 156936
rect 196308 156924 196314 156936
rect 202230 156924 202236 156936
rect 196308 156896 202236 156924
rect 196308 156884 196314 156896
rect 202230 156884 202236 156896
rect 202288 156884 202294 156936
rect 205818 156884 205824 156936
rect 205876 156924 205882 156936
rect 239858 156924 239864 156936
rect 205876 156896 239864 156924
rect 205876 156884 205882 156896
rect 239858 156884 239864 156896
rect 239916 156884 239922 156936
rect 85574 156816 85580 156868
rect 85632 156856 85638 156868
rect 169018 156856 169024 156868
rect 85632 156828 169024 156856
rect 85632 156816 85638 156828
rect 169018 156816 169024 156828
rect 169076 156816 169082 156868
rect 179598 156816 179604 156868
rect 179656 156856 179662 156868
rect 200666 156856 200672 156868
rect 179656 156828 200672 156856
rect 179656 156816 179662 156828
rect 200666 156816 200672 156828
rect 200724 156816 200730 156868
rect 200942 156816 200948 156868
rect 201000 156856 201006 156868
rect 209222 156856 209228 156868
rect 201000 156828 209228 156856
rect 201000 156816 201006 156828
rect 209222 156816 209228 156828
rect 209280 156816 209286 156868
rect 81434 156748 81440 156800
rect 81492 156788 81498 156800
rect 168650 156788 168656 156800
rect 81492 156760 168656 156788
rect 81492 156748 81498 156760
rect 168650 156748 168656 156760
rect 168708 156748 168714 156800
rect 178770 156748 178776 156800
rect 178828 156788 178834 156800
rect 209682 156788 209688 156800
rect 178828 156760 209688 156788
rect 178828 156748 178834 156760
rect 209682 156748 209688 156760
rect 209740 156788 209746 156800
rect 215846 156788 215852 156800
rect 209740 156760 215852 156788
rect 209740 156748 209746 156760
rect 215846 156748 215852 156760
rect 215904 156748 215910 156800
rect 74534 156680 74540 156732
rect 74592 156720 74598 156732
rect 168190 156720 168196 156732
rect 74592 156692 168196 156720
rect 74592 156680 74598 156692
rect 168190 156680 168196 156692
rect 168248 156680 168254 156732
rect 182542 156720 182548 156732
rect 176626 156692 182548 156720
rect 67634 156612 67640 156664
rect 67692 156652 67698 156664
rect 167638 156652 167644 156664
rect 67692 156624 167644 156652
rect 67692 156612 67698 156624
rect 167638 156612 167644 156624
rect 167696 156612 167702 156664
rect 176626 156596 176654 156692
rect 182542 156680 182548 156692
rect 182600 156720 182606 156732
rect 182600 156692 191236 156720
rect 182600 156680 182606 156692
rect 191208 156652 191236 156692
rect 191374 156680 191380 156732
rect 191432 156720 191438 156732
rect 220354 156720 220360 156732
rect 191432 156692 220360 156720
rect 191432 156680 191438 156692
rect 220354 156680 220360 156692
rect 220412 156680 220418 156732
rect 220262 156652 220268 156664
rect 191208 156624 220268 156652
rect 220262 156612 220268 156624
rect 220320 156612 220326 156664
rect 245010 156612 245016 156664
rect 245068 156652 245074 156664
rect 266998 156652 267004 156664
rect 245068 156624 267004 156652
rect 245068 156612 245074 156624
rect 266998 156612 267004 156624
rect 267056 156612 267062 156664
rect 289170 156652 289176 156664
rect 277366 156624 289176 156652
rect 161474 156544 161480 156596
rect 161532 156584 161538 156596
rect 169938 156584 169944 156596
rect 161532 156556 169944 156584
rect 161532 156544 161538 156556
rect 169938 156544 169944 156556
rect 169996 156544 170002 156596
rect 176562 156544 176568 156596
rect 176620 156556 176654 156596
rect 176620 156544 176626 156556
rect 176838 156544 176844 156596
rect 176896 156584 176902 156596
rect 185762 156584 185768 156596
rect 176896 156556 185768 156584
rect 176896 156544 176902 156556
rect 185762 156544 185768 156556
rect 185820 156584 185826 156596
rect 191374 156584 191380 156596
rect 185820 156556 191380 156584
rect 185820 156544 185826 156556
rect 191374 156544 191380 156556
rect 191432 156544 191438 156596
rect 200666 156544 200672 156596
rect 200724 156584 200730 156596
rect 211798 156584 211804 156596
rect 200724 156556 211804 156584
rect 200724 156544 200730 156556
rect 211798 156544 211804 156556
rect 211856 156584 211862 156596
rect 212350 156584 212356 156596
rect 211856 156556 212356 156584
rect 211856 156544 211862 156556
rect 212350 156544 212356 156556
rect 212408 156544 212414 156596
rect 154206 156476 154212 156528
rect 154264 156516 154270 156528
rect 164234 156516 164240 156528
rect 154264 156488 164240 156516
rect 154264 156476 154270 156488
rect 164234 156476 164240 156488
rect 164292 156516 164298 156528
rect 165246 156516 165252 156528
rect 164292 156488 165252 156516
rect 164292 156476 164298 156488
rect 165246 156476 165252 156488
rect 165304 156476 165310 156528
rect 185394 156476 185400 156528
rect 185452 156516 185458 156528
rect 275922 156516 275928 156528
rect 185452 156488 275928 156516
rect 185452 156476 185458 156488
rect 275922 156476 275928 156488
rect 275980 156516 275986 156528
rect 277366 156516 277394 156624
rect 289170 156612 289176 156624
rect 289228 156612 289234 156664
rect 275980 156488 277394 156516
rect 275980 156476 275986 156488
rect 159542 156408 159548 156460
rect 159600 156448 159606 156460
rect 166994 156448 167000 156460
rect 159600 156420 167000 156448
rect 159600 156408 159606 156420
rect 166994 156408 167000 156420
rect 167052 156448 167058 156460
rect 168006 156448 168012 156460
rect 167052 156420 168012 156448
rect 167052 156408 167058 156420
rect 168006 156408 168012 156420
rect 168064 156408 168070 156460
rect 169662 156408 169668 156460
rect 169720 156448 169726 156460
rect 170674 156448 170680 156460
rect 169720 156420 170680 156448
rect 169720 156408 169726 156420
rect 170674 156408 170680 156420
rect 170732 156408 170738 156460
rect 172974 156408 172980 156460
rect 173032 156448 173038 156460
rect 232958 156448 232964 156460
rect 173032 156420 232964 156448
rect 173032 156408 173038 156420
rect 232958 156408 232964 156420
rect 233016 156408 233022 156460
rect 175366 156340 175372 156392
rect 175424 156380 175430 156392
rect 176378 156380 176384 156392
rect 175424 156352 176384 156380
rect 175424 156340 175430 156352
rect 176378 156340 176384 156352
rect 176436 156380 176442 156392
rect 235166 156380 235172 156392
rect 176436 156352 235172 156380
rect 176436 156340 176442 156352
rect 235166 156340 235172 156352
rect 235224 156340 235230 156392
rect 184106 156272 184112 156324
rect 184164 156312 184170 156324
rect 207014 156312 207020 156324
rect 184164 156284 207020 156312
rect 184164 156272 184170 156284
rect 207014 156272 207020 156284
rect 207072 156272 207078 156324
rect 176286 156068 176292 156120
rect 176344 156108 176350 156120
rect 179414 156108 179420 156120
rect 176344 156080 179420 156108
rect 176344 156068 176350 156080
rect 179414 156068 179420 156080
rect 179472 156068 179478 156120
rect 191006 156000 191012 156052
rect 191064 156040 191070 156052
rect 191190 156040 191196 156052
rect 191064 156012 191196 156040
rect 191064 156000 191070 156012
rect 191190 156000 191196 156012
rect 191248 156000 191254 156052
rect 164418 155932 164424 155984
rect 164476 155972 164482 155984
rect 165522 155972 165528 155984
rect 164476 155944 165528 155972
rect 164476 155932 164482 155944
rect 165522 155932 165528 155944
rect 165580 155932 165586 155984
rect 189902 155932 189908 155984
rect 189960 155972 189966 155984
rect 191374 155972 191380 155984
rect 189960 155944 191380 155972
rect 189960 155932 189966 155944
rect 191374 155932 191380 155944
rect 191432 155932 191438 155984
rect 195808 155944 196112 155972
rect 149054 155864 149060 155916
rect 149112 155904 149118 155916
rect 150342 155904 150348 155916
rect 149112 155876 150348 155904
rect 149112 155864 149118 155876
rect 150342 155864 150348 155876
rect 150400 155904 150406 155916
rect 164694 155904 164700 155916
rect 150400 155876 164700 155904
rect 150400 155864 150406 155876
rect 164694 155864 164700 155876
rect 164752 155864 164758 155916
rect 193582 155864 193588 155916
rect 193640 155904 193646 155916
rect 195808 155904 195836 155944
rect 193640 155876 195836 155904
rect 193640 155864 193646 155876
rect 195882 155864 195888 155916
rect 195940 155904 195946 155916
rect 196084 155904 196112 155944
rect 206370 155932 206376 155984
rect 206428 155972 206434 155984
rect 206922 155972 206928 155984
rect 206428 155944 206928 155972
rect 206428 155932 206434 155944
rect 206922 155932 206928 155944
rect 206980 155932 206986 155984
rect 269758 155932 269764 155984
rect 269816 155972 269822 155984
rect 518894 155972 518900 155984
rect 269816 155944 518900 155972
rect 269816 155932 269822 155944
rect 518894 155932 518900 155944
rect 518952 155932 518958 155984
rect 272150 155904 272156 155916
rect 195940 155864 195974 155904
rect 196084 155876 272156 155904
rect 272150 155864 272156 155876
rect 272208 155904 272214 155916
rect 272334 155904 272340 155916
rect 272208 155876 272340 155904
rect 272208 155864 272214 155876
rect 272334 155864 272340 155876
rect 272392 155864 272398 155916
rect 171962 155836 171968 155848
rect 161446 155808 171968 155836
rect 125594 155592 125600 155644
rect 125652 155632 125658 155644
rect 159818 155632 159824 155644
rect 125652 155604 159824 155632
rect 125652 155592 125658 155604
rect 159818 155592 159824 155604
rect 159876 155632 159882 155644
rect 161446 155632 161474 155808
rect 171962 155796 171968 155808
rect 172020 155796 172026 155848
rect 185486 155796 185492 155848
rect 185544 155836 185550 155848
rect 191006 155836 191012 155848
rect 185544 155808 191012 155836
rect 185544 155796 185550 155808
rect 191006 155796 191012 155808
rect 191064 155796 191070 155848
rect 195946 155836 195974 155864
rect 196986 155836 196992 155848
rect 195946 155808 196992 155836
rect 196986 155796 196992 155808
rect 197044 155796 197050 155848
rect 203058 155796 203064 155848
rect 203116 155836 203122 155848
rect 271230 155836 271236 155848
rect 203116 155808 271236 155836
rect 203116 155796 203122 155808
rect 271230 155796 271236 155808
rect 271288 155836 271294 155848
rect 271782 155836 271788 155848
rect 271288 155808 271788 155836
rect 271288 155796 271294 155808
rect 271782 155796 271788 155808
rect 271840 155796 271846 155848
rect 164694 155728 164700 155780
rect 164752 155768 164758 155780
rect 165338 155768 165344 155780
rect 164752 155740 165344 155768
rect 164752 155728 164758 155740
rect 165338 155728 165344 155740
rect 165396 155728 165402 155780
rect 190270 155728 190276 155780
rect 190328 155768 190334 155780
rect 214834 155768 214840 155780
rect 190328 155740 214840 155768
rect 190328 155728 190334 155740
rect 214834 155728 214840 155740
rect 214892 155728 214898 155780
rect 200666 155660 200672 155712
rect 200724 155700 200730 155712
rect 207198 155700 207204 155712
rect 200724 155672 207204 155700
rect 200724 155660 200730 155672
rect 207198 155660 207204 155672
rect 207256 155660 207262 155712
rect 159876 155604 161474 155632
rect 159876 155592 159882 155604
rect 168558 155592 168564 155644
rect 168616 155632 168622 155644
rect 175366 155632 175372 155644
rect 168616 155604 175372 155632
rect 168616 155592 168622 155604
rect 175366 155592 175372 155604
rect 175424 155592 175430 155644
rect 180150 155592 180156 155644
rect 180208 155632 180214 155644
rect 222102 155632 222108 155644
rect 180208 155604 222108 155632
rect 180208 155592 180214 155604
rect 222102 155592 222108 155604
rect 222160 155632 222166 155644
rect 225598 155632 225604 155644
rect 222160 155604 225604 155632
rect 222160 155592 222166 155604
rect 225598 155592 225604 155604
rect 225656 155592 225662 155644
rect 137278 155524 137284 155576
rect 137336 155564 137342 155576
rect 172790 155564 172796 155576
rect 137336 155536 172796 155564
rect 137336 155524 137342 155536
rect 172790 155524 172796 155536
rect 172848 155524 172854 155576
rect 175182 155524 175188 155576
rect 175240 155564 175246 155576
rect 216122 155564 216128 155576
rect 175240 155536 216128 155564
rect 175240 155524 175246 155536
rect 216122 155524 216128 155536
rect 216180 155524 216186 155576
rect 115198 155456 115204 155508
rect 115256 155496 115262 155508
rect 150434 155496 150440 155508
rect 115256 155468 150440 155496
rect 115256 155456 115262 155468
rect 150434 155456 150440 155468
rect 150492 155456 150498 155508
rect 175366 155456 175372 155508
rect 175424 155496 175430 155508
rect 175734 155496 175740 155508
rect 175424 155468 175740 155496
rect 175424 155456 175430 155468
rect 175734 155456 175740 155468
rect 175792 155496 175798 155508
rect 216030 155496 216036 155508
rect 175792 155468 216036 155496
rect 175792 155456 175798 155468
rect 216030 155456 216036 155468
rect 216088 155456 216094 155508
rect 135254 155388 135260 155440
rect 135312 155428 135318 155440
rect 172974 155428 172980 155440
rect 135312 155400 172980 155428
rect 135312 155388 135318 155400
rect 172974 155388 172980 155400
rect 173032 155388 173038 155440
rect 179322 155388 179328 155440
rect 179380 155428 179386 155440
rect 210418 155428 210424 155440
rect 179380 155400 210424 155428
rect 179380 155388 179386 155400
rect 210418 155388 210424 155400
rect 210476 155388 210482 155440
rect 106274 155320 106280 155372
rect 106332 155360 106338 155372
rect 169754 155360 169760 155372
rect 106332 155332 169760 155360
rect 106332 155320 106338 155332
rect 169754 155320 169760 155332
rect 169812 155320 169818 155372
rect 191006 155320 191012 155372
rect 191064 155360 191070 155372
rect 207842 155360 207848 155372
rect 191064 155332 207848 155360
rect 191064 155320 191070 155332
rect 207842 155320 207848 155332
rect 207900 155320 207906 155372
rect 272334 155320 272340 155372
rect 272392 155360 272398 155372
rect 355318 155360 355324 155372
rect 272392 155332 355324 155360
rect 272392 155320 272398 155332
rect 355318 155320 355324 155332
rect 355376 155320 355382 155372
rect 26234 155252 26240 155304
rect 26292 155292 26298 155304
rect 149054 155292 149060 155304
rect 26292 155264 149060 155292
rect 26292 155252 26298 155264
rect 149054 155252 149060 155264
rect 149112 155252 149118 155304
rect 150434 155252 150440 155304
rect 150492 155292 150498 155304
rect 174170 155292 174176 155304
rect 150492 155264 174176 155292
rect 150492 155252 150498 155264
rect 174170 155252 174176 155264
rect 174228 155252 174234 155304
rect 177942 155252 177948 155304
rect 178000 155292 178006 155304
rect 193582 155292 193588 155304
rect 178000 155264 193588 155292
rect 178000 155252 178006 155264
rect 193582 155252 193588 155264
rect 193640 155252 193646 155304
rect 270218 155252 270224 155304
rect 270276 155292 270282 155304
rect 494054 155292 494060 155304
rect 270276 155264 494060 155292
rect 270276 155252 270282 155264
rect 494054 155252 494060 155264
rect 494112 155252 494118 155304
rect 13078 155184 13084 155236
rect 13136 155224 13142 155236
rect 152918 155224 152924 155236
rect 13136 155196 152924 155224
rect 13136 155184 13142 155196
rect 152918 155184 152924 155196
rect 152976 155184 152982 155236
rect 178034 155184 178040 155236
rect 178092 155224 178098 155236
rect 191006 155224 191012 155236
rect 178092 155196 191012 155224
rect 178092 155184 178098 155196
rect 191006 155184 191012 155196
rect 191064 155184 191070 155236
rect 271782 155184 271788 155236
rect 271840 155224 271846 155236
rect 522298 155224 522304 155236
rect 271840 155196 522304 155224
rect 271840 155184 271846 155196
rect 522298 155184 522304 155196
rect 522356 155184 522362 155236
rect 193030 155116 193036 155168
rect 193088 155156 193094 155168
rect 200666 155156 200672 155168
rect 193088 155128 200672 155156
rect 193088 155116 193094 155128
rect 200666 155116 200672 155128
rect 200724 155116 200730 155168
rect 201678 155116 201684 155168
rect 201736 155156 201742 155168
rect 202690 155156 202696 155168
rect 201736 155128 202696 155156
rect 201736 155116 201742 155128
rect 202690 155116 202696 155128
rect 202748 155156 202754 155168
rect 267918 155156 267924 155168
rect 202748 155128 267924 155156
rect 202748 155116 202754 155128
rect 267918 155116 267924 155128
rect 267976 155116 267982 155168
rect 179874 155048 179880 155100
rect 179932 155088 179938 155100
rect 212442 155088 212448 155100
rect 179932 155060 212448 155088
rect 179932 155048 179938 155060
rect 212442 155048 212448 155060
rect 212500 155088 212506 155100
rect 213178 155088 213184 155100
rect 212500 155060 213184 155088
rect 212500 155048 212506 155060
rect 213178 155048 213184 155060
rect 213236 155048 213242 155100
rect 174170 154980 174176 155032
rect 174228 155020 174234 155032
rect 234430 155020 234436 155032
rect 174228 154992 234436 155020
rect 174228 154980 174234 154992
rect 234430 154980 234436 154992
rect 234488 154980 234494 155032
rect 185854 154912 185860 154964
rect 185912 154952 185918 154964
rect 207934 154952 207940 154964
rect 185912 154924 207940 154952
rect 185912 154912 185918 154924
rect 207934 154912 207940 154924
rect 207992 154912 207998 154964
rect 184658 154844 184664 154896
rect 184716 154884 184722 154896
rect 190270 154884 190276 154896
rect 184716 154856 190276 154884
rect 184716 154844 184722 154856
rect 190270 154844 190276 154856
rect 190328 154844 190334 154896
rect 190914 154844 190920 154896
rect 190972 154884 190978 154896
rect 208026 154884 208032 154896
rect 190972 154856 208032 154884
rect 190972 154844 190978 154856
rect 208026 154844 208032 154856
rect 208084 154844 208090 154896
rect 191006 154708 191012 154760
rect 191064 154748 191070 154760
rect 201954 154748 201960 154760
rect 191064 154720 201960 154748
rect 191064 154708 191070 154720
rect 201954 154708 201960 154720
rect 202012 154708 202018 154760
rect 200574 154640 200580 154692
rect 200632 154680 200638 154692
rect 203058 154680 203064 154692
rect 200632 154652 203064 154680
rect 200632 154640 200638 154652
rect 203058 154640 203064 154652
rect 203116 154640 203122 154692
rect 174722 154572 174728 154624
rect 174780 154612 174786 154624
rect 175182 154612 175188 154624
rect 174780 154584 175188 154612
rect 174780 154572 174786 154584
rect 175182 154572 175188 154584
rect 175240 154572 175246 154624
rect 194502 154572 194508 154624
rect 194560 154612 194566 154624
rect 200666 154612 200672 154624
rect 194560 154584 200672 154612
rect 194560 154572 194566 154584
rect 200666 154572 200672 154584
rect 200724 154572 200730 154624
rect 201218 154504 201224 154556
rect 201276 154544 201282 154556
rect 215110 154544 215116 154556
rect 201276 154516 215116 154544
rect 201276 154504 201282 154516
rect 215110 154504 215116 154516
rect 215168 154504 215174 154556
rect 196526 154436 196532 154488
rect 196584 154476 196590 154488
rect 210694 154476 210700 154488
rect 196584 154448 210700 154476
rect 196584 154436 196590 154448
rect 210694 154436 210700 154448
rect 210752 154436 210758 154488
rect 188430 154368 188436 154420
rect 188488 154408 188494 154420
rect 249242 154408 249248 154420
rect 188488 154380 249248 154408
rect 188488 154368 188494 154380
rect 249242 154368 249248 154380
rect 249300 154368 249306 154420
rect 181622 154300 181628 154352
rect 181680 154340 181686 154352
rect 240778 154340 240784 154352
rect 181680 154312 240784 154340
rect 181680 154300 181686 154312
rect 240778 154300 240784 154312
rect 240836 154300 240842 154352
rect 157058 154232 157064 154284
rect 157116 154272 157122 154284
rect 160186 154272 160192 154284
rect 157116 154244 160192 154272
rect 157116 154232 157122 154244
rect 160186 154232 160192 154244
rect 160244 154272 160250 154284
rect 174906 154272 174912 154284
rect 160244 154244 174912 154272
rect 160244 154232 160250 154244
rect 174906 154232 174912 154244
rect 174964 154232 174970 154284
rect 183830 154232 183836 154284
rect 183888 154272 183894 154284
rect 243538 154272 243544 154284
rect 183888 154244 243544 154272
rect 183888 154232 183894 154244
rect 243538 154232 243544 154244
rect 243596 154232 243602 154284
rect 153194 154164 153200 154216
rect 153252 154204 153258 154216
rect 173342 154204 173348 154216
rect 153252 154176 173348 154204
rect 153252 154164 153258 154176
rect 173342 154164 173348 154176
rect 173400 154204 173406 154216
rect 176286 154204 176292 154216
rect 173400 154176 176292 154204
rect 173400 154164 173406 154176
rect 176286 154164 176292 154176
rect 176344 154164 176350 154216
rect 182910 154164 182916 154216
rect 182968 154204 182974 154216
rect 182968 154176 238754 154204
rect 182968 154164 182974 154176
rect 151814 154096 151820 154148
rect 151872 154136 151878 154148
rect 174262 154136 174268 154148
rect 151872 154108 174268 154136
rect 151872 154096 151878 154108
rect 174262 154096 174268 154108
rect 174320 154096 174326 154148
rect 180426 154096 180432 154148
rect 180484 154136 180490 154148
rect 227806 154136 227812 154148
rect 180484 154108 227812 154136
rect 180484 154096 180490 154108
rect 227806 154096 227812 154108
rect 227864 154096 227870 154148
rect 173250 154068 173256 154080
rect 161446 154040 173256 154068
rect 139394 153960 139400 154012
rect 139452 154000 139458 154012
rect 161446 154000 161474 154040
rect 173250 154028 173256 154040
rect 173308 154068 173314 154080
rect 217318 154068 217324 154080
rect 173308 154040 217324 154068
rect 173308 154028 173314 154040
rect 217318 154028 217324 154040
rect 217376 154028 217382 154080
rect 139452 153972 161474 154000
rect 139452 153960 139458 153972
rect 180518 153960 180524 154012
rect 180576 154000 180582 154012
rect 220722 154000 220728 154012
rect 180576 153972 220728 154000
rect 180576 153960 180582 153972
rect 220722 153960 220728 153972
rect 220780 154000 220786 154012
rect 228358 154000 228364 154012
rect 220780 153972 228364 154000
rect 220780 153960 220786 153972
rect 228358 153960 228364 153972
rect 228416 153960 228422 154012
rect 91094 153892 91100 153944
rect 91152 153932 91158 153944
rect 169478 153932 169484 153944
rect 91152 153904 169484 153932
rect 91152 153892 91158 153904
rect 169478 153892 169484 153904
rect 169536 153892 169542 153944
rect 174630 153932 174636 153944
rect 172486 153904 174636 153932
rect 46934 153824 46940 153876
rect 46992 153864 46998 153876
rect 155770 153864 155776 153876
rect 46992 153836 155776 153864
rect 46992 153824 46998 153836
rect 155770 153824 155776 153836
rect 155828 153824 155834 153876
rect 157334 153824 157340 153876
rect 157392 153864 157398 153876
rect 172486 153864 172514 153904
rect 174630 153892 174636 153904
rect 174688 153932 174694 153944
rect 212994 153932 213000 153944
rect 174688 153904 213000 153932
rect 174688 153892 174694 153904
rect 212994 153892 213000 153904
rect 213052 153892 213058 153944
rect 157392 153836 172514 153864
rect 157392 153824 157398 153836
rect 178862 153824 178868 153876
rect 178920 153864 178926 153876
rect 211154 153864 211160 153876
rect 178920 153836 211160 153864
rect 178920 153824 178926 153836
rect 211154 153824 211160 153836
rect 211212 153864 211218 153876
rect 212166 153864 212172 153876
rect 211212 153836 212172 153864
rect 211212 153824 211218 153836
rect 212166 153824 212172 153836
rect 212224 153824 212230 153876
rect 238726 153864 238754 154176
rect 269114 154096 269120 154148
rect 269172 154136 269178 154148
rect 270034 154136 270040 154148
rect 269172 154108 270040 154136
rect 269172 154096 269178 154108
rect 270034 154096 270040 154108
rect 270092 154096 270098 154148
rect 287238 154096 287244 154148
rect 287296 154136 287302 154148
rect 288342 154136 288348 154148
rect 287296 154108 288348 154136
rect 287296 154096 287302 154108
rect 288342 154096 288348 154108
rect 288400 154096 288406 154148
rect 241330 153864 241336 153876
rect 238726 153836 241336 153864
rect 241330 153824 241336 153836
rect 241388 153864 241394 153876
rect 253198 153864 253204 153876
rect 241388 153836 253204 153864
rect 241388 153824 241394 153836
rect 253198 153824 253204 153836
rect 253256 153824 253262 153876
rect 178586 153756 178592 153808
rect 178644 153796 178650 153808
rect 208394 153796 208400 153808
rect 178644 153768 208400 153796
rect 178644 153756 178650 153768
rect 208394 153756 208400 153768
rect 208452 153796 208458 153808
rect 209406 153796 209412 153808
rect 208452 153768 209412 153796
rect 208452 153756 208458 153768
rect 209406 153756 209412 153768
rect 209464 153756 209470 153808
rect 176286 153620 176292 153672
rect 176344 153660 176350 153672
rect 235994 153660 236000 153672
rect 176344 153632 236000 153660
rect 176344 153620 176350 153632
rect 235994 153620 236000 153632
rect 236052 153620 236058 153672
rect 191190 153552 191196 153604
rect 191248 153592 191254 153604
rect 252186 153592 252192 153604
rect 191248 153564 252192 153592
rect 191248 153552 191254 153564
rect 252186 153552 252192 153564
rect 252244 153552 252250 153604
rect 270034 153280 270040 153332
rect 270092 153320 270098 153332
rect 483014 153320 483020 153332
rect 270092 153292 483020 153320
rect 270092 153280 270098 153292
rect 483014 153280 483020 153292
rect 483072 153280 483078 153332
rect 195606 153212 195612 153264
rect 195664 153252 195670 153264
rect 200574 153252 200580 153264
rect 195664 153224 200580 153252
rect 195664 153212 195670 153224
rect 200574 153212 200580 153224
rect 200632 153212 200638 153264
rect 204346 153212 204352 153264
rect 204404 153252 204410 153264
rect 204622 153252 204628 153264
rect 204404 153224 204628 153252
rect 204404 153212 204410 153224
rect 204622 153212 204628 153224
rect 204680 153212 204686 153264
rect 205358 153212 205364 153264
rect 205416 153252 205422 153264
rect 205542 153252 205548 153264
rect 205416 153224 205548 153252
rect 205416 153212 205422 153224
rect 205542 153212 205548 153224
rect 205600 153212 205606 153264
rect 227806 153212 227812 153264
rect 227864 153252 227870 153264
rect 228910 153252 228916 153264
rect 227864 153224 228916 153252
rect 227864 153212 227870 153224
rect 228910 153212 228916 153224
rect 228968 153252 228974 153264
rect 229738 153252 229744 153264
rect 228968 153224 229744 153252
rect 228968 153212 228974 153224
rect 229738 153212 229744 153224
rect 229796 153212 229802 153264
rect 288342 153212 288348 153264
rect 288400 153252 288406 153264
rect 507854 153252 507860 153264
rect 288400 153224 507860 153252
rect 288400 153212 288406 153224
rect 507854 153212 507860 153224
rect 507912 153212 507918 153264
rect 181898 153144 181904 153196
rect 181956 153184 181962 153196
rect 182082 153184 182088 153196
rect 181956 153156 182088 153184
rect 181956 153144 181962 153156
rect 182082 153144 182088 153156
rect 182140 153144 182146 153196
rect 204438 153144 204444 153196
rect 204496 153184 204502 153196
rect 273806 153184 273812 153196
rect 204496 153156 273812 153184
rect 204496 153144 204502 153156
rect 273806 153144 273812 153156
rect 273864 153144 273870 153196
rect 276474 153144 276480 153196
rect 276532 153184 276538 153196
rect 579890 153184 579896 153196
rect 276532 153156 579896 153184
rect 276532 153144 276538 153156
rect 579890 153144 579896 153156
rect 579948 153144 579954 153196
rect 186498 153076 186504 153128
rect 186556 153116 186562 153128
rect 280246 153116 280252 153128
rect 186556 153088 280252 153116
rect 186556 153076 186562 153088
rect 280246 153076 280252 153088
rect 280304 153116 280310 153128
rect 281442 153116 281448 153128
rect 280304 153088 281448 153116
rect 280304 153076 280310 153088
rect 281442 153076 281448 153088
rect 281500 153076 281506 153128
rect 202322 153008 202328 153060
rect 202380 153048 202386 153060
rect 269022 153048 269028 153060
rect 202380 153020 269028 153048
rect 202380 153008 202386 153020
rect 269022 153008 269028 153020
rect 269080 153008 269086 153060
rect 178678 152940 178684 152992
rect 178736 152980 178742 152992
rect 183278 152980 183284 152992
rect 178736 152952 183284 152980
rect 178736 152940 178742 152952
rect 183278 152940 183284 152952
rect 183336 152940 183342 152992
rect 189258 152940 189264 152992
rect 189316 152980 189322 152992
rect 190178 152980 190184 152992
rect 189316 152952 190184 152980
rect 189316 152940 189322 152952
rect 190178 152940 190184 152952
rect 190236 152940 190242 152992
rect 190546 152940 190552 152992
rect 190604 152980 190610 152992
rect 191558 152980 191564 152992
rect 190604 152952 191564 152980
rect 190604 152940 190610 152952
rect 191558 152940 191564 152952
rect 191616 152940 191622 152992
rect 196066 152940 196072 152992
rect 196124 152980 196130 152992
rect 196526 152980 196532 152992
rect 196124 152952 196532 152980
rect 196124 152940 196130 152952
rect 196526 152940 196532 152952
rect 196584 152940 196590 152992
rect 199010 152940 199016 152992
rect 199068 152980 199074 152992
rect 258626 152980 258632 152992
rect 199068 152952 258632 152980
rect 199068 152940 199074 152952
rect 258626 152940 258632 152952
rect 258684 152940 258690 152992
rect 182358 152872 182364 152924
rect 182416 152912 182422 152924
rect 241422 152912 241428 152924
rect 182416 152884 241428 152912
rect 182416 152872 182422 152884
rect 241422 152872 241428 152884
rect 241480 152912 241486 152924
rect 246298 152912 246304 152924
rect 241480 152884 246304 152912
rect 241480 152872 241486 152884
rect 246298 152872 246304 152884
rect 246356 152872 246362 152924
rect 181806 152804 181812 152856
rect 181864 152844 181870 152856
rect 239398 152844 239404 152856
rect 181864 152816 239404 152844
rect 181864 152804 181870 152816
rect 239398 152804 239404 152816
rect 239456 152804 239462 152856
rect 180978 152736 180984 152788
rect 181036 152776 181042 152788
rect 185486 152776 185492 152788
rect 181036 152748 185492 152776
rect 181036 152736 181042 152748
rect 185486 152736 185492 152748
rect 185544 152736 185550 152788
rect 185872 152748 186084 152776
rect 173158 152668 173164 152720
rect 173216 152708 173222 152720
rect 173802 152708 173808 152720
rect 173216 152680 173808 152708
rect 173216 152668 173222 152680
rect 173802 152668 173808 152680
rect 173860 152708 173866 152720
rect 185872 152708 185900 152748
rect 173860 152680 185900 152708
rect 186056 152708 186084 152748
rect 187142 152736 187148 152788
rect 187200 152776 187206 152788
rect 193030 152776 193036 152788
rect 187200 152748 193036 152776
rect 187200 152736 187206 152748
rect 193030 152736 193036 152748
rect 193088 152736 193094 152788
rect 193306 152736 193312 152788
rect 193364 152776 193370 152788
rect 193950 152776 193956 152788
rect 193364 152748 193956 152776
rect 193364 152736 193370 152748
rect 193950 152736 193956 152748
rect 194008 152736 194014 152788
rect 194870 152736 194876 152788
rect 194928 152776 194934 152788
rect 247310 152776 247316 152788
rect 194928 152748 247316 152776
rect 194928 152736 194934 152748
rect 247310 152736 247316 152748
rect 247368 152736 247374 152788
rect 214558 152708 214564 152720
rect 186056 152680 214564 152708
rect 173860 152668 173866 152680
rect 214558 152668 214564 152680
rect 214616 152668 214622 152720
rect 217318 152668 217324 152720
rect 217376 152708 217382 152720
rect 217778 152708 217784 152720
rect 217376 152680 217784 152708
rect 217376 152668 217382 152680
rect 217778 152668 217784 152680
rect 217836 152668 217842 152720
rect 133874 152600 133880 152652
rect 133932 152640 133938 152652
rect 133932 152612 166994 152640
rect 133932 152600 133938 152612
rect 128998 152532 129004 152584
rect 129056 152572 129062 152584
rect 129056 152544 161474 152572
rect 129056 152532 129062 152544
rect 34514 152464 34520 152516
rect 34572 152504 34578 152516
rect 149146 152504 149152 152516
rect 34572 152476 149152 152504
rect 34572 152464 34578 152476
rect 149146 152464 149152 152476
rect 149204 152464 149210 152516
rect 161446 152300 161474 152544
rect 166966 152368 166994 152612
rect 168650 152600 168656 152652
rect 168708 152640 168714 152652
rect 169202 152640 169208 152652
rect 168708 152612 169208 152640
rect 168708 152600 168714 152612
rect 169202 152600 169208 152612
rect 169260 152600 169266 152652
rect 177666 152600 177672 152652
rect 177724 152640 177730 152652
rect 182910 152640 182916 152652
rect 177724 152612 182916 152640
rect 177724 152600 177730 152612
rect 182910 152600 182916 152612
rect 182968 152600 182974 152652
rect 185486 152600 185492 152652
rect 185544 152640 185550 152652
rect 217336 152640 217364 152668
rect 185544 152612 217364 152640
rect 185544 152600 185550 152612
rect 281442 152600 281448 152652
rect 281500 152640 281506 152652
rect 307202 152640 307208 152652
rect 281500 152612 307208 152640
rect 281500 152600 281506 152612
rect 307202 152600 307208 152612
rect 307260 152600 307266 152652
rect 171134 152532 171140 152584
rect 171192 152572 171198 152584
rect 172330 152572 172336 152584
rect 171192 152544 172336 152572
rect 171192 152532 171198 152544
rect 172330 152532 172336 152544
rect 172388 152532 172394 152584
rect 182450 152532 182456 152584
rect 182508 152572 182514 152584
rect 183186 152572 183192 152584
rect 182508 152544 183192 152572
rect 182508 152532 182514 152544
rect 183186 152532 183192 152544
rect 183244 152532 183250 152584
rect 183278 152532 183284 152584
rect 183336 152572 183342 152584
rect 183336 152544 186084 152572
rect 183336 152532 183342 152544
rect 167270 152464 167276 152516
rect 167328 152504 167334 152516
rect 167638 152504 167644 152516
rect 167328 152476 167644 152504
rect 167328 152464 167334 152476
rect 167638 152464 167644 152476
rect 167696 152464 167702 152516
rect 171686 152464 171692 152516
rect 171744 152504 171750 152516
rect 171870 152504 171876 152516
rect 171744 152476 171876 152504
rect 171744 152464 171750 152476
rect 171870 152464 171876 152476
rect 171928 152464 171934 152516
rect 175550 152464 175556 152516
rect 175608 152504 175614 152516
rect 176194 152504 176200 152516
rect 175608 152476 176200 152504
rect 175608 152464 175614 152476
rect 176194 152464 176200 152476
rect 176252 152464 176258 152516
rect 176838 152464 176844 152516
rect 176896 152504 176902 152516
rect 177574 152504 177580 152516
rect 176896 152476 177580 152504
rect 176896 152464 176902 152476
rect 177574 152464 177580 152476
rect 177632 152464 177638 152516
rect 182266 152464 182272 152516
rect 182324 152504 182330 152516
rect 182818 152504 182824 152516
rect 182324 152476 182824 152504
rect 182324 152464 182330 152476
rect 182818 152464 182824 152476
rect 182876 152464 182882 152516
rect 185118 152464 185124 152516
rect 185176 152504 185182 152516
rect 185946 152504 185952 152516
rect 185176 152476 185952 152504
rect 185176 152464 185182 152476
rect 185946 152464 185952 152476
rect 186004 152464 186010 152516
rect 186056 152504 186084 152544
rect 186590 152532 186596 152584
rect 186648 152572 186654 152584
rect 187050 152572 187056 152584
rect 186648 152544 187056 152572
rect 186648 152532 186654 152544
rect 187050 152532 187056 152544
rect 187108 152532 187114 152584
rect 187694 152532 187700 152584
rect 187752 152572 187758 152584
rect 188706 152572 188712 152584
rect 187752 152544 188712 152572
rect 187752 152532 187758 152544
rect 188706 152532 188712 152544
rect 188764 152532 188770 152584
rect 189166 152532 189172 152584
rect 189224 152572 189230 152584
rect 189810 152572 189816 152584
rect 189224 152544 189816 152572
rect 189224 152532 189230 152544
rect 189810 152532 189816 152544
rect 189868 152532 189874 152584
rect 190546 152532 190552 152584
rect 190604 152572 190610 152584
rect 191466 152572 191472 152584
rect 190604 152544 191472 152572
rect 190604 152532 190610 152544
rect 191466 152532 191472 152544
rect 191524 152532 191530 152584
rect 191926 152532 191932 152584
rect 191984 152572 191990 152584
rect 192570 152572 192576 152584
rect 191984 152544 192576 152572
rect 191984 152532 191990 152544
rect 192570 152532 192576 152544
rect 192628 152532 192634 152584
rect 193214 152532 193220 152584
rect 193272 152572 193278 152584
rect 194226 152572 194232 152584
rect 193272 152544 194232 152572
rect 193272 152532 193278 152544
rect 194226 152532 194232 152544
rect 194284 152532 194290 152584
rect 194686 152532 194692 152584
rect 194744 152572 194750 152584
rect 195054 152572 195060 152584
rect 194744 152544 195060 152572
rect 194744 152532 194750 152544
rect 195054 152532 195060 152544
rect 195112 152532 195118 152584
rect 195146 152532 195152 152584
rect 195204 152572 195210 152584
rect 212902 152572 212908 152584
rect 195204 152544 212908 152572
rect 195204 152532 195210 152544
rect 212902 152532 212908 152544
rect 212960 152532 212966 152584
rect 269022 152532 269028 152584
rect 269080 152572 269086 152584
rect 511994 152572 512000 152584
rect 269080 152544 512000 152572
rect 269080 152532 269086 152544
rect 511994 152532 512000 152544
rect 512052 152532 512058 152584
rect 209866 152504 209872 152516
rect 186056 152476 209872 152504
rect 209866 152464 209872 152476
rect 209924 152464 209930 152516
rect 273806 152464 273812 152516
rect 273864 152504 273870 152516
rect 274542 152504 274548 152516
rect 273864 152476 274548 152504
rect 273864 152464 273870 152476
rect 274542 152464 274548 152476
rect 274600 152504 274606 152516
rect 536098 152504 536104 152516
rect 274600 152476 536104 152504
rect 274600 152464 274606 152476
rect 536098 152464 536104 152476
rect 536156 152464 536162 152516
rect 167454 152396 167460 152448
rect 167512 152436 167518 152448
rect 167914 152436 167920 152448
rect 167512 152408 167920 152436
rect 167512 152396 167518 152408
rect 167914 152396 167920 152408
rect 167972 152396 167978 152448
rect 168374 152396 168380 152448
rect 168432 152436 168438 152448
rect 169110 152436 169116 152448
rect 168432 152408 169116 152436
rect 168432 152396 168438 152408
rect 169110 152396 169116 152408
rect 169168 152396 169174 152448
rect 172974 152396 172980 152448
rect 173032 152436 173038 152448
rect 173618 152436 173624 152448
rect 173032 152408 173624 152436
rect 173032 152396 173038 152408
rect 173618 152396 173624 152408
rect 173676 152396 173682 152448
rect 175458 152396 175464 152448
rect 175516 152436 175522 152448
rect 176470 152436 176476 152448
rect 175516 152408 176476 152436
rect 175516 152396 175522 152408
rect 176470 152396 176476 152408
rect 176528 152396 176534 152448
rect 220078 152436 220084 152448
rect 176626 152408 220084 152436
rect 172790 152368 172796 152380
rect 166966 152340 172796 152368
rect 172790 152328 172796 152340
rect 172848 152368 172854 152380
rect 176626 152368 176654 152408
rect 220078 152396 220084 152408
rect 220136 152396 220142 152448
rect 172848 152340 176654 152368
rect 172848 152328 172854 152340
rect 181162 152328 181168 152380
rect 181220 152368 181226 152380
rect 181990 152368 181996 152380
rect 181220 152340 181996 152368
rect 181220 152328 181226 152340
rect 181990 152328 181996 152340
rect 182048 152328 182054 152380
rect 182358 152328 182364 152380
rect 182416 152368 182422 152380
rect 183462 152368 183468 152380
rect 182416 152340 183468 152368
rect 182416 152328 182422 152340
rect 183462 152328 183468 152340
rect 183520 152328 183526 152380
rect 185302 152328 185308 152380
rect 185360 152368 185366 152380
rect 186130 152368 186136 152380
rect 185360 152340 186136 152368
rect 185360 152328 185366 152340
rect 186130 152328 186136 152340
rect 186188 152328 186194 152380
rect 186498 152328 186504 152380
rect 186556 152368 186562 152380
rect 187326 152368 187332 152380
rect 186556 152340 187332 152368
rect 186556 152328 186562 152340
rect 187326 152328 187332 152340
rect 187384 152328 187390 152380
rect 188338 152328 188344 152380
rect 188396 152368 188402 152380
rect 188890 152368 188896 152380
rect 188396 152340 188896 152368
rect 188396 152328 188402 152340
rect 188890 152328 188896 152340
rect 188948 152328 188954 152380
rect 192018 152328 192024 152380
rect 192076 152368 192082 152380
rect 192846 152368 192852 152380
rect 192076 152340 192852 152368
rect 192076 152328 192082 152340
rect 192846 152328 192852 152340
rect 192904 152328 192910 152380
rect 193030 152328 193036 152380
rect 193088 152368 193094 152380
rect 210602 152368 210608 152380
rect 193088 152340 210608 152368
rect 193088 152328 193094 152340
rect 210602 152328 210608 152340
rect 210660 152328 210666 152380
rect 172238 152300 172244 152312
rect 161446 152272 172244 152300
rect 172238 152260 172244 152272
rect 172296 152300 172302 152312
rect 210510 152300 210516 152312
rect 172296 152272 210516 152300
rect 172296 152260 172302 152272
rect 210510 152260 210516 152272
rect 210568 152260 210574 152312
rect 185026 152192 185032 152244
rect 185084 152232 185090 152244
rect 186222 152232 186228 152244
rect 185084 152204 186228 152232
rect 185084 152192 185090 152204
rect 186222 152192 186228 152204
rect 186280 152192 186286 152244
rect 186406 152192 186412 152244
rect 186464 152232 186470 152244
rect 187602 152232 187608 152244
rect 186464 152204 187608 152232
rect 186464 152192 186470 152204
rect 187602 152192 187608 152204
rect 187660 152192 187666 152244
rect 191834 152192 191840 152244
rect 191892 152232 191898 152244
rect 192938 152232 192944 152244
rect 191892 152204 192944 152232
rect 191892 152192 191898 152204
rect 192938 152192 192944 152204
rect 192996 152192 193002 152244
rect 194962 152192 194968 152244
rect 195020 152232 195026 152244
rect 195882 152232 195888 152244
rect 195020 152204 195888 152232
rect 195020 152192 195026 152204
rect 195882 152192 195888 152204
rect 195940 152192 195946 152244
rect 196066 152192 196072 152244
rect 196124 152232 196130 152244
rect 196710 152232 196716 152244
rect 196124 152204 196716 152232
rect 196124 152192 196130 152204
rect 196710 152192 196716 152204
rect 196768 152192 196774 152244
rect 197354 152192 197360 152244
rect 197412 152232 197418 152244
rect 198090 152232 198096 152244
rect 197412 152204 198096 152232
rect 197412 152192 197418 152204
rect 198090 152192 198096 152204
rect 198148 152192 198154 152244
rect 198826 152192 198832 152244
rect 198884 152232 198890 152244
rect 199930 152232 199936 152244
rect 198884 152204 199936 152232
rect 198884 152192 198890 152204
rect 199930 152192 199936 152204
rect 199988 152192 199994 152244
rect 200206 152192 200212 152244
rect 200264 152232 200270 152244
rect 200758 152232 200764 152244
rect 200264 152204 200764 152232
rect 200264 152192 200270 152204
rect 200758 152192 200764 152204
rect 200816 152192 200822 152244
rect 201678 152192 201684 152244
rect 201736 152232 201742 152244
rect 202506 152232 202512 152244
rect 201736 152204 202512 152232
rect 201736 152192 201742 152204
rect 202506 152192 202512 152204
rect 202564 152192 202570 152244
rect 203334 152192 203340 152244
rect 203392 152232 203398 152244
rect 203794 152232 203800 152244
rect 203392 152204 203800 152232
rect 203392 152192 203398 152204
rect 203794 152192 203800 152204
rect 203852 152192 203858 152244
rect 204806 152192 204812 152244
rect 204864 152232 204870 152244
rect 205450 152232 205456 152244
rect 204864 152204 205456 152232
rect 204864 152192 204870 152204
rect 205450 152192 205456 152204
rect 205508 152192 205514 152244
rect 188890 152124 188896 152176
rect 188948 152164 188954 152176
rect 195146 152164 195152 152176
rect 188948 152136 195152 152164
rect 188948 152124 188954 152136
rect 195146 152124 195152 152136
rect 195204 152124 195210 152176
rect 196250 152124 196256 152176
rect 196308 152164 196314 152176
rect 196894 152164 196900 152176
rect 196308 152136 196900 152164
rect 196308 152124 196314 152136
rect 196894 152124 196900 152136
rect 196952 152124 196958 152176
rect 197446 152124 197452 152176
rect 197504 152164 197510 152176
rect 198550 152164 198556 152176
rect 197504 152136 198556 152164
rect 197504 152124 197510 152136
rect 198550 152124 198556 152136
rect 198608 152124 198614 152176
rect 202874 152124 202880 152176
rect 202932 152164 202938 152176
rect 203886 152164 203892 152176
rect 202932 152136 203892 152164
rect 202932 152124 202938 152136
rect 203886 152124 203892 152136
rect 203944 152124 203950 152176
rect 165982 151852 165988 151904
rect 166040 151892 166046 151904
rect 166258 151892 166264 151904
rect 166040 151864 166264 151892
rect 166040 151852 166046 151864
rect 166258 151852 166264 151864
rect 166316 151852 166322 151904
rect 176654 151716 176660 151768
rect 176712 151756 176718 151768
rect 181530 151756 181536 151768
rect 176712 151728 181536 151756
rect 176712 151716 176718 151728
rect 181530 151716 181536 151728
rect 181588 151716 181594 151768
rect 189626 151716 189632 151768
rect 189684 151756 189690 151768
rect 190086 151756 190092 151768
rect 189684 151728 190092 151756
rect 189684 151716 189690 151728
rect 190086 151716 190092 151728
rect 190144 151716 190150 151768
rect 203058 151716 203064 151768
rect 203116 151756 203122 151768
rect 280154 151756 280160 151768
rect 203116 151728 280160 151756
rect 203116 151716 203122 151728
rect 280154 151716 280160 151728
rect 280212 151716 280218 151768
rect 182634 151648 182640 151700
rect 182692 151688 182698 151700
rect 244918 151688 244924 151700
rect 182692 151660 244924 151688
rect 182692 151648 182698 151660
rect 244918 151648 244924 151660
rect 244976 151648 244982 151700
rect 174538 151580 174544 151632
rect 174596 151620 174602 151632
rect 175642 151620 175648 151632
rect 174596 151592 175648 151620
rect 174596 151580 174602 151592
rect 175642 151580 175648 151592
rect 175700 151620 175706 151632
rect 235534 151620 235540 151632
rect 175700 151592 235540 151620
rect 175700 151580 175706 151592
rect 235534 151580 235540 151592
rect 235592 151580 235598 151632
rect 185670 151512 185676 151564
rect 185728 151552 185734 151564
rect 242802 151552 242808 151564
rect 185728 151524 242808 151552
rect 185728 151512 185734 151524
rect 242802 151512 242808 151524
rect 242860 151512 242866 151564
rect 181070 151444 181076 151496
rect 181128 151484 181134 151496
rect 236638 151484 236644 151496
rect 181128 151456 236644 151484
rect 181128 151444 181134 151456
rect 236638 151444 236644 151456
rect 236696 151444 236702 151496
rect 181254 151376 181260 151428
rect 181312 151416 181318 151428
rect 232498 151416 232504 151428
rect 181312 151388 232504 151416
rect 181312 151376 181318 151388
rect 232498 151376 232504 151388
rect 232556 151376 232562 151428
rect 180242 151308 180248 151360
rect 180300 151348 180306 151360
rect 229094 151348 229100 151360
rect 180300 151320 229100 151348
rect 180300 151308 180306 151320
rect 229094 151308 229100 151320
rect 229152 151348 229158 151360
rect 230014 151348 230020 151360
rect 229152 151320 230020 151348
rect 229152 151308 229158 151320
rect 230014 151308 230020 151320
rect 230072 151308 230078 151360
rect 140774 151240 140780 151292
rect 140832 151280 140838 151292
rect 158438 151280 158444 151292
rect 140832 151252 158444 151280
rect 140832 151240 140838 151252
rect 158438 151240 158444 151252
rect 158496 151240 158502 151292
rect 184934 151240 184940 151292
rect 184992 151280 184998 151292
rect 233970 151280 233976 151292
rect 184992 151252 233976 151280
rect 184992 151240 184998 151252
rect 233970 151240 233976 151252
rect 234028 151240 234034 151292
rect 82814 151172 82820 151224
rect 82872 151212 82878 151224
rect 152826 151212 152832 151224
rect 82872 151184 152832 151212
rect 82872 151172 82878 151184
rect 152826 151172 152832 151184
rect 152884 151172 152890 151224
rect 189074 151172 189080 151224
rect 189132 151212 189138 151224
rect 189534 151212 189540 151224
rect 189132 151184 189540 151212
rect 189132 151172 189138 151184
rect 189534 151172 189540 151184
rect 189592 151172 189598 151224
rect 192202 151172 192208 151224
rect 192260 151212 192266 151224
rect 240870 151212 240876 151224
rect 192260 151184 240876 151212
rect 192260 151172 192266 151184
rect 240870 151172 240876 151184
rect 240928 151172 240934 151224
rect 64874 151104 64880 151156
rect 64932 151144 64938 151156
rect 155494 151144 155500 151156
rect 64932 151116 155500 151144
rect 64932 151104 64938 151116
rect 155494 151104 155500 151116
rect 155552 151104 155558 151156
rect 189442 151104 189448 151156
rect 189500 151144 189506 151156
rect 189994 151144 190000 151156
rect 189500 151116 190000 151144
rect 189500 151104 189506 151116
rect 189994 151104 190000 151116
rect 190052 151104 190058 151156
rect 197998 151104 198004 151156
rect 198056 151144 198062 151156
rect 242986 151144 242992 151156
rect 198056 151116 242992 151144
rect 198056 151104 198062 151116
rect 242986 151104 242992 151116
rect 243044 151104 243050 151156
rect 28994 151036 29000 151088
rect 29052 151076 29058 151088
rect 164510 151076 164516 151088
rect 29052 151048 164516 151076
rect 29052 151036 29058 151048
rect 164510 151036 164516 151048
rect 164568 151036 164574 151088
rect 189074 151036 189080 151088
rect 189132 151076 189138 151088
rect 190362 151076 190368 151088
rect 189132 151048 190368 151076
rect 189132 151036 189138 151048
rect 190362 151036 190368 151048
rect 190420 151036 190426 151088
rect 197078 151036 197084 151088
rect 197136 151076 197142 151088
rect 235994 151076 236000 151088
rect 197136 151048 236000 151076
rect 197136 151036 197142 151048
rect 235994 151036 236000 151048
rect 236052 151036 236058 151088
rect 242802 151036 242808 151088
rect 242860 151076 242866 151088
rect 295978 151076 295984 151088
rect 242860 151048 295984 151076
rect 242860 151036 242866 151048
rect 295978 151036 295984 151048
rect 296036 151036 296042 151088
rect 195514 150968 195520 151020
rect 195572 151008 195578 151020
rect 233234 151008 233240 151020
rect 195572 150980 233240 151008
rect 195572 150968 195578 150980
rect 233234 150968 233240 150980
rect 233292 150968 233298 151020
rect 199654 150900 199660 150952
rect 199712 150940 199718 150952
rect 223206 150940 223212 150952
rect 199712 150912 223212 150940
rect 199712 150900 199718 150912
rect 223206 150900 223212 150912
rect 223264 150900 223270 150952
rect 190086 150832 190092 150884
rect 190144 150872 190150 150884
rect 211614 150872 211620 150884
rect 190144 150844 211620 150872
rect 190144 150832 190150 150844
rect 211614 150832 211620 150844
rect 211672 150832 211678 150884
rect 233234 150492 233240 150544
rect 233292 150532 233298 150544
rect 234246 150532 234252 150544
rect 233292 150504 234252 150532
rect 233292 150492 233298 150504
rect 234246 150492 234252 150504
rect 234304 150492 234310 150544
rect 235994 150424 236000 150476
rect 236052 150464 236058 150476
rect 236914 150464 236920 150476
rect 236052 150436 236920 150464
rect 236052 150424 236058 150436
rect 236914 150424 236920 150436
rect 236972 150424 236978 150476
rect 244918 150424 244924 150476
rect 244976 150464 244982 150476
rect 250438 150464 250444 150476
rect 244976 150436 250444 150464
rect 244976 150424 244982 150436
rect 250438 150424 250444 150436
rect 250496 150424 250502 150476
rect 280154 150424 280160 150476
rect 280212 150464 280218 150476
rect 280798 150464 280804 150476
rect 280212 150436 280804 150464
rect 280212 150424 280218 150436
rect 280798 150424 280804 150436
rect 280856 150424 280862 150476
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 11698 150396 11704 150408
rect 3384 150368 11704 150396
rect 3384 150356 3390 150368
rect 11698 150356 11704 150368
rect 11756 150356 11762 150408
rect 186682 150356 186688 150408
rect 186740 150396 186746 150408
rect 215938 150396 215944 150408
rect 186740 150368 215944 150396
rect 186740 150356 186746 150368
rect 215938 150356 215944 150368
rect 215996 150356 216002 150408
rect 204254 150288 204260 150340
rect 204312 150328 204318 150340
rect 291286 150328 291292 150340
rect 204312 150300 291292 150328
rect 204312 150288 204318 150300
rect 291286 150288 291292 150300
rect 291344 150288 291350 150340
rect 187786 150220 187792 150272
rect 187844 150260 187850 150272
rect 272518 150260 272524 150272
rect 187844 150232 272524 150260
rect 187844 150220 187850 150232
rect 272518 150220 272524 150232
rect 272576 150220 272582 150272
rect 187418 150152 187424 150204
rect 187476 150192 187482 150204
rect 259454 150192 259460 150204
rect 187476 150164 259460 150192
rect 187476 150152 187482 150164
rect 259454 150152 259460 150164
rect 259512 150152 259518 150204
rect 174998 150084 175004 150136
rect 175056 150124 175062 150136
rect 235442 150124 235448 150136
rect 175056 150096 235448 150124
rect 175056 150084 175062 150096
rect 235442 150084 235448 150096
rect 235500 150084 235506 150136
rect 197630 150016 197636 150068
rect 197688 150056 197694 150068
rect 257430 150056 257436 150068
rect 197688 150028 257436 150056
rect 197688 150016 197694 150028
rect 257430 150016 257436 150028
rect 257488 150016 257494 150068
rect 196618 149948 196624 150000
rect 196676 149988 196682 150000
rect 252094 149988 252100 150000
rect 196676 149960 252100 149988
rect 196676 149948 196682 149960
rect 252094 149948 252100 149960
rect 252152 149948 252158 150000
rect 181622 149880 181628 149932
rect 181680 149920 181686 149932
rect 235258 149920 235264 149932
rect 181680 149892 235264 149920
rect 181680 149880 181686 149892
rect 235258 149880 235264 149892
rect 235316 149880 235322 149932
rect 177482 149812 177488 149864
rect 177540 149852 177546 149864
rect 218698 149852 218704 149864
rect 177540 149824 218704 149852
rect 177540 149812 177546 149824
rect 218698 149812 218704 149824
rect 218756 149812 218762 149864
rect 56594 149744 56600 149796
rect 56652 149784 56658 149796
rect 165706 149784 165712 149796
rect 56652 149756 165712 149784
rect 56652 149744 56658 149756
rect 165706 149744 165712 149756
rect 165764 149744 165770 149796
rect 179138 149744 179144 149796
rect 179196 149784 179202 149796
rect 213730 149784 213736 149796
rect 179196 149756 213736 149784
rect 179196 149744 179202 149756
rect 213730 149744 213736 149756
rect 213788 149744 213794 149796
rect 215938 149744 215944 149796
rect 215996 149784 216002 149796
rect 234062 149784 234068 149796
rect 215996 149756 234068 149784
rect 215996 149744 216002 149756
rect 234062 149744 234068 149756
rect 234120 149744 234126 149796
rect 272518 149744 272524 149796
rect 272576 149784 272582 149796
rect 327074 149784 327080 149796
rect 272576 149756 327080 149784
rect 272576 149744 272582 149756
rect 327074 149744 327080 149756
rect 327132 149744 327138 149796
rect 15194 149676 15200 149728
rect 15252 149716 15258 149728
rect 163130 149716 163136 149728
rect 15252 149688 163136 149716
rect 15252 149676 15258 149688
rect 163130 149676 163136 149688
rect 163188 149676 163194 149728
rect 186682 149676 186688 149728
rect 186740 149716 186746 149728
rect 186958 149716 186964 149728
rect 186740 149688 186964 149716
rect 186740 149676 186746 149688
rect 186958 149676 186964 149688
rect 187016 149676 187022 149728
rect 201954 149676 201960 149728
rect 202012 149716 202018 149728
rect 232866 149716 232872 149728
rect 202012 149688 232872 149716
rect 202012 149676 202018 149688
rect 232866 149676 232872 149688
rect 232924 149676 232930 149728
rect 291286 149676 291292 149728
rect 291344 149716 291350 149728
rect 451274 149716 451280 149728
rect 291344 149688 451280 149716
rect 291344 149676 291350 149688
rect 451274 149676 451280 149688
rect 451332 149676 451338 149728
rect 188522 149608 188528 149660
rect 188580 149648 188586 149660
rect 217502 149648 217508 149660
rect 188580 149620 217508 149648
rect 188580 149608 188586 149620
rect 217502 149608 217508 149620
rect 217560 149608 217566 149660
rect 184014 149540 184020 149592
rect 184072 149580 184078 149592
rect 274818 149580 274824 149592
rect 184072 149552 274824 149580
rect 184072 149540 184078 149552
rect 274818 149540 274824 149552
rect 274876 149540 274882 149592
rect 172514 149472 172520 149524
rect 172572 149512 172578 149524
rect 175826 149512 175832 149524
rect 172572 149484 175832 149512
rect 172572 149472 172578 149484
rect 175826 149472 175832 149484
rect 175884 149512 175890 149524
rect 214006 149512 214012 149524
rect 175884 149484 214012 149512
rect 175884 149472 175890 149484
rect 214006 149472 214012 149484
rect 214064 149472 214070 149524
rect 187786 149268 187792 149320
rect 187844 149308 187850 149320
rect 188982 149308 188988 149320
rect 187844 149280 188988 149308
rect 187844 149268 187850 149280
rect 188982 149268 188988 149280
rect 189040 149268 189046 149320
rect 213730 149064 213736 149116
rect 213788 149104 213794 149116
rect 214558 149104 214564 149116
rect 213788 149076 214564 149104
rect 213788 149064 213794 149076
rect 214558 149064 214564 149076
rect 214616 149064 214622 149116
rect 259454 149064 259460 149116
rect 259512 149104 259518 149116
rect 260098 149104 260104 149116
rect 259512 149076 260104 149104
rect 259512 149064 259518 149076
rect 260098 149064 260104 149076
rect 260156 149064 260162 149116
rect 274818 149064 274824 149116
rect 274876 149104 274882 149116
rect 275278 149104 275284 149116
rect 274876 149076 275284 149104
rect 274876 149064 274882 149076
rect 275278 149064 275284 149076
rect 275336 149064 275342 149116
rect 181898 148996 181904 149048
rect 181956 149036 181962 149048
rect 217134 149036 217140 149048
rect 181956 149008 217140 149036
rect 181956 148996 181962 149008
rect 217134 148996 217140 149008
rect 217192 149036 217198 149048
rect 220078 149036 220084 149048
rect 217192 149008 220084 149036
rect 217192 148996 217198 149008
rect 220078 148996 220084 149008
rect 220136 148996 220142 149048
rect 183554 148928 183560 148980
rect 183612 148968 183618 148980
rect 271874 148968 271880 148980
rect 183612 148940 271880 148968
rect 183612 148928 183618 148940
rect 271874 148928 271880 148940
rect 271932 148928 271938 148980
rect 186038 148860 186044 148912
rect 186096 148900 186102 148912
rect 267826 148900 267832 148912
rect 186096 148872 267832 148900
rect 186096 148860 186102 148872
rect 267826 148860 267832 148872
rect 267884 148900 267890 148912
rect 268378 148900 268384 148912
rect 267884 148872 268384 148900
rect 267884 148860 267890 148872
rect 268378 148860 268384 148872
rect 268436 148860 268442 148912
rect 182174 148792 182180 148844
rect 182232 148832 182238 148844
rect 243722 148832 243728 148844
rect 182232 148804 243728 148832
rect 182232 148792 182238 148804
rect 243722 148792 243728 148804
rect 243780 148792 243786 148844
rect 184290 148724 184296 148776
rect 184348 148764 184354 148776
rect 244090 148764 244096 148776
rect 184348 148736 244096 148764
rect 184348 148724 184354 148736
rect 244090 148724 244096 148736
rect 244148 148724 244154 148776
rect 182174 148656 182180 148708
rect 182232 148696 182238 148708
rect 182542 148696 182548 148708
rect 182232 148668 182548 148696
rect 182232 148656 182238 148668
rect 182542 148656 182548 148668
rect 182600 148656 182606 148708
rect 184474 148656 184480 148708
rect 184532 148696 184538 148708
rect 243630 148696 243636 148708
rect 184532 148668 243636 148696
rect 184532 148656 184538 148668
rect 243630 148656 243636 148668
rect 243688 148656 243694 148708
rect 194134 148588 194140 148640
rect 194192 148628 194198 148640
rect 252002 148628 252008 148640
rect 194192 148600 252008 148628
rect 194192 148588 194198 148600
rect 252002 148588 252008 148600
rect 252060 148588 252066 148640
rect 191650 148520 191656 148572
rect 191708 148560 191714 148572
rect 246390 148560 246396 148572
rect 191708 148532 246396 148560
rect 191708 148520 191714 148532
rect 246390 148520 246396 148532
rect 246448 148520 246454 148572
rect 189718 148452 189724 148504
rect 189776 148492 189782 148504
rect 244274 148492 244280 148504
rect 189776 148464 244280 148492
rect 189776 148452 189782 148464
rect 244274 148452 244280 148464
rect 244332 148452 244338 148504
rect 271874 148452 271880 148504
rect 271932 148492 271938 148504
rect 272426 148492 272432 148504
rect 271932 148464 272432 148492
rect 271932 148452 271938 148464
rect 272426 148452 272432 148464
rect 272484 148452 272490 148504
rect 144914 148384 144920 148436
rect 144972 148424 144978 148436
rect 173710 148424 173716 148436
rect 144972 148396 173716 148424
rect 144972 148384 144978 148396
rect 173710 148384 173716 148396
rect 173768 148384 173774 148436
rect 202230 148384 202236 148436
rect 202288 148424 202294 148436
rect 256050 148424 256056 148436
rect 202288 148396 256056 148424
rect 202288 148384 202294 148396
rect 256050 148384 256056 148396
rect 256108 148384 256114 148436
rect 57974 148316 57980 148368
rect 58032 148356 58038 148368
rect 165890 148356 165896 148368
rect 58032 148328 165896 148356
rect 58032 148316 58038 148328
rect 165890 148316 165896 148328
rect 165948 148316 165954 148368
rect 192662 148316 192668 148368
rect 192720 148356 192726 148368
rect 237006 148356 237012 148368
rect 192720 148328 237012 148356
rect 192720 148316 192726 148328
rect 237006 148316 237012 148328
rect 237064 148316 237070 148368
rect 244090 148316 244096 148368
rect 244148 148356 244154 148368
rect 278038 148356 278044 148368
rect 244148 148328 278044 148356
rect 244148 148316 244154 148328
rect 278038 148316 278044 148328
rect 278096 148316 278102 148368
rect 345014 148356 345020 148368
rect 287026 148328 345020 148356
rect 191558 148248 191564 148300
rect 191616 148288 191622 148300
rect 230198 148288 230204 148300
rect 191616 148260 230204 148288
rect 191616 148248 191622 148260
rect 230198 148248 230204 148260
rect 230256 148248 230262 148300
rect 179506 148180 179512 148232
rect 179564 148220 179570 148232
rect 215294 148220 215300 148232
rect 179564 148192 215300 148220
rect 179564 148180 179570 148192
rect 215294 148180 215300 148192
rect 215352 148180 215358 148232
rect 190178 148112 190184 148164
rect 190236 148152 190242 148164
rect 278406 148152 278412 148164
rect 190236 148124 278412 148152
rect 190236 148112 190242 148124
rect 278406 148112 278412 148124
rect 278464 148152 278470 148164
rect 287026 148152 287054 148328
rect 345014 148316 345020 148328
rect 345072 148316 345078 148368
rect 278464 148124 287054 148152
rect 278464 148112 278470 148124
rect 244274 147636 244280 147688
rect 244332 147676 244338 147688
rect 244918 147676 244924 147688
rect 244332 147648 244924 147676
rect 244332 147636 244338 147648
rect 244918 147636 244924 147648
rect 244976 147636 244982 147688
rect 200850 147568 200856 147620
rect 200908 147608 200914 147620
rect 228542 147608 228548 147620
rect 200908 147580 228548 147608
rect 200908 147568 200914 147580
rect 228542 147568 228548 147580
rect 228600 147568 228606 147620
rect 201770 147500 201776 147552
rect 201828 147540 201834 147552
rect 287238 147540 287244 147552
rect 201828 147512 287244 147540
rect 201828 147500 201834 147512
rect 287238 147500 287244 147512
rect 287296 147500 287302 147552
rect 194778 147432 194784 147484
rect 194836 147472 194842 147484
rect 278958 147472 278964 147484
rect 194836 147444 278964 147472
rect 194836 147432 194842 147444
rect 278958 147432 278964 147444
rect 279016 147472 279022 147484
rect 279970 147472 279976 147484
rect 279016 147444 279976 147472
rect 279016 147432 279022 147444
rect 279970 147432 279976 147444
rect 280028 147432 280034 147484
rect 182450 147364 182456 147416
rect 182508 147404 182514 147416
rect 260190 147404 260196 147416
rect 182508 147376 260196 147404
rect 182508 147364 182514 147376
rect 260190 147364 260196 147376
rect 260248 147404 260254 147416
rect 264238 147404 264244 147416
rect 260248 147376 264244 147404
rect 260248 147364 260254 147376
rect 264238 147364 264244 147376
rect 264296 147364 264302 147416
rect 168374 147296 168380 147348
rect 168432 147336 168438 147348
rect 168558 147336 168564 147348
rect 168432 147308 168564 147336
rect 168432 147296 168438 147308
rect 168558 147296 168564 147308
rect 168616 147296 168622 147348
rect 184750 147296 184756 147348
rect 184808 147336 184814 147348
rect 245194 147336 245200 147348
rect 184808 147308 245200 147336
rect 184808 147296 184814 147308
rect 245194 147296 245200 147308
rect 245252 147296 245258 147348
rect 185302 147228 185308 147280
rect 185360 147268 185366 147280
rect 246574 147268 246580 147280
rect 185360 147240 246580 147268
rect 185360 147228 185366 147240
rect 246574 147228 246580 147240
rect 246632 147228 246638 147280
rect 190730 147160 190736 147212
rect 190788 147200 190794 147212
rect 251910 147200 251916 147212
rect 190788 147172 251916 147200
rect 190788 147160 190794 147172
rect 251910 147160 251916 147172
rect 251968 147160 251974 147212
rect 188062 147092 188068 147144
rect 188120 147132 188126 147144
rect 247678 147132 247684 147144
rect 188120 147104 247684 147132
rect 188120 147092 188126 147104
rect 247678 147092 247684 147104
rect 247736 147092 247742 147144
rect 153838 147024 153844 147076
rect 153896 147064 153902 147076
rect 175090 147064 175096 147076
rect 153896 147036 175096 147064
rect 153896 147024 153902 147036
rect 175090 147024 175096 147036
rect 175148 147024 175154 147076
rect 196342 147024 196348 147076
rect 196400 147064 196406 147076
rect 255406 147064 255412 147076
rect 196400 147036 255412 147064
rect 196400 147024 196406 147036
rect 255406 147024 255412 147036
rect 255464 147024 255470 147076
rect 126238 146956 126244 147008
rect 126296 146996 126302 147008
rect 161750 146996 161756 147008
rect 126296 146968 161756 146996
rect 126296 146956 126302 146968
rect 161750 146956 161756 146968
rect 161808 146956 161814 147008
rect 191098 146956 191104 147008
rect 191156 146996 191162 147008
rect 250530 146996 250536 147008
rect 191156 146968 250536 146996
rect 191156 146956 191162 146968
rect 250530 146956 250536 146968
rect 250588 146956 250594 147008
rect 316678 146996 316684 147008
rect 277366 146968 316684 146996
rect 104894 146888 104900 146940
rect 104952 146928 104958 146940
rect 170950 146928 170956 146940
rect 104952 146900 170956 146928
rect 104952 146888 104958 146900
rect 170950 146888 170956 146900
rect 171008 146888 171014 146940
rect 189534 146888 189540 146940
rect 189592 146928 189598 146940
rect 235810 146928 235816 146940
rect 189592 146900 235816 146928
rect 189592 146888 189598 146900
rect 235810 146888 235816 146900
rect 235868 146888 235874 146940
rect 179690 146820 179696 146872
rect 179748 146860 179754 146872
rect 222194 146860 222200 146872
rect 179748 146832 222200 146860
rect 179748 146820 179754 146832
rect 222194 146820 222200 146832
rect 222252 146860 222258 146872
rect 223022 146860 223028 146872
rect 222252 146832 223028 146860
rect 222252 146820 222258 146832
rect 223022 146820 223028 146832
rect 223080 146820 223086 146872
rect 215294 146752 215300 146804
rect 215352 146792 215358 146804
rect 216582 146792 216588 146804
rect 215352 146764 216588 146792
rect 215352 146752 215358 146764
rect 216582 146752 216588 146764
rect 216640 146792 216646 146804
rect 239582 146792 239588 146804
rect 216640 146764 239588 146792
rect 216640 146752 216646 146764
rect 239582 146752 239588 146764
rect 239640 146752 239646 146804
rect 187970 146684 187976 146736
rect 188028 146724 188034 146736
rect 276198 146724 276204 146736
rect 188028 146696 276204 146724
rect 188028 146684 188034 146696
rect 276198 146684 276204 146696
rect 276256 146724 276262 146736
rect 277366 146724 277394 146968
rect 316678 146956 316684 146968
rect 316736 146956 316742 147008
rect 279970 146888 279976 146940
rect 280028 146928 280034 146940
rect 415394 146928 415400 146940
rect 280028 146900 415400 146928
rect 280028 146888 280034 146900
rect 415394 146888 415400 146900
rect 415452 146888 415458 146940
rect 276256 146696 277394 146724
rect 276256 146684 276262 146696
rect 177390 146276 177396 146328
rect 177448 146316 177454 146328
rect 180058 146316 180064 146328
rect 177448 146288 180064 146316
rect 177448 146276 177454 146288
rect 180058 146276 180064 146288
rect 180116 146276 180122 146328
rect 201678 146208 201684 146260
rect 201736 146248 201742 146260
rect 294046 146248 294052 146260
rect 201736 146220 294052 146248
rect 201736 146208 201742 146220
rect 294046 146208 294052 146220
rect 294104 146248 294110 146260
rect 294874 146248 294880 146260
rect 294104 146220 294880 146248
rect 294104 146208 294110 146220
rect 294874 146208 294880 146220
rect 294932 146208 294938 146260
rect 183646 146140 183652 146192
rect 183704 146180 183710 146192
rect 245470 146180 245476 146192
rect 183704 146152 245476 146180
rect 183704 146140 183710 146152
rect 245470 146140 245476 146152
rect 245528 146180 245534 146192
rect 282178 146180 282184 146192
rect 245528 146152 282184 146180
rect 245528 146140 245534 146152
rect 282178 146140 282184 146152
rect 282236 146140 282242 146192
rect 189442 146072 189448 146124
rect 189500 146112 189506 146124
rect 251082 146112 251088 146124
rect 189500 146084 251088 146112
rect 189500 146072 189506 146084
rect 251082 146072 251088 146084
rect 251140 146072 251146 146124
rect 190638 146004 190644 146056
rect 190696 146044 190702 146056
rect 250990 146044 250996 146056
rect 190696 146016 250996 146044
rect 190696 146004 190702 146016
rect 250990 146004 250996 146016
rect 251048 146004 251054 146056
rect 195330 145936 195336 145988
rect 195388 145976 195394 145988
rect 253382 145976 253388 145988
rect 195388 145948 253388 145976
rect 195388 145936 195394 145948
rect 253382 145936 253388 145948
rect 253440 145936 253446 145988
rect 196710 145868 196716 145920
rect 196768 145908 196774 145920
rect 254854 145908 254860 145920
rect 196768 145880 254860 145908
rect 196768 145868 196774 145880
rect 254854 145868 254860 145880
rect 254912 145868 254918 145920
rect 197722 145800 197728 145852
rect 197780 145840 197786 145852
rect 254946 145840 254952 145852
rect 197780 145812 254952 145840
rect 197780 145800 197786 145812
rect 254946 145800 254952 145812
rect 255004 145800 255010 145852
rect 199378 145732 199384 145784
rect 199436 145772 199442 145784
rect 255958 145772 255964 145784
rect 199436 145744 255964 145772
rect 199436 145732 199442 145744
rect 255958 145732 255964 145744
rect 256016 145732 256022 145784
rect 251082 145664 251088 145716
rect 251140 145704 251146 145716
rect 356054 145704 356060 145716
rect 251140 145676 356060 145704
rect 251140 145664 251146 145676
rect 356054 145664 356060 145676
rect 356112 145664 356118 145716
rect 138014 145596 138020 145648
rect 138072 145636 138078 145648
rect 172882 145636 172888 145648
rect 138072 145608 172888 145636
rect 138072 145596 138078 145608
rect 172882 145596 172888 145608
rect 172940 145596 172946 145648
rect 250990 145596 250996 145648
rect 251048 145636 251054 145648
rect 369854 145636 369860 145648
rect 251048 145608 369860 145636
rect 251048 145596 251054 145608
rect 369854 145596 369860 145608
rect 369912 145596 369918 145648
rect 46198 145528 46204 145580
rect 46256 145568 46262 145580
rect 152458 145568 152464 145580
rect 46256 145540 152464 145568
rect 46256 145528 46262 145540
rect 152458 145528 152464 145540
rect 152516 145528 152522 145580
rect 155954 145528 155960 145580
rect 156012 145568 156018 145580
rect 174814 145568 174820 145580
rect 156012 145540 174820 145568
rect 156012 145528 156018 145540
rect 174814 145528 174820 145540
rect 174872 145528 174878 145580
rect 202414 145528 202420 145580
rect 202472 145568 202478 145580
rect 257338 145568 257344 145580
rect 202472 145540 257344 145568
rect 202472 145528 202478 145540
rect 257338 145528 257344 145540
rect 257396 145528 257402 145580
rect 294874 145528 294880 145580
rect 294932 145568 294938 145580
rect 514018 145568 514024 145580
rect 294932 145540 514024 145568
rect 294932 145528 294938 145540
rect 514018 145528 514024 145540
rect 514076 145528 514082 145580
rect 170030 145460 170036 145512
rect 170088 145500 170094 145512
rect 170490 145500 170496 145512
rect 170088 145472 170496 145500
rect 170088 145460 170094 145472
rect 170490 145460 170496 145472
rect 170548 145500 170554 145512
rect 222838 145500 222844 145512
rect 170548 145472 222844 145500
rect 170548 145460 170554 145472
rect 222838 145460 222844 145472
rect 222896 145460 222902 145512
rect 200482 145392 200488 145444
rect 200540 145432 200546 145444
rect 251818 145432 251824 145444
rect 200540 145404 251824 145432
rect 200540 145392 200546 145404
rect 251818 145392 251824 145404
rect 251876 145392 251882 145444
rect 199470 145324 199476 145376
rect 199528 145364 199534 145376
rect 226978 145364 226984 145376
rect 199528 145336 226984 145364
rect 199528 145324 199534 145336
rect 226978 145324 226984 145336
rect 227036 145324 227042 145376
rect 200942 145256 200948 145308
rect 201000 145296 201006 145308
rect 254762 145296 254768 145308
rect 201000 145268 254768 145296
rect 201000 145256 201006 145268
rect 254762 145256 254768 145268
rect 254820 145256 254826 145308
rect 200758 145188 200764 145240
rect 200816 145228 200822 145240
rect 254670 145228 254676 145240
rect 200816 145200 254676 145228
rect 200816 145188 200822 145200
rect 254670 145188 254676 145200
rect 254728 145188 254734 145240
rect 196158 144848 196164 144900
rect 196216 144888 196222 144900
rect 289262 144888 289268 144900
rect 196216 144860 289268 144888
rect 196216 144848 196222 144860
rect 289262 144848 289268 144860
rect 289320 144888 289326 144900
rect 289722 144888 289728 144900
rect 289320 144860 289728 144888
rect 289320 144848 289326 144860
rect 289722 144848 289728 144860
rect 289780 144848 289786 144900
rect 185118 144780 185124 144832
rect 185176 144820 185182 144832
rect 278130 144820 278136 144832
rect 185176 144792 278136 144820
rect 185176 144780 185182 144792
rect 278130 144780 278136 144792
rect 278188 144820 278194 144832
rect 284938 144820 284944 144832
rect 278188 144792 284944 144820
rect 278188 144780 278194 144792
rect 284938 144780 284944 144792
rect 284996 144780 285002 144832
rect 189350 144712 189356 144764
rect 189408 144752 189414 144764
rect 274634 144752 274640 144764
rect 189408 144724 274640 144752
rect 189408 144712 189414 144724
rect 274634 144712 274640 144724
rect 274692 144712 274698 144764
rect 175550 144644 175556 144696
rect 175608 144684 175614 144696
rect 176562 144684 176568 144696
rect 175608 144656 176568 144684
rect 175608 144644 175614 144656
rect 176562 144644 176568 144656
rect 176620 144644 176626 144696
rect 202874 144644 202880 144696
rect 202932 144684 202938 144696
rect 270310 144684 270316 144696
rect 202932 144656 270316 144684
rect 202932 144644 202938 144656
rect 270310 144644 270316 144656
rect 270368 144644 270374 144696
rect 198826 144576 198832 144628
rect 198884 144616 198890 144628
rect 260374 144616 260380 144628
rect 198884 144588 260380 144616
rect 198884 144576 198890 144588
rect 260374 144576 260380 144588
rect 260432 144576 260438 144628
rect 175458 144508 175464 144560
rect 175516 144548 175522 144560
rect 176470 144548 176476 144560
rect 175516 144520 176476 144548
rect 175516 144508 175522 144520
rect 176470 144508 176476 144520
rect 176528 144508 176534 144560
rect 238110 144548 238116 144560
rect 177960 144520 238116 144548
rect 177960 144424 177988 144520
rect 238110 144508 238116 144520
rect 238168 144508 238174 144560
rect 196250 144440 196256 144492
rect 196308 144480 196314 144492
rect 257522 144480 257528 144492
rect 196308 144452 257528 144480
rect 196308 144440 196314 144452
rect 257522 144440 257528 144452
rect 257580 144440 257586 144492
rect 176838 144372 176844 144424
rect 176896 144412 176902 144424
rect 177942 144412 177948 144424
rect 176896 144384 177948 144412
rect 176896 144372 176902 144384
rect 177942 144372 177948 144384
rect 178000 144372 178006 144424
rect 185210 144372 185216 144424
rect 185268 144412 185274 144424
rect 245102 144412 245108 144424
rect 185268 144384 245108 144412
rect 185268 144372 185274 144384
rect 245102 144372 245108 144384
rect 245160 144372 245166 144424
rect 205818 144304 205824 144356
rect 205876 144344 205882 144356
rect 206646 144344 206652 144356
rect 205876 144316 206652 144344
rect 205876 144304 205882 144316
rect 206646 144304 206652 144316
rect 206704 144344 206710 144356
rect 265434 144344 265440 144356
rect 206704 144316 265440 144344
rect 206704 144304 206710 144316
rect 265434 144304 265440 144316
rect 265492 144304 265498 144356
rect 274634 144304 274640 144356
rect 274692 144344 274698 144356
rect 341518 144344 341524 144356
rect 274692 144316 341524 144344
rect 274692 144304 274698 144316
rect 341518 144304 341524 144316
rect 341576 144304 341582 144356
rect 142154 144236 142160 144288
rect 142212 144276 142218 144288
rect 173434 144276 173440 144288
rect 142212 144248 173440 144276
rect 142212 144236 142218 144248
rect 173434 144236 173440 144248
rect 173492 144236 173498 144288
rect 177758 144236 177764 144288
rect 177816 144276 177822 144288
rect 231118 144276 231124 144288
rect 177816 144248 231124 144276
rect 177816 144236 177822 144248
rect 231118 144236 231124 144248
rect 231176 144236 231182 144288
rect 289722 144236 289728 144288
rect 289780 144276 289786 144288
rect 436738 144276 436744 144288
rect 289780 144248 436744 144276
rect 289780 144236 289786 144248
rect 436738 144236 436744 144248
rect 436796 144236 436802 144288
rect 75914 144168 75920 144220
rect 75972 144208 75978 144220
rect 166994 144208 167000 144220
rect 75972 144180 167000 144208
rect 75972 144168 75978 144180
rect 166994 144168 167000 144180
rect 167052 144168 167058 144220
rect 176470 144168 176476 144220
rect 176528 144208 176534 144220
rect 225782 144208 225788 144220
rect 176528 144180 225788 144208
rect 176528 144168 176534 144180
rect 225782 144168 225788 144180
rect 225840 144168 225846 144220
rect 270310 144168 270316 144220
rect 270368 144208 270374 144220
rect 532694 144208 532700 144220
rect 270368 144180 532700 144208
rect 270368 144168 270374 144180
rect 532694 144168 532700 144180
rect 532752 144168 532758 144220
rect 222930 144140 222936 144152
rect 190426 144112 222936 144140
rect 176562 143964 176568 144016
rect 176620 144004 176626 144016
rect 190426 144004 190454 144112
rect 222930 144100 222936 144112
rect 222988 144100 222994 144152
rect 176620 143976 190454 144004
rect 176620 143964 176626 143976
rect 177022 143556 177028 143608
rect 177080 143596 177086 143608
rect 177758 143596 177764 143608
rect 177080 143568 177764 143596
rect 177080 143556 177086 143568
rect 177758 143556 177764 143568
rect 177816 143556 177822 143608
rect 193306 143488 193312 143540
rect 193364 143528 193370 143540
rect 288526 143528 288532 143540
rect 193364 143500 288532 143528
rect 193364 143488 193370 143500
rect 288526 143488 288532 143500
rect 288584 143488 288590 143540
rect 186774 143420 186780 143472
rect 186832 143460 186838 143472
rect 277578 143460 277584 143472
rect 186832 143432 277584 143460
rect 186832 143420 186838 143432
rect 277578 143420 277584 143432
rect 277636 143460 277642 143472
rect 278682 143460 278688 143472
rect 277636 143432 278688 143460
rect 277636 143420 277642 143432
rect 278682 143420 278688 143432
rect 278740 143420 278746 143472
rect 197538 143352 197544 143404
rect 197596 143392 197602 143404
rect 282914 143392 282920 143404
rect 197596 143364 282920 143392
rect 197596 143352 197602 143364
rect 282914 143352 282920 143364
rect 282972 143352 282978 143404
rect 193950 143284 193956 143336
rect 194008 143324 194014 143336
rect 273254 143324 273260 143336
rect 194008 143296 273260 143324
rect 194008 143284 194014 143296
rect 273254 143284 273260 143296
rect 273312 143284 273318 143336
rect 203794 143216 203800 143268
rect 203852 143256 203858 143268
rect 271138 143256 271144 143268
rect 203852 143228 271144 143256
rect 203852 143216 203858 143228
rect 271138 143216 271144 143228
rect 271196 143216 271202 143268
rect 182358 143148 182364 143200
rect 182416 143188 182422 143200
rect 244182 143188 244188 143200
rect 182416 143160 244188 143188
rect 182416 143148 182422 143160
rect 244182 143148 244188 143160
rect 244240 143188 244246 143200
rect 244240 143160 248414 143188
rect 244240 143148 244246 143160
rect 177850 143080 177856 143132
rect 177908 143120 177914 143132
rect 220170 143120 220176 143132
rect 177908 143092 220176 143120
rect 177908 143080 177914 143092
rect 220170 143080 220176 143092
rect 220228 143080 220234 143132
rect 204438 143012 204444 143064
rect 204496 143052 204502 143064
rect 205266 143052 205272 143064
rect 204496 143024 205272 143052
rect 204496 143012 204502 143024
rect 205266 143012 205272 143024
rect 205324 143012 205330 143064
rect 118694 142944 118700 142996
rect 118752 142984 118758 142996
rect 172146 142984 172152 142996
rect 118752 142956 172152 142984
rect 118752 142944 118758 142956
rect 172146 142944 172152 142956
rect 172204 142944 172210 142996
rect 174630 142944 174636 142996
rect 174688 142984 174694 142996
rect 224218 142984 224224 142996
rect 174688 142956 224224 142984
rect 174688 142944 174694 142956
rect 224218 142944 224224 142956
rect 224276 142944 224282 142996
rect 60826 142876 60832 142928
rect 60884 142916 60890 142928
rect 167362 142916 167368 142928
rect 60884 142888 167368 142916
rect 60884 142876 60890 142888
rect 167362 142876 167368 142888
rect 167420 142876 167426 142928
rect 177298 142876 177304 142928
rect 177356 142916 177362 142928
rect 177850 142916 177856 142928
rect 177356 142888 177856 142916
rect 177356 142876 177362 142888
rect 177850 142876 177856 142888
rect 177908 142876 177914 142928
rect 229830 142916 229836 142928
rect 186286 142888 229836 142916
rect 35894 142808 35900 142860
rect 35952 142848 35958 142860
rect 164234 142848 164240 142860
rect 35952 142820 164240 142848
rect 35952 142808 35958 142820
rect 164234 142808 164240 142820
rect 164292 142808 164298 142860
rect 176746 142808 176752 142860
rect 176804 142848 176810 142860
rect 179322 142848 179328 142860
rect 176804 142820 179328 142848
rect 176804 142808 176810 142820
rect 179322 142808 179328 142820
rect 179380 142848 179386 142860
rect 186286 142848 186314 142888
rect 229830 142876 229836 142888
rect 229888 142876 229894 142928
rect 248386 142916 248414 143160
rect 278682 142944 278688 142996
rect 278740 142984 278746 142996
rect 309870 142984 309876 142996
rect 278740 142956 309876 142984
rect 278740 142944 278746 142956
rect 309870 142944 309876 142956
rect 309928 142944 309934 142996
rect 261478 142916 261484 142928
rect 248386 142888 261484 142916
rect 261478 142876 261484 142888
rect 261536 142876 261542 142928
rect 273254 142876 273260 142928
rect 273312 142916 273318 142928
rect 380894 142916 380900 142928
rect 273312 142888 380900 142916
rect 273312 142876 273318 142888
rect 380894 142876 380900 142888
rect 380952 142876 380958 142928
rect 179380 142820 186314 142848
rect 179380 142808 179386 142820
rect 205266 142808 205272 142860
rect 205324 142848 205330 142860
rect 263594 142848 263600 142860
rect 205324 142820 263600 142848
rect 205324 142808 205330 142820
rect 263594 142808 263600 142820
rect 263652 142808 263658 142860
rect 282914 142808 282920 142860
rect 282972 142848 282978 142860
rect 283742 142848 283748 142860
rect 282972 142820 283748 142848
rect 282972 142808 282978 142820
rect 283742 142808 283748 142820
rect 283800 142848 283806 142860
rect 449894 142848 449900 142860
rect 283800 142820 449900 142848
rect 283800 142808 283806 142820
rect 449894 142808 449900 142820
rect 449952 142808 449958 142860
rect 202690 142128 202696 142180
rect 202748 142168 202754 142180
rect 260834 142168 260840 142180
rect 202748 142140 260840 142168
rect 202748 142128 202754 142140
rect 260834 142128 260840 142140
rect 260892 142128 260898 142180
rect 193214 142060 193220 142112
rect 193272 142100 193278 142112
rect 285858 142100 285864 142112
rect 193272 142072 285864 142100
rect 193272 142060 193278 142072
rect 285858 142060 285864 142072
rect 285916 142060 285922 142112
rect 194686 141992 194692 142044
rect 194744 142032 194750 142044
rect 287514 142032 287520 142044
rect 194744 142004 287520 142032
rect 194744 141992 194750 142004
rect 287514 141992 287520 142004
rect 287572 141992 287578 142044
rect 198458 141924 198464 141976
rect 198516 141964 198522 141976
rect 287790 141964 287796 141976
rect 198516 141936 287796 141964
rect 198516 141924 198522 141936
rect 287790 141924 287796 141936
rect 287848 141924 287854 141976
rect 204898 141856 204904 141908
rect 204956 141896 204962 141908
rect 267734 141896 267740 141908
rect 204956 141868 267740 141896
rect 204956 141856 204962 141868
rect 267734 141856 267740 141868
rect 267792 141896 267798 141908
rect 269022 141896 269028 141908
rect 267792 141868 269028 141896
rect 267792 141856 267798 141868
rect 269022 141856 269028 141868
rect 269080 141856 269086 141908
rect 185026 141788 185032 141840
rect 185084 141828 185090 141840
rect 246942 141828 246948 141840
rect 185084 141800 246948 141828
rect 185084 141788 185090 141800
rect 246942 141788 246948 141800
rect 247000 141788 247006 141840
rect 164418 141720 164424 141772
rect 164476 141760 164482 141772
rect 223850 141760 223856 141772
rect 164476 141732 223856 141760
rect 164476 141720 164482 141732
rect 223850 141720 223856 141732
rect 223908 141720 223914 141772
rect 188982 141652 188988 141704
rect 189040 141692 189046 141704
rect 225874 141692 225880 141704
rect 189040 141664 225880 141692
rect 189040 141652 189046 141664
rect 225874 141652 225880 141664
rect 225932 141652 225938 141704
rect 189258 141584 189264 141636
rect 189316 141624 189322 141636
rect 190362 141624 190368 141636
rect 189316 141596 190368 141624
rect 189316 141584 189322 141596
rect 190362 141584 190368 141596
rect 190420 141624 190426 141636
rect 227070 141624 227076 141636
rect 190420 141596 227076 141624
rect 190420 141584 190426 141596
rect 227070 141584 227076 141596
rect 227128 141584 227134 141636
rect 246942 141584 246948 141636
rect 247000 141624 247006 141636
rect 302878 141624 302884 141636
rect 247000 141596 302884 141624
rect 247000 141584 247006 141596
rect 302878 141584 302884 141596
rect 302936 141584 302942 141636
rect 287514 141516 287520 141568
rect 287572 141556 287578 141568
rect 419534 141556 419540 141568
rect 287572 141528 419540 141556
rect 287572 141516 287578 141528
rect 419534 141516 419540 141528
rect 419592 141516 419598 141568
rect 92474 141448 92480 141500
rect 92532 141488 92538 141500
rect 168926 141488 168932 141500
rect 92532 141460 168932 141488
rect 92532 141448 92538 141460
rect 168926 141448 168932 141460
rect 168984 141448 168990 141500
rect 187786 141448 187792 141500
rect 187844 141488 187850 141500
rect 323578 141488 323584 141500
rect 187844 141460 323584 141488
rect 187844 141448 187850 141460
rect 323578 141448 323584 141460
rect 323636 141448 323642 141500
rect 48314 141380 48320 141432
rect 48372 141420 48378 141432
rect 165798 141420 165804 141432
rect 48372 141392 165804 141420
rect 48372 141380 48378 141392
rect 165798 141380 165804 141392
rect 165856 141380 165862 141432
rect 187878 141380 187884 141432
rect 187936 141420 187942 141432
rect 188982 141420 188988 141432
rect 187936 141392 188988 141420
rect 187936 141380 187942 141392
rect 188982 141380 188988 141392
rect 189040 141380 189046 141432
rect 269022 141380 269028 141432
rect 269080 141420 269086 141432
rect 550634 141420 550640 141432
rect 269080 141392 550640 141420
rect 269080 141380 269086 141392
rect 550634 141380 550640 141392
rect 550692 141380 550698 141432
rect 285858 140768 285864 140820
rect 285916 140808 285922 140820
rect 286318 140808 286324 140820
rect 285916 140780 286324 140808
rect 285916 140768 285922 140780
rect 286318 140768 286324 140780
rect 286376 140768 286382 140820
rect 182266 140700 182272 140752
rect 182324 140740 182330 140752
rect 183370 140740 183376 140752
rect 182324 140712 183376 140740
rect 182324 140700 182330 140712
rect 183370 140700 183376 140712
rect 183428 140700 183434 140752
rect 186590 140700 186596 140752
rect 186648 140740 186654 140752
rect 281534 140740 281540 140752
rect 186648 140712 281540 140740
rect 186648 140700 186654 140712
rect 281534 140700 281540 140712
rect 281592 140700 281598 140752
rect 197354 140632 197360 140684
rect 197412 140672 197418 140684
rect 261570 140672 261576 140684
rect 197412 140644 261576 140672
rect 197412 140632 197418 140644
rect 261570 140632 261576 140644
rect 261628 140632 261634 140684
rect 198642 140564 198648 140616
rect 198700 140604 198706 140616
rect 258810 140604 258816 140616
rect 198700 140576 258816 140604
rect 198700 140564 198706 140576
rect 258810 140564 258816 140576
rect 258868 140564 258874 140616
rect 183370 140496 183376 140548
rect 183428 140536 183434 140548
rect 241790 140536 241796 140548
rect 183428 140508 241796 140536
rect 183428 140496 183434 140508
rect 241790 140496 241796 140508
rect 241848 140496 241854 140548
rect 191650 140428 191656 140480
rect 191708 140468 191714 140480
rect 231210 140468 231216 140480
rect 191708 140440 231216 140468
rect 191708 140428 191714 140440
rect 231210 140428 231216 140440
rect 231268 140428 231274 140480
rect 189994 140360 190000 140412
rect 190052 140400 190058 140412
rect 225966 140400 225972 140412
rect 190052 140372 225972 140400
rect 190052 140360 190058 140372
rect 225966 140360 225972 140372
rect 226024 140360 226030 140412
rect 281534 140088 281540 140140
rect 281592 140128 281598 140140
rect 314010 140128 314016 140140
rect 281592 140100 314016 140128
rect 281592 140088 281598 140100
rect 314010 140088 314016 140100
rect 314068 140088 314074 140140
rect 20714 140020 20720 140072
rect 20772 140060 20778 140072
rect 162854 140060 162860 140072
rect 20772 140032 162860 140060
rect 20772 140020 20778 140032
rect 162854 140020 162860 140032
rect 162912 140020 162918 140072
rect 280798 140020 280804 140072
rect 280856 140060 280862 140072
rect 363598 140060 363604 140072
rect 280856 140032 363604 140060
rect 280856 140020 280862 140032
rect 363598 140020 363604 140032
rect 363656 140020 363662 140072
rect 186498 139340 186504 139392
rect 186556 139380 186562 139392
rect 282270 139380 282276 139392
rect 186556 139352 282276 139380
rect 186556 139340 186562 139352
rect 282270 139340 282276 139352
rect 282328 139340 282334 139392
rect 192110 139272 192116 139324
rect 192168 139312 192174 139324
rect 284386 139312 284392 139324
rect 192168 139284 284392 139312
rect 192168 139272 192174 139284
rect 284386 139272 284392 139284
rect 284444 139272 284450 139324
rect 184842 139204 184848 139256
rect 184900 139244 184906 139256
rect 244734 139244 244740 139256
rect 184900 139216 244740 139244
rect 184900 139204 184906 139216
rect 244734 139204 244740 139216
rect 244792 139244 244798 139256
rect 249058 139244 249064 139256
rect 244792 139216 249064 139244
rect 244792 139204 244798 139216
rect 249058 139204 249064 139216
rect 249116 139204 249122 139256
rect 167270 139136 167276 139188
rect 167328 139176 167334 139188
rect 167638 139176 167644 139188
rect 167328 139148 167644 139176
rect 167328 139136 167334 139148
rect 167638 139136 167644 139148
rect 167696 139176 167702 139188
rect 227714 139176 227720 139188
rect 167696 139148 227720 139176
rect 167696 139136 167702 139148
rect 227714 139136 227720 139148
rect 227772 139136 227778 139188
rect 166442 139068 166448 139120
rect 166500 139108 166506 139120
rect 225690 139108 225696 139120
rect 166500 139080 225696 139108
rect 166500 139068 166506 139080
rect 225690 139068 225696 139080
rect 225748 139068 225754 139120
rect 168558 139000 168564 139052
rect 168616 139040 168622 139052
rect 169110 139040 169116 139052
rect 168616 139012 169116 139040
rect 168616 139000 168622 139012
rect 169110 139000 169116 139012
rect 169168 139040 169174 139052
rect 228450 139040 228456 139052
rect 169168 139012 228456 139040
rect 169168 139000 169174 139012
rect 228450 139000 228456 139012
rect 228508 139000 228514 139052
rect 122834 138728 122840 138780
rect 122892 138768 122898 138780
rect 171686 138768 171692 138780
rect 122892 138740 171692 138768
rect 122892 138728 122898 138740
rect 171686 138728 171692 138740
rect 171744 138728 171750 138780
rect 282270 138728 282276 138780
rect 282328 138768 282334 138780
rect 320174 138768 320180 138780
rect 282328 138740 320180 138768
rect 282328 138728 282334 138740
rect 320174 138728 320180 138740
rect 320232 138728 320238 138780
rect 40034 138660 40040 138712
rect 40092 138700 40098 138712
rect 164418 138700 164424 138712
rect 40092 138672 164424 138700
rect 40092 138660 40098 138672
rect 164418 138660 164424 138672
rect 164476 138660 164482 138712
rect 284386 138660 284392 138712
rect 284444 138700 284450 138712
rect 383654 138700 383660 138712
rect 284444 138672 383660 138700
rect 284444 138660 284450 138672
rect 383654 138660 383660 138672
rect 383712 138660 383718 138712
rect 3050 137912 3056 137964
rect 3108 137952 3114 137964
rect 159358 137952 159364 137964
rect 3108 137924 159364 137952
rect 3108 137912 3114 137924
rect 159358 137912 159364 137924
rect 159416 137912 159422 137964
rect 187694 137912 187700 137964
rect 187752 137952 187758 137964
rect 282914 137952 282920 137964
rect 187752 137924 282920 137952
rect 187752 137912 187758 137924
rect 282914 137912 282920 137924
rect 282972 137912 282978 137964
rect 205174 137844 205180 137896
rect 205232 137884 205238 137896
rect 272702 137884 272708 137896
rect 205232 137856 272708 137884
rect 205232 137844 205238 137856
rect 272702 137844 272708 137856
rect 272760 137844 272766 137896
rect 167730 137776 167736 137828
rect 167788 137816 167794 137828
rect 168006 137816 168012 137828
rect 167788 137788 168012 137816
rect 167788 137776 167794 137788
rect 168006 137776 168012 137788
rect 168064 137816 168070 137828
rect 223758 137816 223764 137828
rect 168064 137788 223764 137816
rect 168064 137776 168070 137788
rect 223758 137776 223764 137788
rect 223816 137776 223822 137828
rect 282914 137368 282920 137420
rect 282972 137408 282978 137420
rect 283558 137408 283564 137420
rect 282972 137380 283564 137408
rect 282972 137368 282978 137380
rect 283558 137368 283564 137380
rect 283616 137408 283622 137420
rect 338114 137408 338120 137420
rect 283616 137380 338120 137408
rect 283616 137368 283622 137380
rect 338114 137368 338120 137380
rect 338172 137368 338178 137420
rect 288526 137300 288532 137352
rect 288584 137340 288590 137352
rect 405734 137340 405740 137352
rect 288584 137312 405740 137340
rect 288584 137300 288590 137312
rect 405734 137300 405740 137312
rect 405792 137300 405798 137352
rect 146294 137232 146300 137284
rect 146352 137272 146358 137284
rect 173158 137272 173164 137284
rect 146352 137244 173164 137272
rect 146352 137232 146358 137244
rect 173158 137232 173164 137244
rect 173216 137232 173222 137284
rect 180610 137232 180616 137284
rect 180668 137272 180674 137284
rect 219434 137272 219440 137284
rect 180668 137244 219440 137272
rect 180668 137232 180674 137244
rect 219434 137232 219440 137244
rect 219492 137232 219498 137284
rect 272702 137232 272708 137284
rect 272760 137272 272766 137284
rect 554774 137272 554780 137284
rect 272760 137244 554780 137272
rect 272760 137232 272766 137244
rect 554774 137232 554780 137244
rect 554832 137232 554838 137284
rect 205726 136552 205732 136604
rect 205784 136592 205790 136604
rect 272242 136592 272248 136604
rect 205784 136564 272248 136592
rect 205784 136552 205790 136564
rect 272242 136552 272248 136564
rect 272300 136552 272306 136604
rect 196066 136484 196072 136536
rect 196124 136524 196130 136536
rect 255866 136524 255872 136536
rect 196124 136496 255872 136524
rect 196124 136484 196130 136496
rect 255866 136484 255872 136496
rect 255924 136484 255930 136536
rect 189166 136416 189172 136468
rect 189224 136456 189230 136468
rect 247310 136456 247316 136468
rect 189224 136428 247316 136456
rect 189224 136416 189230 136428
rect 247310 136416 247316 136428
rect 247368 136416 247374 136468
rect 79318 135940 79324 135992
rect 79376 135980 79382 135992
rect 168558 135980 168564 135992
rect 79376 135952 168564 135980
rect 79376 135940 79382 135952
rect 168558 135940 168564 135952
rect 168616 135940 168622 135992
rect 247310 135940 247316 135992
rect 247368 135980 247374 135992
rect 248230 135980 248236 135992
rect 247368 135952 248236 135980
rect 247368 135940 247374 135952
rect 248230 135940 248236 135952
rect 248288 135980 248294 135992
rect 351914 135980 351920 135992
rect 248288 135952 351920 135980
rect 248288 135940 248294 135952
rect 351914 135940 351920 135952
rect 351972 135940 351978 135992
rect 55214 135872 55220 135924
rect 55272 135912 55278 135924
rect 166442 135912 166448 135924
rect 55272 135884 166448 135912
rect 55272 135872 55278 135884
rect 166442 135872 166448 135884
rect 166500 135872 166506 135924
rect 255866 135872 255872 135924
rect 255924 135912 255930 135924
rect 256602 135912 256608 135924
rect 255924 135884 256608 135912
rect 255924 135872 255930 135884
rect 256602 135872 256608 135884
rect 256660 135912 256666 135924
rect 440234 135912 440240 135924
rect 256660 135884 440240 135912
rect 256660 135872 256666 135884
rect 440234 135872 440240 135884
rect 440292 135872 440298 135924
rect 272242 135260 272248 135312
rect 272300 135300 272306 135312
rect 568574 135300 568580 135312
rect 272300 135272 568580 135300
rect 272300 135260 272306 135272
rect 568574 135260 568580 135272
rect 568632 135260 568638 135312
rect 206370 135192 206376 135244
rect 206428 135232 206434 135244
rect 270494 135232 270500 135244
rect 206428 135204 270500 135232
rect 206428 135192 206434 135204
rect 270494 135192 270500 135204
rect 270552 135232 270558 135244
rect 271782 135232 271788 135244
rect 270552 135204 271788 135232
rect 270552 135192 270558 135204
rect 271782 135192 271788 135204
rect 271840 135192 271846 135244
rect 190546 135124 190552 135176
rect 190604 135164 190610 135176
rect 249702 135164 249708 135176
rect 190604 135136 249708 135164
rect 190604 135124 190610 135136
rect 249702 135124 249708 135136
rect 249760 135124 249766 135176
rect 249702 134648 249708 134700
rect 249760 134688 249766 134700
rect 351178 134688 351184 134700
rect 249760 134660 351184 134688
rect 249760 134648 249766 134660
rect 351178 134648 351184 134660
rect 351236 134648 351242 134700
rect 287790 134580 287796 134632
rect 287848 134620 287854 134632
rect 455414 134620 455420 134632
rect 287848 134592 455420 134620
rect 287848 134580 287854 134592
rect 455414 134580 455420 134592
rect 455472 134580 455478 134632
rect 18598 134512 18604 134564
rect 18656 134552 18662 134564
rect 161658 134552 161664 134564
rect 18656 134524 161664 134552
rect 18656 134512 18662 134524
rect 161658 134512 161664 134524
rect 161716 134512 161722 134564
rect 181990 134512 181996 134564
rect 182048 134552 182054 134564
rect 241514 134552 241520 134564
rect 182048 134524 241520 134552
rect 182048 134512 182054 134524
rect 241514 134512 241520 134524
rect 241572 134512 241578 134564
rect 271782 134512 271788 134564
rect 271840 134552 271846 134564
rect 549898 134552 549904 134564
rect 271840 134524 549904 134552
rect 271840 134512 271846 134524
rect 549898 134512 549904 134524
rect 549956 134512 549962 134564
rect 192018 133832 192024 133884
rect 192076 133872 192082 133884
rect 252462 133872 252468 133884
rect 192076 133844 252468 133872
rect 192076 133832 192082 133844
rect 252462 133832 252468 133844
rect 252520 133832 252526 133884
rect 102134 133220 102140 133272
rect 102192 133260 102198 133272
rect 169846 133260 169852 133272
rect 102192 133232 169852 133260
rect 102192 133220 102198 133232
rect 169846 133220 169852 133232
rect 169904 133220 169910 133272
rect 252462 133220 252468 133272
rect 252520 133260 252526 133272
rect 390554 133260 390560 133272
rect 252520 133232 390560 133260
rect 252520 133220 252526 133232
rect 390554 133220 390560 133232
rect 390612 133220 390618 133272
rect 8294 133152 8300 133204
rect 8352 133192 8358 133204
rect 163682 133192 163688 133204
rect 8352 133164 163688 133192
rect 8352 133152 8358 133164
rect 163682 133152 163688 133164
rect 163740 133152 163746 133204
rect 208118 133152 208124 133204
rect 208176 133192 208182 133204
rect 575474 133192 575480 133204
rect 208176 133164 575480 133192
rect 208176 133152 208182 133164
rect 575474 133152 575480 133164
rect 575532 133152 575538 133204
rect 191926 132404 191932 132456
rect 191984 132444 191990 132456
rect 287146 132444 287152 132456
rect 191984 132416 287152 132444
rect 191984 132404 191990 132416
rect 287146 132404 287152 132416
rect 287204 132444 287210 132456
rect 288342 132444 288348 132456
rect 287204 132416 288348 132444
rect 287204 132404 287210 132416
rect 288342 132404 288348 132416
rect 288400 132404 288406 132456
rect 186406 132336 186412 132388
rect 186464 132376 186470 132388
rect 248322 132376 248328 132388
rect 186464 132348 248328 132376
rect 186464 132336 186470 132348
rect 248322 132336 248328 132348
rect 248380 132336 248386 132388
rect 248322 131792 248328 131844
rect 248380 131832 248386 131844
rect 287698 131832 287704 131844
rect 248380 131804 287704 131832
rect 248380 131792 248386 131804
rect 287698 131792 287704 131804
rect 287756 131792 287762 131844
rect 111794 131724 111800 131776
rect 111852 131764 111858 131776
rect 172330 131764 172336 131776
rect 111852 131736 172336 131764
rect 111852 131724 111858 131736
rect 172330 131724 172336 131736
rect 172388 131724 172394 131776
rect 288342 131724 288348 131776
rect 288400 131764 288406 131776
rect 387794 131764 387800 131776
rect 288400 131736 387800 131764
rect 288400 131724 288406 131736
rect 387794 131724 387800 131736
rect 387852 131724 387858 131776
rect 84194 130364 84200 130416
rect 84252 130404 84258 130416
rect 169202 130404 169208 130416
rect 84252 130376 169208 130404
rect 84252 130364 84258 130376
rect 169202 130364 169208 130376
rect 169260 130364 169266 130416
rect 286318 130364 286324 130416
rect 286376 130404 286382 130416
rect 408494 130404 408500 130416
rect 286376 130376 408500 130404
rect 286376 130364 286382 130376
rect 408494 130364 408500 130376
rect 408552 130364 408558 130416
rect 199838 129684 199844 129736
rect 199896 129724 199902 129736
rect 270402 129724 270408 129736
rect 199896 129696 270408 129724
rect 199896 129684 199902 129696
rect 270402 129684 270408 129696
rect 270460 129684 270466 129736
rect 195606 129616 195612 129668
rect 195664 129656 195670 129668
rect 253842 129656 253848 129668
rect 195664 129628 253848 129656
rect 195664 129616 195670 129628
rect 253842 129616 253848 129628
rect 253900 129616 253906 129668
rect 97994 129072 98000 129124
rect 98052 129112 98058 129124
rect 170490 129112 170496 129124
rect 98052 129084 170496 129112
rect 98052 129072 98058 129084
rect 170490 129072 170496 129084
rect 170548 129072 170554 129124
rect 253842 129072 253848 129124
rect 253900 129112 253906 129124
rect 422938 129112 422944 129124
rect 253900 129084 422944 129112
rect 253900 129072 253906 129084
rect 422938 129072 422944 129084
rect 422996 129072 423002 129124
rect 25498 129004 25504 129056
rect 25556 129044 25562 129056
rect 163038 129044 163044 129056
rect 25556 129016 163044 129044
rect 25556 129004 25562 129016
rect 163038 129004 163044 129016
rect 163096 129004 163102 129056
rect 182082 129004 182088 129056
rect 182140 129044 182146 129056
rect 237374 129044 237380 129056
rect 182140 129016 237380 129044
rect 182140 129004 182146 129016
rect 237374 129004 237380 129016
rect 237432 129004 237438 129056
rect 270402 129004 270408 129056
rect 270460 129044 270466 129056
rect 480254 129044 480260 129056
rect 270460 129016 480260 129044
rect 270460 129004 270466 129016
rect 480254 129004 480260 129016
rect 480312 129004 480318 129056
rect 189074 128256 189080 128308
rect 189132 128296 189138 128308
rect 284294 128296 284300 128308
rect 189132 128268 284300 128296
rect 189132 128256 189138 128268
rect 284294 128256 284300 128268
rect 284352 128256 284358 128308
rect 195974 128188 195980 128240
rect 196032 128228 196038 128240
rect 291194 128228 291200 128240
rect 196032 128200 291200 128228
rect 196032 128188 196038 128200
rect 291194 128188 291200 128200
rect 291252 128228 291258 128240
rect 291654 128228 291660 128240
rect 291252 128200 291660 128228
rect 291252 128188 291258 128200
rect 291654 128188 291660 128200
rect 291712 128188 291718 128240
rect 117314 127644 117320 127696
rect 117372 127684 117378 127696
rect 171410 127684 171416 127696
rect 117372 127656 171416 127684
rect 117372 127644 117378 127656
rect 171410 127644 171416 127656
rect 171468 127644 171474 127696
rect 284294 127644 284300 127696
rect 284352 127684 284358 127696
rect 358814 127684 358820 127696
rect 284352 127656 358820 127684
rect 284352 127644 284358 127656
rect 358814 127644 358820 127656
rect 358872 127644 358878 127696
rect 66254 127576 66260 127628
rect 66312 127616 66318 127628
rect 167638 127616 167644 127628
rect 66312 127588 167644 127616
rect 66312 127576 66318 127588
rect 167638 127576 167644 127588
rect 167696 127576 167702 127628
rect 291654 127576 291660 127628
rect 291712 127616 291718 127628
rect 444374 127616 444380 127628
rect 291712 127588 444380 127616
rect 291712 127576 291718 127588
rect 444374 127576 444380 127588
rect 444432 127576 444438 127628
rect 200114 126896 200120 126948
rect 200172 126936 200178 126948
rect 273898 126936 273904 126948
rect 200172 126908 273904 126936
rect 200172 126896 200178 126908
rect 273898 126896 273904 126908
rect 273956 126936 273962 126948
rect 274082 126936 274088 126948
rect 273956 126908 274088 126936
rect 273956 126896 273962 126908
rect 274082 126896 274088 126908
rect 274140 126896 274146 126948
rect 261570 126284 261576 126336
rect 261628 126324 261634 126336
rect 458174 126324 458180 126336
rect 261628 126296 458180 126324
rect 261628 126284 261634 126296
rect 458174 126284 458180 126296
rect 458232 126284 458238 126336
rect 69014 126216 69020 126268
rect 69072 126256 69078 126268
rect 167822 126256 167828 126268
rect 69072 126228 167828 126256
rect 69072 126216 69078 126228
rect 167822 126216 167828 126228
rect 167880 126216 167886 126268
rect 274082 126216 274088 126268
rect 274140 126256 274146 126268
rect 489914 126256 489920 126268
rect 274140 126228 489920 126256
rect 274140 126216 274146 126228
rect 489914 126216 489920 126228
rect 489972 126216 489978 126268
rect 190454 125536 190460 125588
rect 190512 125576 190518 125588
rect 285766 125576 285772 125588
rect 190512 125548 285772 125576
rect 190512 125536 190518 125548
rect 285766 125536 285772 125548
rect 285824 125576 285830 125588
rect 286226 125576 286232 125588
rect 285824 125548 286232 125576
rect 285824 125536 285830 125548
rect 286226 125536 286232 125548
rect 286284 125536 286290 125588
rect 115934 124924 115940 124976
rect 115992 124964 115998 124976
rect 171318 124964 171324 124976
rect 115992 124936 171324 124964
rect 115992 124924 115998 124936
rect 171318 124924 171324 124936
rect 171376 124924 171382 124976
rect 15838 124856 15844 124908
rect 15896 124896 15902 124908
rect 162946 124896 162952 124908
rect 15896 124868 162952 124896
rect 15896 124856 15902 124868
rect 162946 124856 162952 124868
rect 163004 124856 163010 124908
rect 286226 124856 286232 124908
rect 286284 124896 286290 124908
rect 376754 124896 376760 124908
rect 286284 124868 376760 124896
rect 286284 124856 286290 124868
rect 376754 124856 376760 124868
rect 376812 124856 376818 124908
rect 201586 124108 201592 124160
rect 201644 124148 201650 124160
rect 294506 124148 294512 124160
rect 201644 124120 294512 124148
rect 201644 124108 201650 124120
rect 294506 124108 294512 124120
rect 294564 124108 294570 124160
rect 111058 123496 111064 123548
rect 111116 123536 111122 123548
rect 170766 123536 170772 123548
rect 111116 123508 170772 123536
rect 111116 123496 111122 123508
rect 170766 123496 170772 123508
rect 170824 123496 170830 123548
rect 191834 123496 191840 123548
rect 191892 123536 191898 123548
rect 394694 123536 394700 123548
rect 191892 123508 394700 123536
rect 191892 123496 191898 123508
rect 394694 123496 394700 123508
rect 394752 123496 394758 123548
rect 14458 123428 14464 123480
rect 14516 123468 14522 123480
rect 161566 123468 161572 123480
rect 14516 123440 161572 123468
rect 14516 123428 14522 123440
rect 161566 123428 161572 123440
rect 161624 123428 161630 123480
rect 294506 123428 294512 123480
rect 294564 123468 294570 123480
rect 503714 123468 503720 123480
rect 294564 123440 503720 123468
rect 294564 123428 294570 123440
rect 503714 123428 503720 123440
rect 503772 123428 503778 123480
rect 86954 122068 86960 122120
rect 87012 122108 87018 122120
rect 169018 122108 169024 122120
rect 87012 122080 169024 122108
rect 87012 122068 87018 122080
rect 169018 122068 169024 122080
rect 169076 122068 169082 122120
rect 203886 122068 203892 122120
rect 203944 122108 203950 122120
rect 520918 122108 520924 122120
rect 203944 122080 520924 122108
rect 203944 122068 203950 122080
rect 520918 122068 520924 122080
rect 520976 122068 520982 122120
rect 23474 120708 23480 120760
rect 23532 120748 23538 120760
rect 164602 120748 164608 120760
rect 23532 120720 164608 120748
rect 23532 120708 23538 120720
rect 164602 120708 164608 120720
rect 164660 120708 164666 120760
rect 205266 120708 205272 120760
rect 205324 120748 205330 120760
rect 539686 120748 539692 120760
rect 205324 120720 539692 120748
rect 205324 120708 205330 120720
rect 539686 120708 539692 120720
rect 539744 120708 539750 120760
rect 19334 119348 19340 119400
rect 19392 119388 19398 119400
rect 161014 119388 161020 119400
rect 19392 119360 161020 119388
rect 19392 119348 19398 119360
rect 161014 119348 161020 119360
rect 161072 119348 161078 119400
rect 22738 117920 22744 117972
rect 22796 117960 22802 117972
rect 163406 117960 163412 117972
rect 22796 117932 163412 117960
rect 22796 117920 22802 117932
rect 163406 117920 163412 117932
rect 163464 117920 163470 117972
rect 163498 117920 163504 117972
rect 163556 117960 163562 117972
rect 174814 117960 174820 117972
rect 163556 117932 174820 117960
rect 163556 117920 163562 117932
rect 174814 117920 174820 117932
rect 174872 117920 174878 117972
rect 187510 116628 187516 116680
rect 187568 116668 187574 116680
rect 307846 116668 307852 116680
rect 187568 116640 307852 116668
rect 187568 116628 187574 116640
rect 307846 116628 307852 116640
rect 307904 116628 307910 116680
rect 22094 116560 22100 116612
rect 22152 116600 22158 116612
rect 163590 116600 163596 116612
rect 22152 116572 163596 116600
rect 22152 116560 22158 116572
rect 163590 116560 163596 116572
rect 163648 116560 163654 116612
rect 198550 116560 198556 116612
rect 198608 116600 198614 116612
rect 462314 116600 462320 116612
rect 198608 116572 462320 116600
rect 198608 116560 198614 116572
rect 462314 116560 462320 116572
rect 462372 116560 462378 116612
rect 39298 115200 39304 115252
rect 39356 115240 39362 115252
rect 164694 115240 164700 115252
rect 39356 115212 164700 115240
rect 39356 115200 39362 115212
rect 164694 115200 164700 115212
rect 164752 115200 164758 115252
rect 166350 112412 166356 112464
rect 166408 112452 166414 112464
rect 174078 112452 174084 112464
rect 166408 112424 174084 112452
rect 166408 112412 166414 112424
rect 174078 112412 174084 112424
rect 174136 112412 174142 112464
rect 194410 112412 194416 112464
rect 194468 112452 194474 112464
rect 404354 112452 404360 112464
rect 194468 112424 404360 112452
rect 194468 112412 194474 112424
rect 404354 112412 404360 112424
rect 404412 112412 404418 112464
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 142798 111772 142804 111784
rect 3384 111744 142804 111772
rect 3384 111732 3390 111744
rect 142798 111732 142804 111744
rect 142856 111732 142862 111784
rect 183370 111052 183376 111104
rect 183428 111092 183434 111104
rect 262214 111092 262220 111104
rect 183428 111064 262220 111092
rect 183428 111052 183434 111064
rect 262214 111052 262220 111064
rect 262272 111052 262278 111104
rect 9674 109692 9680 109744
rect 9732 109732 9738 109744
rect 163314 109732 163320 109744
rect 9732 109704 163320 109732
rect 9732 109692 9738 109704
rect 163314 109692 163320 109704
rect 163372 109692 163378 109744
rect 49694 108264 49700 108316
rect 49752 108304 49758 108316
rect 166074 108304 166080 108316
rect 49752 108276 166080 108304
rect 49752 108264 49758 108276
rect 166074 108264 166080 108276
rect 166132 108264 166138 108316
rect 178034 108264 178040 108316
rect 178092 108304 178098 108316
rect 200758 108304 200764 108316
rect 178092 108276 200764 108304
rect 178092 108264 178098 108276
rect 200758 108264 200764 108276
rect 200816 108264 200822 108316
rect 201310 108264 201316 108316
rect 201368 108304 201374 108316
rect 492674 108304 492680 108316
rect 201368 108276 492680 108304
rect 201368 108264 201374 108276
rect 492674 108264 492680 108276
rect 492732 108264 492738 108316
rect 63494 106904 63500 106956
rect 63552 106944 63558 106956
rect 167546 106944 167552 106956
rect 63552 106916 167552 106944
rect 63552 106904 63558 106916
rect 167546 106904 167552 106916
rect 167604 106904 167610 106956
rect 167638 106904 167644 106956
rect 167696 106944 167702 106956
rect 174722 106944 174728 106956
rect 167696 106916 174728 106944
rect 167696 106904 167702 106916
rect 174722 106904 174728 106916
rect 174780 106904 174786 106956
rect 70394 105544 70400 105596
rect 70452 105584 70458 105596
rect 167454 105584 167460 105596
rect 70452 105556 167460 105584
rect 70452 105544 70458 105556
rect 167454 105544 167460 105556
rect 167512 105544 167518 105596
rect 201402 105544 201408 105596
rect 201460 105584 201466 105596
rect 499574 105584 499580 105596
rect 201460 105556 499580 105584
rect 201460 105544 201466 105556
rect 499574 105544 499580 105556
rect 499632 105544 499638 105596
rect 88334 104116 88340 104168
rect 88392 104156 88398 104168
rect 168742 104156 168748 104168
rect 88392 104128 168748 104156
rect 88392 104116 88398 104128
rect 168742 104116 168748 104128
rect 168800 104116 168806 104168
rect 177666 104116 177672 104168
rect 177724 104156 177730 104168
rect 189718 104156 189724 104168
rect 177724 104128 189724 104156
rect 177724 104116 177730 104128
rect 189718 104116 189724 104128
rect 189776 104116 189782 104168
rect 190362 104116 190368 104168
rect 190420 104156 190426 104168
rect 347774 104156 347780 104168
rect 190420 104128 347780 104156
rect 190420 104116 190426 104128
rect 347774 104116 347780 104128
rect 347832 104116 347838 104168
rect 102226 102756 102232 102808
rect 102284 102796 102290 102808
rect 171042 102796 171048 102808
rect 102284 102768 171048 102796
rect 102284 102756 102290 102768
rect 171042 102756 171048 102768
rect 171100 102756 171106 102808
rect 202690 102756 202696 102808
rect 202748 102796 202754 102808
rect 510614 102796 510620 102808
rect 202748 102768 510620 102796
rect 202748 102756 202754 102768
rect 510614 102756 510620 102768
rect 510672 102756 510678 102808
rect 120074 101396 120080 101448
rect 120132 101436 120138 101448
rect 171870 101436 171876 101448
rect 120132 101408 171876 101436
rect 120132 101396 120138 101408
rect 171870 101396 171876 101408
rect 171928 101396 171934 101448
rect 337378 100648 337384 100700
rect 337436 100688 337442 100700
rect 580166 100688 580172 100700
rect 337436 100660 580172 100688
rect 337436 100648 337442 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 31754 99968 31760 100020
rect 31812 100008 31818 100020
rect 164970 100008 164976 100020
rect 31812 99980 164976 100008
rect 31812 99968 31818 99980
rect 164970 99968 164976 99980
rect 165028 99968 165034 100020
rect 176470 99288 176476 99340
rect 176528 99328 176534 99340
rect 180794 99328 180800 99340
rect 176528 99300 180800 99328
rect 176528 99288 176534 99300
rect 180794 99288 180800 99300
rect 180852 99288 180858 99340
rect 27614 98608 27620 98660
rect 27672 98648 27678 98660
rect 158346 98648 158352 98660
rect 27672 98620 158352 98648
rect 27672 98608 27678 98620
rect 158346 98608 158352 98620
rect 158404 98608 158410 98660
rect 53834 97316 53840 97368
rect 53892 97356 53898 97368
rect 165614 97356 165620 97368
rect 53892 97328 165620 97356
rect 53892 97316 53898 97328
rect 165614 97316 165620 97328
rect 165672 97316 165678 97368
rect 161934 97248 161940 97300
rect 161992 97288 161998 97300
rect 580258 97288 580264 97300
rect 161992 97260 580264 97288
rect 161992 97248 161998 97260
rect 580258 97248 580264 97260
rect 580316 97248 580322 97300
rect 11698 95888 11704 95940
rect 11756 95928 11762 95940
rect 163222 95928 163228 95940
rect 11756 95900 163228 95928
rect 11756 95888 11762 95900
rect 163222 95888 163228 95900
rect 163280 95888 163286 95940
rect 183462 94528 183468 94580
rect 183520 94568 183526 94580
rect 269114 94568 269120 94580
rect 183520 94540 269120 94568
rect 183520 94528 183526 94540
rect 269114 94528 269120 94540
rect 269172 94528 269178 94580
rect 42794 94460 42800 94512
rect 42852 94500 42858 94512
rect 148318 94500 148324 94512
rect 42852 94472 148324 94500
rect 42852 94460 42858 94472
rect 148318 94460 148324 94472
rect 148376 94460 148382 94512
rect 203978 94460 203984 94512
rect 204036 94500 204042 94512
rect 535454 94500 535460 94512
rect 204036 94472 535460 94500
rect 204036 94460 204042 94472
rect 535454 94460 535460 94472
rect 535512 94460 535518 94512
rect 180702 93168 180708 93220
rect 180760 93208 180766 93220
rect 234706 93208 234712 93220
rect 180760 93180 234712 93208
rect 180760 93168 180766 93180
rect 234706 93168 234712 93180
rect 234764 93168 234770 93220
rect 204346 93100 204352 93152
rect 204404 93140 204410 93152
rect 542354 93140 542360 93152
rect 204404 93112 542360 93140
rect 204404 93100 204410 93112
rect 542354 93100 542360 93112
rect 542412 93100 542418 93152
rect 205450 91740 205456 91792
rect 205508 91780 205514 91792
rect 546494 91780 546500 91792
rect 205508 91752 546500 91780
rect 205508 91740 205514 91752
rect 546494 91740 546500 91752
rect 546552 91740 546558 91792
rect 206646 88952 206652 89004
rect 206704 88992 206710 89004
rect 552658 88992 552664 89004
rect 206704 88964 552664 88992
rect 206704 88952 206710 88964
rect 552658 88952 552664 88964
rect 552716 88952 552722 89004
rect 205542 87592 205548 87644
rect 205600 87632 205606 87644
rect 553394 87632 553400 87644
rect 205600 87604 553400 87632
rect 205600 87592 205606 87604
rect 553394 87592 553400 87604
rect 553452 87592 553458 87644
rect 206554 86232 206560 86284
rect 206612 86272 206618 86284
rect 560294 86272 560300 86284
rect 206612 86244 560300 86272
rect 206612 86232 206618 86244
rect 560294 86232 560300 86244
rect 560352 86232 560358 86284
rect 208210 83444 208216 83496
rect 208268 83484 208274 83496
rect 574094 83484 574100 83496
rect 208268 83456 574100 83484
rect 208268 83444 208274 83456
rect 574094 83444 574100 83456
rect 574152 83444 574158 83496
rect 206830 82084 206836 82136
rect 206888 82124 206894 82136
rect 567194 82124 567200 82136
rect 206888 82096 567200 82124
rect 206888 82084 206894 82096
rect 567194 82084 567200 82096
rect 567252 82084 567258 82136
rect 208302 80656 208308 80708
rect 208360 80696 208366 80708
rect 578234 80696 578240 80708
rect 208360 80668 578240 80696
rect 208360 80656 208366 80668
rect 578234 80656 578240 80668
rect 578292 80656 578298 80708
rect 194502 79296 194508 79348
rect 194560 79336 194566 79348
rect 400214 79336 400220 79348
rect 194560 79308 400220 79336
rect 194560 79296 194566 79308
rect 400214 79296 400220 79308
rect 400272 79296 400278 79348
rect 162026 73788 162032 73840
rect 162084 73828 162090 73840
rect 580258 73828 580264 73840
rect 162084 73800 580264 73828
rect 162084 73788 162090 73800
rect 580258 73788 580264 73800
rect 580316 73788 580322 73840
rect 188890 72428 188896 72480
rect 188948 72468 188954 72480
rect 331858 72468 331864 72480
rect 188948 72440 331864 72468
rect 188948 72428 188954 72440
rect 331858 72428 331864 72440
rect 331916 72428 331922 72480
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 120718 71720 120724 71732
rect 3568 71692 120724 71720
rect 3568 71680 3574 71692
rect 120718 71680 120724 71692
rect 120776 71680 120782 71732
rect 177758 66852 177764 66904
rect 177816 66892 177822 66904
rect 187694 66892 187700 66904
rect 177816 66864 187700 66892
rect 177816 66852 177822 66864
rect 187694 66852 187700 66864
rect 187752 66852 187758 66904
rect 95970 59984 95976 60036
rect 96028 60024 96034 60036
rect 170582 60024 170588 60036
rect 96028 59996 170588 60024
rect 96028 59984 96034 59996
rect 170582 59984 170588 59996
rect 170640 59984 170646 60036
rect 177850 59984 177856 60036
rect 177908 60024 177914 60036
rect 191098 60024 191104 60036
rect 177908 59996 191104 60024
rect 177908 59984 177914 59996
rect 191098 59984 191104 59996
rect 191156 59984 191162 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 95878 59344 95884 59356
rect 3108 59316 95884 59344
rect 3108 59304 3114 59316
rect 95878 59304 95884 59316
rect 95936 59304 95942 59356
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 155218 45540 155224 45552
rect 3568 45512 155224 45540
rect 3568 45500 3574 45512
rect 155218 45500 155224 45512
rect 155276 45500 155282 45552
rect 75178 37884 75184 37936
rect 75236 37924 75242 37936
rect 167730 37924 167736 37936
rect 75236 37896 167736 37924
rect 75236 37884 75242 37896
rect 167730 37884 167736 37896
rect 167788 37884 167794 37936
rect 204070 36524 204076 36576
rect 204128 36564 204134 36576
rect 525794 36564 525800 36576
rect 204128 36536 525800 36564
rect 204128 36524 204134 36536
rect 525794 36524 525800 36536
rect 525852 36524 525858 36576
rect 179230 33736 179236 33788
rect 179288 33776 179294 33788
rect 205634 33776 205640 33788
rect 179288 33748 205640 33776
rect 179288 33736 179294 33748
rect 205634 33736 205640 33748
rect 205692 33736 205698 33788
rect 206922 33736 206928 33788
rect 206980 33776 206986 33788
rect 564526 33776 564532 33788
rect 206980 33748 564532 33776
rect 206980 33736 206986 33748
rect 564526 33736 564532 33748
rect 564584 33736 564590 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 43438 33096 43444 33108
rect 2924 33068 43444 33096
rect 2924 33056 2930 33068
rect 43438 33056 43444 33068
rect 43496 33056 43502 33108
rect 280062 33056 280068 33108
rect 280120 33096 280126 33108
rect 580166 33096 580172 33108
rect 280120 33068 580172 33096
rect 280120 33056 280126 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 203610 28228 203616 28280
rect 203668 28268 203674 28280
rect 524414 28268 524420 28280
rect 203668 28240 524420 28268
rect 203668 28228 203674 28240
rect 524414 28228 524420 28240
rect 524472 28228 524478 28280
rect 175918 23468 175924 23520
rect 175976 23508 175982 23520
rect 176654 23508 176660 23520
rect 175976 23480 176660 23508
rect 175976 23468 175982 23480
rect 176654 23468 176660 23480
rect 176712 23468 176718 23520
rect 187602 22720 187608 22772
rect 187660 22760 187666 22772
rect 315390 22760 315396 22772
rect 187660 22732 315396 22760
rect 187660 22720 187666 22732
rect 315390 22720 315396 22732
rect 315448 22720 315454 22772
rect 334618 20612 334624 20664
rect 334676 20652 334682 20664
rect 580074 20652 580080 20664
rect 334676 20624 580080 20652
rect 334676 20612 334682 20624
rect 580074 20612 580080 20624
rect 580132 20612 580138 20664
rect 202782 17212 202788 17264
rect 202840 17252 202846 17264
rect 505094 17252 505100 17264
rect 202840 17224 505100 17252
rect 202840 17212 202846 17224
rect 505094 17212 505100 17224
rect 505152 17212 505158 17264
rect 39114 15852 39120 15904
rect 39172 15892 39178 15904
rect 164786 15892 164792 15904
rect 39172 15864 164792 15892
rect 39172 15852 39178 15864
rect 164786 15852 164792 15864
rect 164844 15852 164850 15904
rect 177942 15852 177948 15904
rect 178000 15892 178006 15904
rect 195146 15892 195152 15904
rect 178000 15864 195152 15892
rect 178000 15852 178006 15864
rect 195146 15852 195152 15864
rect 195204 15852 195210 15904
rect 195790 15852 195796 15904
rect 195848 15892 195854 15904
rect 429194 15892 429200 15904
rect 195848 15864 429200 15892
rect 195848 15852 195854 15864
rect 429194 15852 429200 15864
rect 429252 15852 429258 15904
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 124858 14464 124864 14476
rect 11204 14436 124864 14464
rect 11204 14424 11210 14436
rect 124858 14424 124864 14436
rect 124916 14424 124922 14476
rect 25314 13064 25320 13116
rect 25372 13104 25378 13116
rect 164878 13104 164884 13116
rect 25372 13076 164884 13104
rect 25372 13064 25378 13076
rect 164878 13064 164884 13076
rect 164936 13064 164942 13116
rect 197446 13064 197452 13116
rect 197504 13104 197510 13116
rect 465166 13104 465172 13116
rect 197504 13076 465172 13104
rect 197504 13064 197510 13076
rect 465166 13064 465172 13076
rect 465224 13064 465230 13116
rect 160094 11772 160100 11824
rect 160152 11812 160158 11824
rect 161290 11812 161296 11824
rect 160152 11784 161296 11812
rect 160152 11772 160158 11784
rect 161290 11772 161296 11784
rect 161348 11772 161354 11824
rect 46106 11704 46112 11756
rect 46164 11744 46170 11756
rect 166258 11744 166264 11756
rect 46164 11716 166264 11744
rect 46164 11704 46170 11716
rect 166258 11704 166264 11716
rect 166316 11704 166322 11756
rect 198734 11704 198740 11756
rect 198792 11744 198798 11756
rect 478874 11744 478880 11756
rect 198792 11716 478880 11744
rect 198792 11704 198798 11716
rect 478874 11704 478880 11716
rect 478932 11704 478938 11756
rect 35986 10276 35992 10328
rect 36044 10316 36050 10328
rect 151078 10316 151084 10328
rect 36044 10288 151084 10316
rect 36044 10276 36050 10288
rect 151078 10276 151084 10288
rect 151136 10276 151142 10328
rect 200022 10276 200028 10328
rect 200080 10316 200086 10328
rect 472250 10316 472256 10328
rect 200080 10288 472256 10316
rect 200080 10276 200086 10288
rect 472250 10276 472256 10288
rect 472308 10276 472314 10328
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 193122 8984 193128 9036
rect 193180 9024 193186 9036
rect 383562 9024 383568 9036
rect 193180 8996 383568 9024
rect 193180 8984 193186 8996
rect 383562 8984 383568 8996
rect 383620 8984 383626 9036
rect 110506 8916 110512 8968
rect 110564 8956 110570 8968
rect 170398 8956 170404 8968
rect 110564 8928 170404 8956
rect 110564 8916 110570 8928
rect 170398 8916 170404 8928
rect 170456 8916 170462 8968
rect 195882 8916 195888 8968
rect 195940 8956 195946 8968
rect 418982 8956 418988 8968
rect 195940 8928 418988 8956
rect 195940 8916 195946 8928
rect 418982 8916 418988 8928
rect 419040 8916 419046 8968
rect 176562 8236 176568 8288
rect 176620 8276 176626 8288
rect 177850 8276 177856 8288
rect 176620 8248 177856 8276
rect 176620 8236 176626 8248
rect 177850 8236 177856 8248
rect 177908 8236 177914 8288
rect 78582 7556 78588 7608
rect 78640 7596 78646 7608
rect 168466 7596 168472 7608
rect 78640 7568 168472 7596
rect 78640 7556 78646 7568
rect 168466 7556 168472 7568
rect 168524 7556 168530 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 146938 6848 146944 6860
rect 3476 6820 146944 6848
rect 3476 6808 3482 6820
rect 146938 6808 146944 6820
rect 146996 6808 147002 6860
rect 191742 6264 191748 6316
rect 191800 6304 191806 6316
rect 369394 6304 369400 6316
rect 191800 6276 369400 6304
rect 191800 6264 191806 6276
rect 369394 6264 369400 6276
rect 369452 6264 369458 6316
rect 191650 6196 191656 6248
rect 191708 6236 191714 6248
rect 372890 6236 372896 6248
rect 191708 6208 372896 6236
rect 191708 6196 191714 6208
rect 372890 6196 372896 6208
rect 372948 6196 372954 6248
rect 197262 6128 197268 6180
rect 197320 6168 197326 6180
rect 436646 6168 436652 6180
rect 197320 6140 436652 6168
rect 197320 6128 197326 6140
rect 436646 6128 436652 6140
rect 436704 6128 436710 6180
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 156598 4808 156604 4820
rect 19484 4780 156604 4808
rect 19484 4768 19490 4780
rect 156598 4768 156604 4780
rect 156656 4768 156662 4820
rect 188982 4768 188988 4820
rect 189040 4808 189046 4820
rect 330386 4808 330392 4820
rect 189040 4780 330392 4808
rect 189040 4768 189046 4780
rect 330386 4768 330392 4780
rect 330444 4768 330450 4820
rect 315298 4156 315304 4208
rect 315356 4196 315362 4208
rect 315356 4168 316264 4196
rect 315356 4156 315362 4168
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 149514 4088 149520 4140
rect 149572 4128 149578 4140
rect 153838 4128 153844 4140
rect 149572 4100 153844 4128
rect 149572 4088 149578 4100
rect 153838 4088 153844 4100
rect 153896 4088 153902 4140
rect 209682 4088 209688 4140
rect 209740 4128 209746 4140
rect 210970 4128 210976 4140
rect 209740 4100 210976 4128
rect 209740 4088 209746 4100
rect 210970 4088 210976 4100
rect 211028 4088 211034 4140
rect 243722 4088 243728 4140
rect 243780 4128 243786 4140
rect 254670 4128 254676 4140
rect 243780 4100 254676 4128
rect 243780 4088 243786 4100
rect 254670 4088 254676 4100
rect 254728 4088 254734 4140
rect 275278 4088 275284 4140
rect 275336 4128 275342 4140
rect 278314 4128 278320 4140
rect 275336 4100 278320 4128
rect 275336 4088 275342 4100
rect 278314 4088 278320 4100
rect 278372 4088 278378 4140
rect 315390 4088 315396 4140
rect 315448 4128 315454 4140
rect 316034 4128 316040 4140
rect 315448 4100 316040 4128
rect 315448 4088 315454 4100
rect 316034 4088 316040 4100
rect 316092 4088 316098 4140
rect 171410 4020 171416 4072
rect 171468 4060 171474 4072
rect 171778 4060 171784 4072
rect 171468 4032 171784 4060
rect 171468 4020 171474 4032
rect 171778 4020 171784 4032
rect 171836 4020 171842 4072
rect 193858 4020 193864 4072
rect 193916 4060 193922 4072
rect 200298 4060 200304 4072
rect 193916 4032 200304 4060
rect 193916 4020 193922 4032
rect 200298 4020 200304 4032
rect 200356 4020 200362 4072
rect 240870 4020 240876 4072
rect 240928 4060 240934 4072
rect 251174 4060 251180 4072
rect 240928 4032 251180 4060
rect 240928 4020 240934 4032
rect 251174 4020 251180 4032
rect 251232 4020 251238 4072
rect 314010 4020 314016 4072
rect 314068 4060 314074 4072
rect 316236 4060 316264 4168
rect 316678 4088 316684 4140
rect 316736 4128 316742 4140
rect 323670 4128 323676 4140
rect 316736 4100 323676 4128
rect 316736 4088 316742 4100
rect 323670 4088 323676 4100
rect 323728 4088 323734 4140
rect 571978 4088 571984 4140
rect 572036 4128 572042 4140
rect 577406 4128 577412 4140
rect 572036 4100 577412 4128
rect 572036 4088 572042 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 326798 4060 326804 4072
rect 314068 4032 316172 4060
rect 316236 4032 326804 4060
rect 314068 4020 314074 4032
rect 239398 3952 239404 4004
rect 239456 3992 239462 4004
rect 249978 3992 249984 4004
rect 239456 3964 249984 3992
rect 239456 3952 239462 3964
rect 249978 3952 249984 3964
rect 250036 3952 250042 4004
rect 250438 3952 250444 4004
rect 250496 3992 250502 4004
rect 260650 3992 260656 4004
rect 250496 3964 260656 3992
rect 250496 3952 250502 3964
rect 260650 3952 260656 3964
rect 260708 3952 260714 4004
rect 313182 3952 313188 4004
rect 313240 3992 313246 4004
rect 316144 3992 316172 4032
rect 326798 4020 326804 4032
rect 326856 4020 326862 4072
rect 507118 4020 507124 4072
rect 507176 4060 507182 4072
rect 510062 4060 510068 4072
rect 507176 4032 510068 4060
rect 507176 4020 507182 4032
rect 510062 4020 510068 4032
rect 510120 4020 510126 4072
rect 317322 3992 317328 4004
rect 313240 3964 316080 3992
rect 316144 3964 317328 3992
rect 313240 3952 313246 3964
rect 235258 3884 235264 3936
rect 235316 3924 235322 3936
rect 246390 3924 246396 3936
rect 235316 3896 246396 3924
rect 235316 3884 235322 3896
rect 246390 3884 246396 3896
rect 246448 3884 246454 3936
rect 246574 3884 246580 3936
rect 246632 3924 246638 3936
rect 257062 3924 257068 3936
rect 246632 3896 257068 3924
rect 246632 3884 246638 3896
rect 257062 3884 257068 3896
rect 257120 3884 257126 3936
rect 264238 3884 264244 3936
rect 264296 3924 264302 3936
rect 267734 3924 267740 3936
rect 264296 3896 267740 3924
rect 264296 3884 264302 3896
rect 267734 3884 267740 3896
rect 267792 3884 267798 3936
rect 302878 3884 302884 3936
rect 302936 3924 302942 3936
rect 306742 3924 306748 3936
rect 302936 3896 306748 3924
rect 302936 3884 302942 3896
rect 306742 3884 306748 3896
rect 306800 3884 306806 3936
rect 316052 3924 316080 3964
rect 317322 3952 317328 3964
rect 317380 3952 317386 4004
rect 325602 3992 325608 4004
rect 320744 3964 325608 3992
rect 320744 3924 320772 3964
rect 325602 3952 325608 3964
rect 325660 3952 325666 4004
rect 431218 3952 431224 4004
rect 431276 3992 431282 4004
rect 434438 3992 434444 4004
rect 431276 3964 434444 3992
rect 431276 3952 431282 3964
rect 434438 3952 434444 3964
rect 434496 3952 434502 4004
rect 316052 3896 320772 3924
rect 323670 3884 323676 3936
rect 323728 3924 323734 3936
rect 331582 3924 331588 3936
rect 323728 3896 331588 3924
rect 323728 3884 323734 3896
rect 331582 3884 331588 3896
rect 331640 3884 331646 3936
rect 363598 3884 363604 3936
rect 363656 3924 363662 3936
rect 367002 3924 367008 3936
rect 363656 3896 367008 3924
rect 363656 3884 363662 3896
rect 367002 3884 367008 3896
rect 367060 3884 367066 3936
rect 44266 3816 44272 3868
rect 44324 3856 44330 3868
rect 46198 3856 46204 3868
rect 44324 3828 46204 3856
rect 44324 3816 44330 3828
rect 46198 3816 46204 3828
rect 46256 3816 46262 3868
rect 244918 3816 244924 3868
rect 244976 3856 244982 3868
rect 258258 3856 258264 3868
rect 244976 3828 258264 3856
rect 244976 3816 244982 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 261478 3816 261484 3868
rect 261536 3856 261542 3868
rect 271230 3856 271236 3868
rect 261536 3828 271236 3856
rect 261536 3816 261542 3828
rect 271230 3816 271236 3828
rect 271288 3816 271294 3868
rect 305638 3816 305644 3868
rect 305696 3856 305702 3868
rect 314010 3856 314016 3868
rect 305696 3828 314016 3856
rect 305696 3816 305702 3828
rect 314010 3816 314016 3828
rect 314068 3816 314074 3868
rect 323578 3816 323584 3868
rect 323636 3856 323642 3868
rect 342162 3856 342168 3868
rect 323636 3828 342168 3856
rect 323636 3816 323642 3828
rect 342162 3816 342168 3828
rect 342220 3816 342226 3868
rect 179322 3748 179328 3800
rect 179380 3788 179386 3800
rect 184934 3788 184940 3800
rect 179380 3760 184940 3788
rect 179380 3748 179386 3760
rect 184934 3748 184940 3760
rect 184992 3748 184998 3800
rect 213178 3748 213184 3800
rect 213236 3788 213242 3800
rect 225138 3788 225144 3800
rect 213236 3760 225144 3788
rect 213236 3748 213242 3760
rect 225138 3748 225144 3760
rect 225196 3748 225202 3800
rect 236638 3748 236644 3800
rect 236696 3788 236702 3800
rect 240502 3788 240508 3800
rect 236696 3760 240508 3788
rect 236696 3748 236702 3760
rect 240502 3748 240508 3760
rect 240560 3748 240566 3800
rect 242158 3748 242164 3800
rect 242216 3788 242222 3800
rect 265342 3788 265348 3800
rect 242216 3760 265348 3788
rect 242216 3748 242222 3760
rect 265342 3748 265348 3760
rect 265400 3748 265406 3800
rect 268378 3748 268384 3800
rect 268436 3788 268442 3800
rect 283098 3788 283104 3800
rect 268436 3760 283104 3788
rect 268436 3748 268442 3760
rect 283098 3748 283104 3760
rect 283156 3748 283162 3800
rect 307110 3748 307116 3800
rect 307168 3788 307174 3800
rect 329190 3788 329196 3800
rect 307168 3760 329196 3788
rect 307168 3748 307174 3760
rect 329190 3748 329196 3760
rect 329248 3748 329254 3800
rect 118786 3680 118792 3732
rect 118844 3720 118850 3732
rect 127618 3720 127624 3732
rect 118844 3692 127624 3720
rect 118844 3680 118850 3692
rect 127618 3680 127624 3692
rect 127676 3680 127682 3732
rect 189810 3680 189816 3732
rect 189868 3720 189874 3732
rect 194410 3720 194416 3732
rect 189868 3692 194416 3720
rect 189868 3680 189874 3692
rect 194410 3680 194416 3692
rect 194468 3680 194474 3732
rect 211798 3680 211804 3732
rect 211856 3720 211862 3732
rect 221550 3720 221556 3732
rect 211856 3692 221556 3720
rect 211856 3680 211862 3692
rect 221550 3680 221556 3692
rect 221608 3680 221614 3732
rect 228358 3680 228364 3732
rect 228416 3720 228422 3732
rect 235810 3720 235816 3732
rect 228416 3692 235816 3720
rect 228416 3680 228422 3692
rect 235810 3680 235816 3692
rect 235868 3680 235874 3732
rect 243630 3680 243636 3732
rect 243688 3720 243694 3732
rect 268838 3720 268844 3732
rect 243688 3692 268844 3720
rect 243688 3680 243694 3692
rect 268838 3680 268844 3692
rect 268896 3680 268902 3732
rect 284938 3680 284944 3732
rect 284996 3720 285002 3732
rect 303154 3720 303160 3732
rect 284996 3692 303160 3720
rect 284996 3680 285002 3692
rect 303154 3680 303160 3692
rect 303212 3680 303218 3732
rect 308398 3680 308404 3732
rect 308456 3720 308462 3732
rect 332594 3720 332600 3732
rect 308456 3692 332600 3720
rect 308456 3680 308462 3692
rect 332594 3680 332600 3692
rect 332652 3680 332658 3732
rect 374086 3680 374092 3732
rect 374144 3720 374150 3732
rect 375282 3720 375288 3732
rect 374144 3692 375288 3720
rect 374144 3680 374150 3692
rect 375282 3680 375288 3692
rect 375340 3680 375346 3732
rect 376018 3680 376024 3732
rect 376076 3720 376082 3732
rect 398834 3720 398840 3732
rect 376076 3692 398840 3720
rect 376076 3680 376082 3692
rect 398834 3680 398840 3692
rect 398892 3680 398898 3732
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 11698 3652 11704 3664
rect 6512 3624 11704 3652
rect 6512 3612 6518 3624
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 14458 3652 14464 3664
rect 11808 3624 14464 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 11808 3584 11836 3624
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 25498 3652 25504 3664
rect 14792 3624 25504 3652
rect 14792 3612 14798 3624
rect 25498 3612 25504 3624
rect 25556 3612 25562 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 130378 3652 130384 3664
rect 96304 3624 130384 3652
rect 96304 3612 96310 3624
rect 130378 3612 130384 3624
rect 130436 3612 130442 3664
rect 180150 3612 180156 3664
rect 180208 3652 180214 3664
rect 190822 3652 190828 3664
rect 180208 3624 190828 3652
rect 180208 3612 180214 3624
rect 190822 3612 190828 3624
rect 190880 3612 190886 3664
rect 196802 3652 196808 3664
rect 190932 3624 196808 3652
rect 1728 3556 11836 3584
rect 1728 3544 1734 3556
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 15838 3584 15844 3596
rect 13596 3556 15844 3584
rect 13596 3544 13602 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 60734 3544 60740 3596
rect 60792 3584 60798 3596
rect 61654 3584 61660 3596
rect 60792 3556 61660 3584
rect 60792 3544 60798 3556
rect 61654 3544 61660 3556
rect 61712 3544 61718 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 71038 3584 71044 3596
rect 69164 3556 71044 3584
rect 69164 3544 69170 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 86862 3544 86868 3596
rect 86920 3584 86926 3596
rect 88978 3584 88984 3596
rect 86920 3556 88984 3584
rect 86920 3544 86926 3556
rect 88978 3544 88984 3556
rect 89036 3544 89042 3596
rect 95142 3544 95148 3596
rect 95200 3584 95206 3596
rect 95970 3584 95976 3596
rect 95200 3556 95976 3584
rect 95200 3544 95206 3556
rect 95970 3544 95976 3556
rect 96028 3544 96034 3596
rect 110414 3544 110420 3596
rect 110472 3584 110478 3596
rect 111610 3584 111616 3596
rect 110472 3556 111616 3584
rect 110472 3544 110478 3556
rect 111610 3544 111616 3556
rect 111668 3544 111674 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 115198 3584 115204 3596
rect 114060 3556 115204 3584
rect 114060 3544 114066 3556
rect 115198 3544 115204 3556
rect 115256 3544 115262 3596
rect 118694 3544 118700 3596
rect 118752 3584 118758 3596
rect 119890 3584 119896 3596
rect 118752 3556 119896 3584
rect 118752 3544 118758 3556
rect 119890 3544 119896 3556
rect 119948 3544 119954 3596
rect 124674 3544 124680 3596
rect 124732 3584 124738 3596
rect 160738 3584 160744 3596
rect 124732 3556 160744 3584
rect 124732 3544 124738 3556
rect 160738 3544 160744 3556
rect 160796 3544 160802 3596
rect 162762 3544 162768 3596
rect 162820 3584 162826 3596
rect 166074 3584 166080 3596
rect 162820 3556 166080 3584
rect 162820 3544 162826 3556
rect 166074 3544 166080 3556
rect 166132 3544 166138 3596
rect 180058 3544 180064 3596
rect 180116 3544 180122 3596
rect 182910 3544 182916 3596
rect 182968 3584 182974 3596
rect 190932 3584 190960 3624
rect 196802 3612 196808 3624
rect 196860 3612 196866 3664
rect 220078 3612 220084 3664
rect 220136 3652 220142 3664
rect 220136 3624 229094 3652
rect 220136 3612 220142 3624
rect 193214 3584 193220 3596
rect 182968 3556 190960 3584
rect 191024 3556 193220 3584
rect 182968 3544 182974 3556
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 18598 3516 18604 3528
rect 4120 3488 18604 3516
rect 4120 3476 4126 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 31294 3476 31300 3528
rect 31352 3516 31358 3528
rect 32398 3516 32404 3528
rect 31352 3488 32404 3516
rect 31352 3476 31358 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 39298 3516 39304 3528
rect 38436 3488 39304 3516
rect 38436 3476 38442 3488
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 53742 3476 53748 3528
rect 53800 3516 53806 3528
rect 162118 3516 162124 3528
rect 53800 3488 162124 3516
rect 53800 3476 53806 3488
rect 162118 3476 162124 3488
rect 162176 3476 162182 3528
rect 162486 3476 162492 3528
rect 162544 3516 162550 3528
rect 163498 3516 163504 3528
rect 162544 3488 163504 3516
rect 162544 3476 162550 3488
rect 163498 3476 163504 3488
rect 163556 3476 163562 3528
rect 164878 3476 164884 3528
rect 164936 3516 164942 3528
rect 167638 3516 167644 3528
rect 164936 3488 167644 3516
rect 164936 3476 164942 3488
rect 167638 3476 167644 3488
rect 167696 3476 167702 3528
rect 170766 3476 170772 3528
rect 170824 3516 170830 3528
rect 174630 3516 174636 3528
rect 170824 3488 174636 3516
rect 170824 3476 170830 3488
rect 174630 3476 174636 3488
rect 174688 3476 174694 3528
rect 180076 3516 180104 3544
rect 191024 3516 191052 3556
rect 193214 3544 193220 3556
rect 193272 3544 193278 3596
rect 225598 3544 225604 3596
rect 225656 3584 225662 3596
rect 228726 3584 228732 3596
rect 225656 3556 228732 3584
rect 225656 3544 225662 3556
rect 228726 3544 228732 3556
rect 228784 3544 228790 3596
rect 229066 3584 229094 3624
rect 232498 3612 232504 3664
rect 232556 3652 232562 3664
rect 242894 3652 242900 3664
rect 232556 3624 242900 3652
rect 232556 3612 232562 3624
rect 242894 3612 242900 3624
rect 242952 3612 242958 3664
rect 243538 3612 243544 3664
rect 243596 3652 243602 3664
rect 276014 3652 276020 3664
rect 243596 3624 276020 3652
rect 243596 3612 243602 3624
rect 276014 3612 276020 3624
rect 276072 3612 276078 3664
rect 287698 3612 287704 3664
rect 287756 3652 287762 3664
rect 324406 3652 324412 3664
rect 287756 3624 324412 3652
rect 287756 3612 287762 3624
rect 324406 3612 324412 3624
rect 324464 3612 324470 3664
rect 327718 3612 327724 3664
rect 327776 3652 327782 3664
rect 339862 3652 339868 3664
rect 327776 3624 339868 3652
rect 327776 3612 327782 3624
rect 339862 3612 339868 3624
rect 339920 3612 339926 3664
rect 341518 3612 341524 3664
rect 341576 3652 341582 3664
rect 349154 3652 349160 3664
rect 341576 3624 349160 3652
rect 341576 3612 341582 3624
rect 349154 3612 349160 3624
rect 349212 3612 349218 3664
rect 355318 3612 355324 3664
rect 355376 3652 355382 3664
rect 402514 3652 402520 3664
rect 355376 3624 402520 3652
rect 355376 3612 355382 3624
rect 402514 3612 402520 3624
rect 402572 3612 402578 3664
rect 423766 3612 423772 3664
rect 423824 3652 423830 3664
rect 424962 3652 424968 3664
rect 423824 3624 424968 3652
rect 423824 3612 423830 3624
rect 424962 3612 424968 3624
rect 425020 3612 425026 3664
rect 448606 3612 448612 3664
rect 448664 3652 448670 3664
rect 449802 3652 449808 3664
rect 448664 3624 449808 3652
rect 448664 3612 448670 3624
rect 449802 3612 449808 3624
rect 449860 3612 449866 3664
rect 552658 3612 552664 3664
rect 552716 3652 552722 3664
rect 557350 3652 557356 3664
rect 552716 3624 557356 3652
rect 552716 3612 552722 3624
rect 557350 3612 557356 3624
rect 557408 3612 557414 3664
rect 253474 3584 253480 3596
rect 229066 3556 253480 3584
rect 253474 3544 253480 3556
rect 253532 3544 253538 3596
rect 253566 3544 253572 3596
rect 253624 3584 253630 3596
rect 260006 3584 260012 3596
rect 253624 3556 260012 3584
rect 253624 3544 253630 3556
rect 260006 3544 260012 3556
rect 260064 3544 260070 3596
rect 260098 3544 260104 3596
rect 260156 3584 260162 3596
rect 261754 3584 261760 3596
rect 260156 3556 261760 3584
rect 260156 3544 260162 3556
rect 261754 3544 261760 3556
rect 261812 3544 261818 3596
rect 265618 3544 265624 3596
rect 265676 3584 265682 3596
rect 266538 3584 266544 3596
rect 265676 3556 266544 3584
rect 265676 3544 265682 3556
rect 266538 3544 266544 3556
rect 266596 3544 266602 3596
rect 266998 3544 267004 3596
rect 267056 3584 267062 3596
rect 292574 3584 292580 3596
rect 267056 3556 292580 3584
rect 267056 3544 267062 3556
rect 292574 3544 292580 3556
rect 292632 3544 292638 3596
rect 295978 3544 295984 3596
rect 296036 3584 296042 3596
rect 299658 3584 299664 3596
rect 296036 3556 299664 3584
rect 296036 3544 296042 3556
rect 299658 3544 299664 3556
rect 299716 3544 299722 3596
rect 307846 3544 307852 3596
rect 307904 3584 307910 3596
rect 309042 3584 309048 3596
rect 307904 3556 309048 3584
rect 307904 3544 307910 3556
rect 309042 3544 309048 3556
rect 309100 3544 309106 3596
rect 311434 3584 311440 3596
rect 311084 3556 311440 3584
rect 180076 3488 191052 3516
rect 191098 3476 191104 3528
rect 191156 3516 191162 3528
rect 192018 3516 192024 3528
rect 191156 3488 192024 3516
rect 191156 3476 191162 3488
rect 192018 3476 192024 3488
rect 192076 3476 192082 3528
rect 197998 3476 198004 3528
rect 198056 3516 198062 3528
rect 199102 3516 199108 3528
rect 198056 3488 199108 3516
rect 198056 3476 198062 3488
rect 199102 3476 199108 3488
rect 199160 3476 199166 3528
rect 217318 3476 217324 3528
rect 217376 3516 217382 3528
rect 239306 3516 239312 3528
rect 217376 3488 239312 3516
rect 217376 3476 217382 3488
rect 239306 3476 239312 3488
rect 239364 3476 239370 3528
rect 240778 3476 240784 3528
rect 240836 3516 240842 3528
rect 247586 3516 247592 3528
rect 240836 3488 247592 3516
rect 240836 3476 240842 3488
rect 247586 3476 247592 3488
rect 247644 3476 247650 3528
rect 249058 3476 249064 3528
rect 249116 3516 249122 3528
rect 288986 3516 288992 3528
rect 249116 3488 288992 3516
rect 249116 3476 249122 3488
rect 288986 3476 288992 3488
rect 289044 3476 289050 3528
rect 289078 3476 289084 3528
rect 289136 3516 289142 3528
rect 290182 3516 290188 3528
rect 289136 3488 290188 3516
rect 289136 3476 289142 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 305730 3476 305736 3528
rect 305788 3516 305794 3528
rect 311084 3516 311112 3556
rect 311434 3544 311440 3556
rect 311492 3544 311498 3596
rect 320818 3544 320824 3596
rect 320876 3584 320882 3596
rect 346946 3584 346952 3596
rect 320876 3556 346952 3584
rect 320876 3544 320882 3556
rect 346946 3544 346952 3556
rect 347004 3544 347010 3596
rect 349246 3544 349252 3596
rect 349304 3584 349310 3596
rect 350442 3584 350448 3596
rect 349304 3556 350448 3584
rect 349304 3544 349310 3556
rect 350442 3544 350448 3556
rect 350500 3544 350506 3596
rect 351270 3544 351276 3596
rect 351328 3584 351334 3596
rect 374086 3584 374092 3596
rect 351328 3556 374092 3584
rect 351328 3544 351334 3556
rect 374086 3544 374092 3556
rect 374144 3544 374150 3596
rect 378042 3544 378048 3596
rect 378100 3584 378106 3596
rect 463970 3584 463976 3596
rect 378100 3556 463976 3584
rect 378100 3544 378106 3556
rect 463970 3544 463976 3556
rect 464028 3544 464034 3596
rect 471238 3544 471244 3596
rect 471296 3584 471302 3596
rect 474550 3584 474556 3596
rect 471296 3556 474556 3584
rect 471296 3544 471302 3556
rect 474550 3544 474556 3556
rect 474608 3544 474614 3596
rect 547874 3544 547880 3596
rect 547932 3584 547938 3596
rect 548702 3584 548708 3596
rect 547932 3556 548708 3584
rect 547932 3544 547938 3556
rect 548702 3544 548708 3556
rect 548760 3544 548766 3596
rect 549898 3544 549904 3596
rect 549956 3584 549962 3596
rect 572714 3584 572720 3596
rect 549956 3556 572720 3584
rect 549956 3544 549962 3556
rect 572714 3544 572720 3556
rect 572772 3544 572778 3596
rect 305788 3488 311112 3516
rect 305788 3476 305794 3488
rect 311158 3476 311164 3528
rect 311216 3516 311222 3528
rect 312630 3516 312636 3528
rect 311216 3488 312636 3516
rect 311216 3476 311222 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 313918 3476 313924 3528
rect 313976 3516 313982 3528
rect 313976 3488 415256 3516
rect 313976 3476 313982 3488
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 126238 3448 126244 3460
rect 2924 3420 126244 3448
rect 2924 3408 2930 3420
rect 126238 3408 126244 3420
rect 126296 3408 126302 3460
rect 126974 3408 126980 3460
rect 127032 3448 127038 3460
rect 128170 3448 128176 3460
rect 127032 3420 128176 3448
rect 127032 3408 127038 3420
rect 128170 3408 128176 3420
rect 128228 3408 128234 3460
rect 135254 3408 135260 3460
rect 135312 3448 135318 3460
rect 136450 3448 136456 3460
rect 135312 3420 136456 3448
rect 135312 3408 135318 3420
rect 136450 3408 136456 3420
rect 136508 3408 136514 3460
rect 169570 3408 169576 3460
rect 169628 3448 169634 3460
rect 174538 3448 174544 3460
rect 169628 3420 174544 3448
rect 169628 3408 169634 3420
rect 174538 3408 174544 3420
rect 174596 3408 174602 3460
rect 181530 3408 181536 3460
rect 181588 3448 181594 3460
rect 183738 3448 183744 3460
rect 181588 3420 183744 3448
rect 181588 3408 181594 3420
rect 183738 3408 183744 3420
rect 183796 3408 183802 3460
rect 207382 3448 207388 3460
rect 190426 3420 207388 3448
rect 109310 3340 109316 3392
rect 109368 3380 109374 3392
rect 111058 3380 111064 3392
rect 109368 3352 111064 3380
rect 109368 3340 109374 3352
rect 111058 3340 111064 3352
rect 111116 3340 111122 3392
rect 182818 3340 182824 3392
rect 182876 3380 182882 3392
rect 190426 3380 190454 3420
rect 207382 3408 207388 3420
rect 207440 3408 207446 3460
rect 210418 3408 210424 3460
rect 210476 3448 210482 3460
rect 218054 3448 218060 3460
rect 210476 3420 218060 3448
rect 210476 3408 210482 3420
rect 218054 3408 218060 3420
rect 218112 3408 218118 3460
rect 219406 3420 354674 3448
rect 182876 3352 190454 3380
rect 182876 3340 182882 3352
rect 215938 3340 215944 3392
rect 215996 3380 216002 3392
rect 219406 3380 219434 3420
rect 215996 3352 219434 3380
rect 215996 3340 216002 3352
rect 258718 3340 258724 3392
rect 258776 3380 258782 3392
rect 259454 3380 259460 3392
rect 258776 3352 259460 3380
rect 258776 3340 258782 3352
rect 259454 3340 259460 3352
rect 259512 3340 259518 3392
rect 260006 3340 260012 3392
rect 260064 3380 260070 3392
rect 264146 3380 264152 3392
rect 260064 3352 264152 3380
rect 260064 3340 260070 3352
rect 264146 3340 264152 3352
rect 264204 3340 264210 3392
rect 271138 3340 271144 3392
rect 271196 3380 271202 3392
rect 274818 3380 274824 3392
rect 271196 3352 274824 3380
rect 271196 3340 271202 3352
rect 274818 3340 274824 3352
rect 274876 3340 274882 3392
rect 278038 3340 278044 3392
rect 278096 3380 278102 3392
rect 281902 3380 281908 3392
rect 278096 3352 281908 3380
rect 278096 3340 278102 3352
rect 281902 3340 281908 3352
rect 281960 3340 281966 3392
rect 309870 3340 309876 3392
rect 309928 3380 309934 3392
rect 313826 3380 313832 3392
rect 309928 3352 313832 3380
rect 309928 3340 309934 3352
rect 313826 3340 313832 3352
rect 313884 3340 313890 3392
rect 320818 3380 320824 3392
rect 313936 3352 320824 3380
rect 18230 3272 18236 3324
rect 18288 3312 18294 3324
rect 22738 3312 22744 3324
rect 18288 3284 22744 3312
rect 18288 3272 18294 3284
rect 22738 3272 22744 3284
rect 22796 3272 22802 3324
rect 77386 3272 77392 3324
rect 77444 3312 77450 3324
rect 79318 3312 79324 3324
rect 77444 3284 79324 3312
rect 77444 3272 77450 3284
rect 79318 3272 79324 3284
rect 79376 3272 79382 3324
rect 126974 3272 126980 3324
rect 127032 3312 127038 3324
rect 128998 3312 129004 3324
rect 127032 3284 129004 3312
rect 127032 3272 127038 3284
rect 128998 3272 129004 3284
rect 129056 3272 129062 3324
rect 135254 3272 135260 3324
rect 135312 3312 135318 3324
rect 137278 3312 137284 3324
rect 135312 3284 137284 3312
rect 135312 3272 135318 3284
rect 137278 3272 137284 3284
rect 137336 3272 137342 3324
rect 214558 3272 214564 3324
rect 214616 3312 214622 3324
rect 215662 3312 215668 3324
rect 214616 3284 215668 3312
rect 214616 3272 214622 3284
rect 215662 3272 215668 3284
rect 215720 3272 215726 3324
rect 309778 3272 309784 3324
rect 309836 3312 309842 3324
rect 313936 3312 313964 3352
rect 320818 3340 320824 3352
rect 320876 3340 320882 3392
rect 332686 3340 332692 3392
rect 332744 3380 332750 3392
rect 333882 3380 333888 3392
rect 332744 3352 333888 3380
rect 332744 3340 332750 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 354646 3380 354674 3420
rect 357526 3408 357532 3460
rect 357584 3448 357590 3460
rect 358722 3448 358728 3460
rect 357584 3420 358728 3448
rect 357584 3408 357590 3420
rect 358722 3408 358728 3420
rect 358780 3408 358786 3460
rect 390554 3408 390560 3460
rect 390612 3448 390618 3460
rect 391842 3448 391848 3460
rect 390612 3420 391848 3448
rect 390612 3408 390618 3420
rect 391842 3408 391848 3420
rect 391900 3408 391906 3460
rect 393286 3420 412634 3448
rect 363506 3380 363512 3392
rect 354646 3352 363512 3380
rect 363506 3340 363512 3352
rect 363564 3340 363570 3392
rect 387058 3340 387064 3392
rect 387116 3380 387122 3392
rect 393286 3380 393314 3420
rect 387116 3352 393314 3380
rect 387116 3340 387122 3352
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 309836 3284 313964 3312
rect 412606 3312 412634 3420
rect 415228 3380 415256 3488
rect 415394 3476 415400 3528
rect 415452 3516 415458 3528
rect 416682 3516 416688 3528
rect 415452 3488 416688 3516
rect 415452 3476 415458 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 422938 3476 422944 3528
rect 422996 3516 423002 3528
rect 423766 3516 423772 3528
rect 422996 3488 423772 3516
rect 422996 3476 423002 3488
rect 423766 3476 423772 3488
rect 423824 3476 423830 3528
rect 432046 3476 432052 3528
rect 432104 3516 432110 3528
rect 433242 3516 433248 3528
rect 432104 3488 433248 3516
rect 432104 3476 432110 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 436738 3476 436744 3528
rect 436796 3516 436802 3528
rect 437934 3516 437940 3528
rect 436796 3488 437940 3516
rect 436796 3476 436802 3488
rect 437934 3476 437940 3488
rect 437992 3476 437998 3528
rect 440234 3476 440240 3528
rect 440292 3516 440298 3528
rect 441522 3516 441528 3528
rect 440292 3488 441528 3516
rect 440292 3476 440298 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 447778 3476 447784 3528
rect 447836 3516 447842 3528
rect 448606 3516 448612 3528
rect 447836 3488 448612 3516
rect 447836 3476 447842 3488
rect 448606 3476 448612 3488
rect 448664 3476 448670 3528
rect 456886 3476 456892 3528
rect 456944 3516 456950 3528
rect 458082 3516 458088 3528
rect 456944 3488 458088 3516
rect 456944 3476 456950 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 465074 3476 465080 3528
rect 465132 3516 465138 3528
rect 465902 3516 465908 3528
rect 465132 3488 465908 3516
rect 465132 3476 465138 3488
rect 465902 3476 465908 3488
rect 465960 3476 465966 3528
rect 468478 3476 468484 3528
rect 468536 3516 468542 3528
rect 469858 3516 469864 3528
rect 468536 3488 469864 3516
rect 468536 3476 468542 3488
rect 469858 3476 469864 3488
rect 469916 3476 469922 3528
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 473446 3516 473452 3528
rect 472676 3488 473452 3516
rect 472676 3476 472682 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 520918 3476 520924 3528
rect 520976 3516 520982 3528
rect 521838 3516 521844 3528
rect 520976 3488 521844 3516
rect 520976 3476 520982 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 522298 3476 522304 3528
rect 522356 3516 522362 3528
rect 523034 3516 523040 3528
rect 522356 3488 523040 3516
rect 522356 3476 522362 3488
rect 523034 3476 523040 3488
rect 523092 3476 523098 3528
rect 527910 3476 527916 3528
rect 527968 3516 527974 3528
rect 552658 3516 552664 3528
rect 527968 3488 552664 3516
rect 527968 3476 527974 3488
rect 552658 3476 552664 3488
rect 552716 3476 552722 3528
rect 566826 3448 566832 3460
rect 422266 3420 566832 3448
rect 421374 3380 421380 3392
rect 415228 3352 421380 3380
rect 421374 3340 421380 3352
rect 421432 3340 421438 3392
rect 422266 3312 422294 3420
rect 566826 3408 566832 3420
rect 566884 3408 566890 3460
rect 412606 3284 422294 3312
rect 309836 3272 309842 3284
rect 27706 3204 27712 3256
rect 27764 3244 27770 3256
rect 31018 3244 31024 3256
rect 27764 3216 31024 3244
rect 27764 3204 27770 3216
rect 31018 3204 31024 3216
rect 31076 3204 31082 3256
rect 163682 3204 163688 3256
rect 163740 3244 163746 3256
rect 166350 3244 166356 3256
rect 163740 3216 166356 3244
rect 163740 3204 163746 3216
rect 166350 3204 166356 3216
rect 166408 3204 166414 3256
rect 175274 3204 175280 3256
rect 175332 3244 175338 3256
rect 179046 3244 179052 3256
rect 175332 3216 179052 3244
rect 175332 3204 175338 3216
rect 179046 3204 179052 3216
rect 179104 3204 179110 3256
rect 314010 3204 314016 3256
rect 314068 3244 314074 3256
rect 318518 3244 318524 3256
rect 314068 3216 318524 3244
rect 314068 3204 314074 3216
rect 318518 3204 318524 3216
rect 318576 3204 318582 3256
rect 216582 3136 216588 3188
rect 216640 3176 216646 3188
rect 219250 3176 219256 3188
rect 216640 3148 219256 3176
rect 216640 3136 216646 3148
rect 219250 3136 219256 3148
rect 219308 3136 219314 3188
rect 282178 3136 282184 3188
rect 282236 3176 282242 3188
rect 285398 3176 285404 3188
rect 282236 3148 285404 3176
rect 282236 3136 282242 3148
rect 285398 3136 285404 3148
rect 285456 3136 285462 3188
rect 307202 3136 307208 3188
rect 307260 3176 307266 3188
rect 310238 3176 310244 3188
rect 307260 3148 310244 3176
rect 307260 3136 307266 3148
rect 310238 3136 310244 3148
rect 310296 3136 310302 3188
rect 331858 3136 331864 3188
rect 331916 3176 331922 3188
rect 335078 3176 335084 3188
rect 331916 3148 335084 3176
rect 331916 3136 331922 3148
rect 335078 3136 335084 3148
rect 335136 3136 335142 3188
rect 12342 3068 12348 3120
rect 12400 3108 12406 3120
rect 13078 3108 13084 3120
rect 12400 3080 13084 3108
rect 12400 3068 12406 3080
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 229738 3068 229744 3120
rect 229796 3108 229802 3120
rect 232222 3108 232228 3120
rect 229796 3080 232228 3108
rect 229796 3068 229802 3080
rect 232222 3068 232228 3080
rect 232280 3068 232286 3120
rect 247678 3068 247684 3120
rect 247736 3108 247742 3120
rect 248782 3108 248788 3120
rect 247736 3080 248788 3108
rect 247736 3068 247742 3080
rect 248782 3068 248788 3080
rect 248840 3068 248846 3120
rect 542998 3068 543004 3120
rect 543056 3108 543062 3120
rect 545482 3108 545488 3120
rect 543056 3080 545488 3108
rect 543056 3068 543062 3080
rect 545482 3068 545488 3080
rect 545540 3068 545546 3120
rect 41874 3000 41880 3052
rect 41932 3040 41938 3052
rect 44818 3040 44824 3052
rect 41932 3012 44824 3040
rect 41932 3000 41938 3012
rect 44818 3000 44824 3012
rect 44876 3000 44882 3052
rect 167178 3000 167184 3052
rect 167236 3040 167242 3052
rect 171410 3040 171416 3052
rect 167236 3012 171416 3040
rect 167236 3000 167242 3012
rect 171410 3000 171416 3012
rect 171468 3000 171474 3052
rect 181438 3000 181444 3052
rect 181496 3040 181502 3052
rect 189718 3040 189724 3052
rect 181496 3012 189724 3040
rect 181496 3000 181502 3012
rect 189718 3000 189724 3012
rect 189776 3000 189782 3052
rect 196618 3000 196624 3052
rect 196676 3040 196682 3052
rect 197906 3040 197912 3052
rect 196676 3012 197912 3040
rect 196676 3000 196682 3012
rect 197906 3000 197912 3012
rect 197964 3000 197970 3052
rect 200758 3000 200764 3052
rect 200816 3040 200822 3052
rect 202690 3040 202696 3052
rect 200816 3012 202696 3040
rect 200816 3000 200822 3012
rect 202690 3000 202696 3012
rect 202748 3000 202754 3052
rect 289170 3000 289176 3052
rect 289228 3040 289234 3052
rect 296070 3040 296076 3052
rect 289228 3012 296076 3040
rect 289228 3000 289234 3012
rect 296070 3000 296076 3012
rect 296128 3000 296134 3052
rect 307018 3000 307024 3052
rect 307076 3040 307082 3052
rect 315022 3040 315028 3052
rect 307076 3012 315028 3040
rect 307076 3000 307082 3012
rect 315022 3000 315028 3012
rect 315080 3000 315086 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 536190 3000 536196 3052
rect 536248 3040 536254 3052
rect 540790 3040 540796 3052
rect 536248 3012 540796 3040
rect 536248 3000 536254 3012
rect 540790 3000 540796 3012
rect 540848 3000 540854 3052
rect 291838 2932 291844 2984
rect 291896 2972 291902 2984
rect 293678 2972 293684 2984
rect 291896 2944 293684 2972
rect 291896 2932 291902 2944
rect 293678 2932 293684 2944
rect 293736 2932 293742 2984
rect 548518 2932 548524 2984
rect 548576 2972 548582 2984
rect 550266 2972 550272 2984
rect 548576 2944 550272 2972
rect 548576 2932 548582 2944
rect 550266 2932 550272 2944
rect 550324 2932 550330 2984
rect 115198 2864 115204 2916
rect 115256 2904 115262 2916
rect 116578 2904 116584 2916
rect 115256 2876 116584 2904
rect 115256 2864 115262 2876
rect 116578 2864 116584 2876
rect 116636 2864 116642 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 348792 700340 348844 700392
rect 364524 700340 364576 700392
rect 24308 700272 24360 700324
rect 280804 700272 280856 700324
rect 283840 700272 283892 700324
rect 304264 700272 304316 700324
rect 332508 700272 332560 700324
rect 364432 700272 364484 700324
rect 218980 699660 219032 699712
rect 220084 699660 220136 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 363604 698640 363656 698692
rect 364984 698640 365036 698692
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 378784 696940 378836 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 369860 683136 369912 683188
rect 3516 670692 3568 670744
rect 298744 670692 298796 670744
rect 360108 670692 360160 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 10324 656888 10376 656940
rect 359464 643084 359516 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 371240 632068 371292 632120
rect 359556 630640 359608 630692
rect 579988 630640 580040 630692
rect 3148 618264 3200 618316
rect 311164 618264 311216 618316
rect 382924 616836 382976 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 180064 605820 180116 605872
rect 367744 590656 367796 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 372620 579640 372672 579692
rect 358084 576852 358136 576904
rect 580172 576852 580224 576904
rect 376024 563048 376076 563100
rect 580172 563048 580224 563100
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 377404 536800 377456 536852
rect 579896 536800 579948 536852
rect 2964 527144 3016 527196
rect 374000 527144 374052 527196
rect 392584 524424 392636 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 262864 514768 262916 514820
rect 361488 511232 361540 511284
rect 580264 511232 580316 511284
rect 3056 500964 3108 501016
rect 51724 500964 51776 501016
rect 355324 484372 355376 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 374460 474716 374512 474768
rect 363972 473968 364024 474020
rect 412640 473968 412692 474020
rect 356704 472608 356756 472660
rect 392584 472608 392636 472660
rect 367836 470568 367888 470620
rect 580080 470568 580132 470620
rect 360844 469820 360896 469872
rect 527180 469820 527232 469872
rect 357716 468460 357768 468512
rect 367744 468460 367796 468512
rect 40040 467100 40092 467152
rect 368572 467100 368624 467152
rect 104900 465672 104952 465724
rect 273260 465672 273312 465724
rect 362224 465672 362276 465724
rect 477500 465672 477552 465724
rect 273260 465060 273312 465112
rect 274548 465060 274600 465112
rect 368480 465060 368532 465112
rect 169760 464312 169812 464364
rect 281448 464312 281500 464364
rect 362316 464312 362368 464364
rect 542360 464312 542412 464364
rect 281448 463700 281500 463752
rect 367284 463700 367336 463752
rect 356796 462952 356848 463004
rect 377404 462952 377456 463004
rect 3516 462340 3568 462392
rect 315304 462340 315356 462392
rect 364156 461660 364208 461712
rect 396724 461660 396776 461712
rect 234620 461592 234672 461644
rect 365720 461592 365772 461644
rect 357348 460232 357400 460284
rect 367836 460232 367888 460284
rect 363144 460164 363196 460216
rect 429200 460164 429252 460216
rect 361120 458804 361172 458856
rect 558920 458804 558972 458856
rect 334716 457240 334768 457292
rect 373540 457240 373592 457292
rect 323768 457172 323820 457224
rect 384212 457172 384264 457224
rect 320916 457104 320968 457156
rect 381084 457104 381136 457156
rect 315304 457036 315356 457088
rect 375748 457036 375800 457088
rect 320824 456968 320876 457020
rect 381268 456968 381320 457020
rect 311164 456900 311216 456952
rect 311808 456900 311860 456952
rect 372712 456900 372764 456952
rect 298744 456764 298796 456816
rect 299388 456764 299440 456816
rect 371424 456832 371476 456884
rect 355968 456764 356020 456816
rect 580172 456764 580224 456816
rect 357624 456084 357676 456136
rect 382924 456084 382976 456136
rect 362868 456016 362920 456068
rect 462320 456016 462372 456068
rect 361672 455948 361724 456000
rect 362316 455948 362368 456000
rect 334624 455880 334676 455932
rect 355508 455880 355560 455932
rect 332140 455812 332192 455864
rect 356152 455812 356204 455864
rect 357348 455812 357400 455864
rect 332048 455744 332100 455796
rect 359556 455744 359608 455796
rect 333336 455676 333388 455728
rect 361672 455676 361724 455728
rect 332232 455608 332284 455660
rect 364432 455608 364484 455660
rect 333428 455540 333480 455592
rect 380164 455540 380216 455592
rect 302884 455472 302936 455524
rect 362224 455472 362276 455524
rect 322296 455404 322348 455456
rect 383108 455404 383160 455456
rect 281356 454928 281408 454980
rect 351920 454928 351972 454980
rect 319536 454860 319588 454912
rect 379796 454860 379848 454912
rect 294696 454792 294748 454844
rect 354680 454792 354732 454844
rect 357440 454792 357492 454844
rect 376024 454792 376076 454844
rect 337936 454724 337988 454776
rect 357624 454724 357676 454776
rect 358452 454724 358504 454776
rect 337292 454656 337344 454708
rect 362040 454656 362092 454708
rect 494060 454656 494112 454708
rect 337384 454588 337436 454640
rect 363144 454588 363196 454640
rect 319628 454520 319680 454572
rect 376760 454520 376812 454572
rect 319720 454452 319772 454504
rect 378692 454452 378744 454504
rect 293868 454384 293920 454436
rect 353300 454384 353352 454436
rect 318248 454316 318300 454368
rect 378324 454316 378376 454368
rect 316868 454248 316920 454300
rect 376944 454248 376996 454300
rect 340696 454180 340748 454232
rect 357440 454180 357492 454232
rect 336464 454112 336516 454164
rect 355048 454112 355100 454164
rect 337476 454044 337528 454096
rect 374276 454044 374328 454096
rect 323584 453568 323636 453620
rect 383844 453568 383896 453620
rect 318064 453500 318116 453552
rect 378416 453500 378468 453552
rect 335268 453432 335320 453484
rect 359096 453432 359148 453484
rect 361396 453432 361448 453484
rect 378784 453432 378836 453484
rect 299480 453364 299532 453416
rect 365076 453364 365128 453416
rect 356244 453296 356296 453348
rect 580356 453296 580408 453348
rect 335176 453228 335228 453280
rect 362408 453228 362460 453280
rect 362868 453228 362920 453280
rect 315396 453160 315448 453212
rect 367100 453160 367152 453212
rect 316684 453092 316736 453144
rect 371332 453092 371384 453144
rect 318156 453024 318208 453076
rect 377220 453024 377272 453076
rect 316776 452956 316828 453008
rect 376116 452956 376168 453008
rect 294788 452888 294840 452940
rect 354128 452888 354180 452940
rect 322204 452820 322256 452872
rect 381636 452820 381688 452872
rect 324964 452752 325016 452804
rect 385040 452752 385092 452804
rect 341984 452684 342036 452736
rect 353024 452684 353076 452736
rect 340052 452616 340104 452668
rect 356244 452616 356296 452668
rect 355416 452548 355468 452600
rect 355968 452548 356020 452600
rect 376760 452548 376812 452600
rect 379060 452548 379112 452600
rect 278596 452140 278648 452192
rect 348516 452140 348568 452192
rect 294604 452072 294656 452124
rect 350632 452072 350684 452124
rect 340144 452004 340196 452056
rect 385684 452004 385736 452056
rect 308496 451936 308548 451988
rect 367192 451936 367244 451988
rect 371332 451936 371384 451988
rect 376760 451936 376812 451988
rect 300124 451868 300176 451920
rect 355416 451868 355468 451920
rect 363328 451868 363380 451920
rect 365720 451868 365772 451920
rect 366180 451868 366232 451920
rect 342168 451800 342220 451852
rect 353668 451800 353720 451852
rect 363604 451800 363656 451852
rect 364064 451800 364116 451852
rect 342352 451732 342404 451784
rect 365812 451732 365864 451784
rect 341524 451664 341576 451716
rect 374644 451664 374696 451716
rect 340972 451596 341024 451648
rect 309784 451528 309836 451580
rect 352656 451528 352708 451580
rect 354588 451528 354640 451580
rect 337568 451460 337620 451512
rect 349252 451460 349304 451512
rect 384580 451528 384632 451580
rect 366548 451460 366600 451512
rect 341708 451392 341760 451444
rect 382372 451392 382424 451444
rect 339408 451324 339460 451376
rect 352564 451324 352616 451376
rect 352656 451324 352708 451376
rect 364708 451324 364760 451376
rect 367100 451324 367152 451376
rect 375380 451324 375432 451376
rect 338856 451256 338908 451308
rect 351460 451256 351512 451308
rect 355048 451256 355100 451308
rect 357440 451256 357492 451308
rect 365720 451256 365772 451308
rect 369952 451256 370004 451308
rect 297456 450780 297508 450832
rect 357716 450780 357768 450832
rect 300308 450712 300360 450764
rect 360200 450712 360252 450764
rect 361396 450712 361448 450764
rect 266360 450644 266412 450696
rect 305000 450644 305052 450696
rect 321008 450644 321060 450696
rect 380532 450644 380584 450696
rect 201500 450576 201552 450628
rect 136640 450508 136692 450560
rect 319444 450576 319496 450628
rect 379428 450576 379480 450628
rect 306380 450508 306432 450560
rect 354588 450508 354640 450560
rect 357440 450508 357492 450560
rect 580264 450508 580316 450560
rect 323676 450440 323728 450492
rect 382740 450440 382792 450492
rect 314016 450372 314068 450424
rect 373172 450372 373224 450424
rect 301504 450304 301556 450356
rect 361028 450304 361080 450356
rect 297364 450236 297416 450288
rect 356888 450236 356940 450288
rect 279884 450168 279936 450220
rect 367882 450168 367934 450220
rect 371240 450168 371292 450220
rect 371700 450168 371752 450220
rect 338764 450100 338816 450152
rect 349114 450100 349166 450152
rect 354128 450100 354180 450152
rect 388444 450100 388496 450152
rect 305000 450032 305052 450084
rect 365444 450032 365496 450084
rect 340328 449964 340380 450016
rect 372068 449964 372120 450016
rect 340788 449896 340840 449948
rect 348148 449896 348200 449948
rect 354864 449896 354916 449948
rect 389824 449896 389876 449948
rect 363328 449556 363380 449608
rect 307024 449284 307076 449336
rect 342444 449420 342496 449472
rect 349620 449420 349672 449472
rect 342076 449284 342128 449336
rect 351092 449420 351144 449472
rect 369860 449420 369912 449472
rect 370596 449420 370648 449472
rect 358084 449352 358136 449404
rect 304356 449216 304408 449268
rect 330208 449216 330260 449268
rect 298744 449148 298796 449200
rect 330208 449080 330260 449132
rect 363972 449352 364024 449404
rect 3148 448536 3200 448588
rect 8944 448536 8996 448588
rect 277768 448536 277820 448588
rect 342444 448536 342496 448588
rect 325056 445000 325108 445052
rect 340972 445000 341024 445052
rect 322388 438132 322440 438184
rect 340972 438132 341024 438184
rect 287704 435344 287756 435396
rect 340880 435344 340932 435396
rect 389824 431876 389876 431928
rect 580172 431876 580224 431928
rect 3516 422288 3568 422340
rect 311164 422288 311216 422340
rect 289728 418752 289780 418804
rect 337568 418752 337620 418804
rect 262864 417392 262916 417444
rect 315488 417392 315540 417444
rect 8944 416712 8996 416764
rect 314752 416712 314804 416764
rect 315396 416712 315448 416764
rect 311164 415420 311216 415472
rect 316776 415420 316828 415472
rect 51724 414672 51776 414724
rect 313924 414672 313976 414724
rect 313924 413924 313976 413976
rect 337476 413924 337528 413976
rect 4804 413856 4856 413908
rect 313280 413856 313332 413908
rect 314016 413856 314068 413908
rect 180064 411884 180116 411936
rect 311900 411884 311952 411936
rect 311900 411204 311952 411256
rect 312636 411204 312688 411256
rect 340328 411204 340380 411256
rect 10324 410524 10376 410576
rect 311256 410524 311308 410576
rect 286416 409096 286468 409148
rect 340236 409096 340288 409148
rect 326344 407736 326396 407788
rect 340144 407736 340196 407788
rect 291936 406444 291988 406496
rect 338856 406444 338908 406496
rect 88340 406376 88392 406428
rect 309968 406376 310020 406428
rect 4160 405628 4212 405680
rect 316040 405628 316092 405680
rect 316868 405628 316920 405680
rect 388996 405628 389048 405680
rect 580172 405628 580224 405680
rect 309968 405560 310020 405612
rect 334808 405560 334860 405612
rect 315488 404268 315540 404320
rect 340972 404268 341024 404320
rect 299388 403588 299440 403640
rect 310520 403588 310572 403640
rect 3424 402228 3476 402280
rect 313280 402228 313332 402280
rect 316132 401616 316184 401668
rect 316776 401616 316828 401668
rect 313280 401548 313332 401600
rect 314016 401548 314068 401600
rect 334716 401548 334768 401600
rect 341800 400936 341852 400988
rect 341432 400800 341484 400852
rect 341524 400800 341576 400852
rect 342260 400800 342312 400852
rect 281264 400528 281316 400580
rect 341892 400528 341944 400580
rect 279976 400460 280028 400512
rect 342260 400460 342312 400512
rect 271696 400392 271748 400444
rect 277124 400324 277176 400376
rect 341432 400324 341484 400376
rect 281080 400256 281132 400308
rect 341892 400256 341944 400308
rect 342260 400324 342312 400376
rect 274272 400188 274324 400240
rect 341340 400120 341392 400172
rect 331864 399644 331916 399696
rect 339868 400052 339920 400104
rect 341616 400052 341668 400104
rect 341524 399916 341576 399968
rect 342352 399848 342404 399900
rect 342582 399848 342634 399900
rect 342766 399848 342818 399900
rect 343686 399848 343738 399900
rect 340328 399712 340380 399764
rect 341248 399644 341300 399696
rect 344054 399848 344106 399900
rect 344146 399848 344198 399900
rect 344514 399848 344566 399900
rect 344606 399848 344658 399900
rect 344790 399848 344842 399900
rect 345342 399848 345394 399900
rect 346170 399848 346222 399900
rect 346354 399848 346406 399900
rect 346722 399848 346774 399900
rect 346998 399848 347050 399900
rect 347182 399848 347234 399900
rect 347366 399848 347418 399900
rect 347826 399848 347878 399900
rect 347918 399848 347970 399900
rect 348194 399848 348246 399900
rect 348286 399848 348338 399900
rect 310060 399576 310112 399628
rect 341800 399576 341852 399628
rect 344422 399780 344474 399832
rect 344376 399644 344428 399696
rect 344192 399576 344244 399628
rect 344744 399712 344796 399764
rect 344652 399644 344704 399696
rect 345986 399780 346038 399832
rect 311164 399508 311216 399560
rect 342260 399508 342312 399560
rect 342812 399508 342864 399560
rect 343824 399508 343876 399560
rect 344008 399508 344060 399560
rect 345296 399508 345348 399560
rect 345940 399576 345992 399628
rect 345572 399508 345624 399560
rect 347550 399780 347602 399832
rect 347642 399780 347694 399832
rect 347228 399712 347280 399764
rect 347320 399712 347372 399764
rect 347504 399644 347556 399696
rect 347780 399712 347832 399764
rect 348240 399712 348292 399764
rect 348838 399848 348890 399900
rect 350586 399848 350638 399900
rect 350678 399848 350730 399900
rect 350954 399848 351006 399900
rect 351414 399848 351466 399900
rect 348746 399780 348798 399832
rect 347872 399644 347924 399696
rect 348148 399644 348200 399696
rect 348332 399644 348384 399696
rect 347596 399576 347648 399628
rect 349022 399780 349074 399832
rect 349482 399780 349534 399832
rect 349574 399780 349626 399832
rect 349666 399780 349718 399832
rect 349850 399780 349902 399832
rect 349942 399780 349994 399832
rect 350126 399780 350178 399832
rect 350310 399780 350362 399832
rect 350494 399780 350546 399832
rect 348792 399644 348844 399696
rect 349068 399644 349120 399696
rect 349160 399644 349212 399696
rect 349528 399644 349580 399696
rect 348976 399576 349028 399628
rect 349436 399576 349488 399628
rect 312728 399440 312780 399492
rect 277216 399372 277268 399424
rect 344560 399440 344612 399492
rect 347136 399508 347188 399560
rect 348424 399508 348476 399560
rect 348516 399508 348568 399560
rect 349804 399508 349856 399560
rect 346308 399440 346360 399492
rect 348056 399440 348108 399492
rect 350080 399644 350132 399696
rect 275928 399304 275980 399356
rect 346768 399372 346820 399424
rect 346952 399372 347004 399424
rect 349896 399440 349948 399492
rect 350264 399440 350316 399492
rect 350632 399712 350684 399764
rect 350724 399712 350776 399764
rect 351230 399780 351282 399832
rect 350448 399576 350500 399628
rect 351000 399576 351052 399628
rect 351690 399848 351742 399900
rect 351874 399848 351926 399900
rect 351966 399848 352018 399900
rect 351644 399712 351696 399764
rect 351736 399644 351788 399696
rect 352242 399848 352294 399900
rect 352426 399848 352478 399900
rect 352518 399848 352570 399900
rect 352150 399780 352202 399832
rect 352104 399644 352156 399696
rect 352196 399576 352248 399628
rect 352380 399576 352432 399628
rect 351184 399508 351236 399560
rect 352012 399508 352064 399560
rect 352472 399440 352524 399492
rect 353254 399848 353306 399900
rect 353300 399644 353352 399696
rect 353622 399848 353674 399900
rect 353806 399848 353858 399900
rect 353898 399780 353950 399832
rect 352748 399508 352800 399560
rect 349620 399372 349672 399424
rect 350908 399372 350960 399424
rect 353668 399576 353720 399628
rect 353852 399508 353904 399560
rect 354266 399848 354318 399900
rect 354082 399780 354134 399832
rect 354220 399576 354272 399628
rect 354128 399508 354180 399560
rect 353944 399440 353996 399492
rect 354450 399780 354502 399832
rect 354726 399848 354778 399900
rect 354910 399848 354962 399900
rect 354634 399780 354686 399832
rect 354680 399644 354732 399696
rect 355094 399780 355146 399832
rect 354772 399576 354824 399628
rect 354864 399576 354916 399628
rect 354404 399372 354456 399424
rect 354772 399372 354824 399424
rect 355554 399848 355606 399900
rect 355922 399848 355974 399900
rect 355508 399644 355560 399696
rect 355416 399508 355468 399560
rect 355232 399440 355284 399492
rect 354588 399304 354640 399356
rect 355140 399304 355192 399356
rect 355876 399508 355928 399560
rect 356290 399848 356342 399900
rect 356566 399848 356618 399900
rect 356842 399848 356894 399900
rect 357118 399848 357170 399900
rect 356152 399508 356204 399560
rect 356612 399712 356664 399764
rect 356520 399508 356572 399560
rect 356336 399440 356388 399492
rect 356428 399440 356480 399492
rect 356796 399440 356848 399492
rect 355876 399372 355928 399424
rect 357348 399508 357400 399560
rect 355692 399304 355744 399356
rect 356244 399304 356296 399356
rect 356428 399304 356480 399356
rect 357578 399848 357630 399900
rect 357762 399848 357814 399900
rect 357854 399848 357906 399900
rect 357946 399848 357998 399900
rect 358222 399848 358274 399900
rect 358406 399848 358458 399900
rect 358682 399848 358734 399900
rect 358866 399848 358918 399900
rect 359234 399848 359286 399900
rect 359418 399848 359470 399900
rect 359602 399848 359654 399900
rect 360062 399848 360114 399900
rect 360246 399848 360298 399900
rect 360338 399848 360390 399900
rect 360706 399848 360758 399900
rect 360798 399848 360850 399900
rect 357624 399508 357676 399560
rect 348424 399236 348476 399288
rect 357164 399236 357216 399288
rect 357992 399644 358044 399696
rect 358268 399644 358320 399696
rect 358498 399780 358550 399832
rect 358544 399644 358596 399696
rect 358452 399576 358504 399628
rect 358176 399508 358228 399560
rect 359142 399780 359194 399832
rect 359280 399576 359332 399628
rect 359694 399780 359746 399832
rect 359786 399780 359838 399832
rect 359878 399780 359930 399832
rect 359648 399644 359700 399696
rect 359740 399576 359792 399628
rect 359832 399576 359884 399628
rect 359372 399508 359424 399560
rect 359464 399508 359516 399560
rect 360016 399508 360068 399560
rect 360108 399440 360160 399492
rect 360292 399576 360344 399628
rect 360660 399440 360712 399492
rect 361074 399848 361126 399900
rect 361166 399848 361218 399900
rect 361258 399848 361310 399900
rect 361534 399848 361586 399900
rect 360936 399508 360988 399560
rect 360844 399440 360896 399492
rect 359096 399372 359148 399424
rect 358728 399304 358780 399356
rect 358084 399236 358136 399288
rect 360752 399236 360804 399288
rect 361442 399780 361494 399832
rect 361626 399780 361678 399832
rect 361902 399848 361954 399900
rect 361396 399508 361448 399560
rect 361580 399508 361632 399560
rect 361764 399508 361816 399560
rect 362730 399848 362782 399900
rect 362914 399848 362966 399900
rect 361994 399780 362046 399832
rect 362270 399780 362322 399832
rect 362362 399780 362414 399832
rect 362454 399780 362506 399832
rect 362132 399508 362184 399560
rect 361488 399440 361540 399492
rect 361672 399372 361724 399424
rect 362316 399644 362368 399696
rect 362592 399644 362644 399696
rect 362408 399576 362460 399628
rect 362500 399508 362552 399560
rect 363098 399848 363150 399900
rect 363558 399848 363610 399900
rect 363650 399848 363702 399900
rect 364018 399848 364070 399900
rect 364294 399848 364346 399900
rect 364386 399848 364438 399900
rect 364570 399848 364622 399900
rect 365030 399848 365082 399900
rect 365214 399848 365266 399900
rect 365306 399848 365358 399900
rect 365490 399848 365542 399900
rect 366042 399848 366094 399900
rect 366134 399848 366186 399900
rect 366226 399848 366278 399900
rect 363052 399508 363104 399560
rect 363236 399372 363288 399424
rect 363328 399372 363380 399424
rect 363972 399644 364024 399696
rect 364432 399644 364484 399696
rect 364340 399576 364392 399628
rect 364064 399508 364116 399560
rect 364754 399780 364806 399832
rect 361304 399304 361356 399356
rect 364892 399508 364944 399560
rect 365260 399712 365312 399764
rect 365168 399644 365220 399696
rect 365444 399644 365496 399696
rect 365536 399576 365588 399628
rect 366088 399576 366140 399628
rect 365720 399508 365772 399560
rect 365812 399508 365864 399560
rect 387800 400460 387852 400512
rect 392124 400460 392176 400512
rect 390192 400324 390244 400376
rect 394792 400324 394844 400376
rect 366594 399848 366646 399900
rect 366870 399848 366922 399900
rect 366548 399712 366600 399764
rect 366364 399644 366416 399696
rect 366456 399508 366508 399560
rect 366732 399712 366784 399764
rect 366824 399712 366876 399764
rect 366640 399576 366692 399628
rect 366732 399508 366784 399560
rect 366548 399440 366600 399492
rect 367606 399848 367658 399900
rect 368710 399848 368762 399900
rect 368802 399848 368854 399900
rect 369170 399848 369222 399900
rect 369906 399848 369958 399900
rect 370090 399848 370142 399900
rect 370366 399848 370418 399900
rect 370734 399848 370786 399900
rect 370918 399848 370970 399900
rect 371286 399848 371338 399900
rect 371654 399848 371706 399900
rect 367422 399780 367474 399832
rect 367468 399644 367520 399696
rect 368250 399780 368302 399832
rect 368342 399780 368394 399832
rect 367928 399576 367980 399628
rect 368204 399576 368256 399628
rect 368664 399644 368716 399696
rect 368296 399508 368348 399560
rect 368940 399508 368992 399560
rect 367376 399372 367428 399424
rect 367560 399372 367612 399424
rect 364064 399236 364116 399288
rect 367560 399236 367612 399288
rect 337752 399168 337804 399220
rect 348700 399168 348752 399220
rect 349620 399168 349672 399220
rect 353484 399168 353536 399220
rect 354036 399168 354088 399220
rect 368388 399236 368440 399288
rect 369676 399372 369728 399424
rect 369998 399780 370050 399832
rect 370044 399508 370096 399560
rect 369584 399304 369636 399356
rect 370228 399440 370280 399492
rect 370550 399780 370602 399832
rect 370504 399576 370556 399628
rect 370688 399576 370740 399628
rect 370596 399440 370648 399492
rect 370688 399372 370740 399424
rect 371332 399712 371384 399764
rect 371700 399712 371752 399764
rect 370964 399508 371016 399560
rect 371056 399372 371108 399424
rect 371516 399304 371568 399356
rect 372022 399848 372074 399900
rect 372114 399848 372166 399900
rect 372298 399848 372350 399900
rect 372666 399848 372718 399900
rect 372850 399848 372902 399900
rect 373034 399848 373086 399900
rect 373218 399848 373270 399900
rect 372482 399780 372534 399832
rect 372344 399644 372396 399696
rect 372436 399644 372488 399696
rect 372528 399576 372580 399628
rect 371976 399508 372028 399560
rect 372804 399644 372856 399696
rect 373494 399780 373546 399832
rect 373586 399780 373638 399832
rect 373678 399780 373730 399832
rect 373770 399780 373822 399832
rect 373862 399780 373914 399832
rect 373540 399576 373592 399628
rect 373448 399508 373500 399560
rect 373908 399644 373960 399696
rect 373724 399576 373776 399628
rect 374230 399848 374282 399900
rect 374414 399848 374466 399900
rect 374690 399848 374742 399900
rect 374598 399780 374650 399832
rect 374276 399576 374328 399628
rect 373816 399508 373868 399560
rect 374460 399508 374512 399560
rect 373632 399440 373684 399492
rect 374092 399440 374144 399492
rect 374782 399780 374834 399832
rect 374828 399576 374880 399628
rect 374736 399440 374788 399492
rect 374460 399372 374512 399424
rect 375242 399848 375294 399900
rect 375886 399848 375938 399900
rect 376070 399848 376122 399900
rect 376346 399848 376398 399900
rect 376438 399848 376490 399900
rect 376806 399848 376858 399900
rect 377726 399848 377778 399900
rect 377818 399848 377870 399900
rect 378186 399848 378238 399900
rect 378278 399848 378330 399900
rect 378922 399848 378974 399900
rect 375058 399780 375110 399832
rect 375150 399780 375202 399832
rect 375196 399644 375248 399696
rect 375104 399576 375156 399628
rect 375196 399508 375248 399560
rect 375610 399780 375662 399832
rect 374920 399440 374972 399492
rect 375380 399440 375432 399492
rect 375748 399508 375800 399560
rect 376208 399576 376260 399628
rect 377082 399780 377134 399832
rect 377174 399780 377226 399832
rect 377358 399780 377410 399832
rect 377450 399780 377502 399832
rect 376944 399644 376996 399696
rect 377036 399644 377088 399696
rect 376392 399508 376444 399560
rect 376300 399236 376352 399288
rect 377312 399644 377364 399696
rect 377680 399712 377732 399764
rect 377772 399712 377824 399764
rect 377404 399508 377456 399560
rect 378600 399508 378652 399560
rect 378600 399372 378652 399424
rect 387892 400052 387944 400104
rect 379106 399848 379158 399900
rect 379382 399848 379434 399900
rect 379750 399848 379802 399900
rect 380302 399848 380354 399900
rect 380670 399848 380722 399900
rect 381222 399848 381274 399900
rect 381498 399848 381550 399900
rect 381590 399848 381642 399900
rect 381958 399848 382010 399900
rect 382234 399848 382286 399900
rect 382602 399848 382654 399900
rect 382786 399848 382838 399900
rect 383430 399848 383482 399900
rect 383706 399848 383758 399900
rect 383798 399848 383850 399900
rect 384166 399848 384218 399900
rect 384258 399848 384310 399900
rect 384442 399848 384494 399900
rect 379336 399712 379388 399764
rect 379704 399712 379756 399764
rect 379980 399712 380032 399764
rect 379428 399644 379480 399696
rect 379612 399644 379664 399696
rect 379152 399508 379204 399560
rect 379796 399508 379848 399560
rect 380486 399780 380538 399832
rect 380532 399644 380584 399696
rect 380440 399576 380492 399628
rect 380900 399508 380952 399560
rect 381360 399576 381412 399628
rect 381544 399508 381596 399560
rect 381912 399508 381964 399560
rect 382648 399712 382700 399764
rect 383568 399644 383620 399696
rect 383936 399644 383988 399696
rect 384304 399644 384356 399696
rect 385086 399780 385138 399832
rect 384718 399712 384770 399764
rect 382372 399508 382424 399560
rect 383292 399508 383344 399560
rect 380256 399440 380308 399492
rect 384580 399508 384632 399560
rect 384764 399440 384816 399492
rect 387984 399984 388036 400036
rect 390192 399916 390244 399968
rect 385546 399848 385598 399900
rect 385914 399848 385966 399900
rect 386006 399848 386058 399900
rect 386558 399848 386610 399900
rect 387018 399848 387070 399900
rect 387202 399848 387254 399900
rect 387524 399848 387576 399900
rect 385638 399780 385690 399832
rect 385684 399644 385736 399696
rect 385868 399644 385920 399696
rect 385776 399576 385828 399628
rect 386190 399780 386242 399832
rect 386236 399576 386288 399628
rect 386420 399576 386472 399628
rect 386742 399780 386794 399832
rect 387110 399780 387162 399832
rect 386788 399644 386840 399696
rect 386880 399576 386932 399628
rect 389180 399508 389232 399560
rect 385592 399440 385644 399492
rect 387800 399372 387852 399424
rect 378692 399304 378744 399356
rect 379244 399304 379296 399356
rect 377680 399236 377732 399288
rect 379612 399168 379664 399220
rect 338028 399100 338080 399152
rect 366180 399100 366232 399152
rect 334992 399032 335044 399084
rect 278688 398964 278740 399016
rect 348516 398964 348568 399016
rect 349988 398964 350040 399016
rect 362868 399032 362920 399084
rect 364524 399032 364576 399084
rect 379244 399100 379296 399152
rect 381636 399100 381688 399152
rect 381912 399100 381964 399152
rect 340512 398896 340564 398948
rect 355968 398896 356020 398948
rect 356152 398896 356204 398948
rect 356520 398896 356572 398948
rect 366180 398964 366232 399016
rect 365904 398896 365956 398948
rect 375748 398896 375800 398948
rect 381176 398896 381228 398948
rect 382188 398896 382240 398948
rect 382464 398896 382516 398948
rect 340420 398828 340472 398880
rect 349988 398828 350040 398880
rect 354404 398828 354456 398880
rect 355876 398828 355928 398880
rect 339132 398760 339184 398812
rect 348148 398760 348200 398812
rect 348700 398760 348752 398812
rect 352104 398760 352156 398812
rect 354036 398760 354088 398812
rect 355416 398760 355468 398812
rect 356520 398760 356572 398812
rect 374276 398828 374328 398880
rect 375472 398828 375524 398880
rect 383016 398828 383068 398880
rect 383568 398828 383620 398880
rect 385684 398828 385736 398880
rect 394700 398828 394752 398880
rect 363696 398760 363748 398812
rect 364064 398760 364116 398812
rect 365628 398760 365680 398812
rect 343824 398692 343876 398744
rect 344836 398692 344888 398744
rect 330760 398624 330812 398676
rect 346032 398692 346084 398744
rect 347780 398692 347832 398744
rect 348516 398692 348568 398744
rect 356428 398692 356480 398744
rect 359188 398692 359240 398744
rect 359556 398692 359608 398744
rect 376944 398760 376996 398812
rect 379060 398760 379112 398812
rect 381084 398692 381136 398744
rect 365536 398624 365588 398676
rect 382556 398624 382608 398676
rect 388076 398624 388128 398676
rect 305092 398556 305144 398608
rect 340328 398556 340380 398608
rect 303620 398488 303672 398540
rect 342904 398488 342956 398540
rect 295340 398420 295392 398472
rect 343916 398420 343968 398472
rect 349252 398556 349304 398608
rect 351552 398556 351604 398608
rect 371424 398556 371476 398608
rect 382372 398556 382424 398608
rect 389272 398556 389324 398608
rect 345020 398488 345072 398540
rect 345940 398488 345992 398540
rect 346124 398488 346176 398540
rect 345664 398420 345716 398472
rect 354404 398420 354456 398472
rect 355508 398488 355560 398540
rect 357348 398488 357400 398540
rect 359556 398488 359608 398540
rect 363144 398488 363196 398540
rect 380992 398488 381044 398540
rect 390652 398488 390704 398540
rect 360660 398420 360712 398472
rect 382924 398420 382976 398472
rect 389548 398420 389600 398472
rect 289084 398352 289136 398404
rect 344100 398352 344152 398404
rect 344928 398352 344980 398404
rect 348332 398352 348384 398404
rect 362684 398352 362736 398404
rect 373816 398352 373868 398404
rect 384488 398352 384540 398404
rect 386604 398352 386656 398404
rect 392032 398352 392084 398404
rect 260748 398216 260800 398268
rect 341892 398284 341944 398336
rect 304264 398148 304316 398200
rect 305644 398148 305696 398200
rect 345112 398284 345164 398336
rect 342904 398216 342956 398268
rect 346124 398284 346176 398336
rect 348148 398284 348200 398336
rect 352104 398284 352156 398336
rect 354588 398284 354640 398336
rect 360384 398284 360436 398336
rect 371424 398284 371476 398336
rect 372436 398284 372488 398336
rect 363512 398216 363564 398268
rect 365996 398216 366048 398268
rect 378784 398216 378836 398268
rect 390560 398216 390612 398268
rect 257988 398080 258040 398132
rect 341156 398080 341208 398132
rect 354496 398148 354548 398200
rect 372436 398148 372488 398200
rect 376852 398148 376904 398200
rect 386972 398148 387024 398200
rect 353484 398080 353536 398132
rect 358544 398080 358596 398132
rect 341892 398012 341944 398064
rect 357808 398012 357860 398064
rect 376852 398012 376904 398064
rect 377312 398012 377364 398064
rect 377588 398012 377640 398064
rect 378784 398012 378836 398064
rect 386512 398012 386564 398064
rect 386972 398012 387024 398064
rect 387708 398012 387760 398064
rect 342444 397944 342496 397996
rect 343364 397944 343416 397996
rect 346032 397944 346084 397996
rect 352472 397944 352524 397996
rect 352840 397944 352892 397996
rect 333244 397740 333296 397792
rect 344836 397876 344888 397928
rect 351092 397876 351144 397928
rect 352104 397876 352156 397928
rect 354588 397876 354640 397928
rect 341524 397808 341576 397860
rect 343088 397808 343140 397860
rect 349620 397808 349672 397860
rect 350080 397808 350132 397860
rect 348424 397740 348476 397792
rect 352380 397740 352432 397792
rect 274456 397672 274508 397724
rect 277032 397604 277084 397656
rect 333244 397604 333296 397656
rect 345664 397672 345716 397724
rect 345848 397672 345900 397724
rect 349436 397672 349488 397724
rect 350080 397672 350132 397724
rect 367836 397944 367888 397996
rect 374184 397944 374236 397996
rect 382924 397944 382976 397996
rect 381544 397876 381596 397928
rect 381912 397876 381964 397928
rect 372252 397740 372304 397792
rect 374368 397740 374420 397792
rect 381268 397740 381320 397792
rect 381544 397740 381596 397792
rect 356428 397672 356480 397724
rect 356888 397672 356940 397724
rect 361120 397672 361172 397724
rect 361488 397672 361540 397724
rect 338948 397604 339000 397656
rect 355048 397604 355100 397656
rect 330852 397536 330904 397588
rect 353484 397536 353536 397588
rect 355600 397536 355652 397588
rect 357808 397536 357860 397588
rect 360936 397536 360988 397588
rect 363604 397536 363656 397588
rect 340972 397468 341024 397520
rect 346952 397468 347004 397520
rect 349436 397468 349488 397520
rect 349712 397468 349764 397520
rect 351092 397468 351144 397520
rect 351368 397468 351420 397520
rect 356796 397468 356848 397520
rect 357992 397468 358044 397520
rect 358360 397468 358412 397520
rect 362316 397468 362368 397520
rect 376760 397672 376812 397724
rect 386420 397672 386472 397724
rect 387340 397672 387392 397724
rect 385316 397468 385368 397520
rect 389456 397468 389508 397520
rect 334716 397400 334768 397452
rect 359096 397400 359148 397452
rect 372068 397400 372120 397452
rect 386420 397400 386472 397452
rect 387524 397400 387576 397452
rect 345664 397332 345716 397384
rect 362500 397332 362552 397384
rect 364524 397332 364576 397384
rect 364708 397332 364760 397384
rect 365996 397332 366048 397384
rect 366180 397332 366232 397384
rect 382372 397332 382424 397384
rect 382740 397332 382792 397384
rect 385684 397332 385736 397384
rect 385960 397332 386012 397384
rect 332324 397264 332376 397316
rect 359648 397264 359700 397316
rect 330668 397196 330720 397248
rect 358636 397196 358688 397248
rect 383752 397196 383804 397248
rect 389364 397196 389416 397248
rect 337844 397128 337896 397180
rect 380624 397128 380676 397180
rect 380992 397128 381044 397180
rect 382648 397128 382700 397180
rect 384304 397128 384356 397180
rect 384580 397128 384632 397180
rect 336188 397060 336240 397112
rect 383292 397060 383344 397112
rect 306288 396992 306340 397044
rect 366364 396992 366416 397044
rect 386696 396992 386748 397044
rect 387248 396992 387300 397044
rect 276940 396924 276992 396976
rect 339868 396924 339920 396976
rect 349160 396924 349212 396976
rect 349528 396924 349580 396976
rect 377864 396924 377916 396976
rect 381084 396924 381136 396976
rect 280988 396856 281040 396908
rect 350448 396856 350500 396908
rect 355692 396856 355744 396908
rect 360844 396856 360896 396908
rect 362316 396856 362368 396908
rect 371976 396856 372028 396908
rect 378508 396856 378560 396908
rect 381268 396856 381320 396908
rect 390008 396856 390060 396908
rect 394884 396856 394936 396908
rect 271512 396788 271564 396840
rect 353116 396788 353168 396840
rect 354496 396788 354548 396840
rect 354956 396788 355008 396840
rect 377864 396788 377916 396840
rect 379704 396788 379756 396840
rect 340604 396720 340656 396772
rect 345664 396720 345716 396772
rect 355140 396720 355192 396772
rect 360752 396720 360804 396772
rect 367928 396720 367980 396772
rect 368664 396720 368716 396772
rect 377312 396720 377364 396772
rect 381452 396720 381504 396772
rect 346032 396652 346084 396704
rect 351184 396652 351236 396704
rect 358268 396652 358320 396704
rect 358820 396652 358872 396704
rect 363512 396652 363564 396704
rect 363972 396652 364024 396704
rect 377404 396652 377456 396704
rect 377680 396652 377732 396704
rect 383936 396652 383988 396704
rect 384120 396652 384172 396704
rect 385224 396652 385276 396704
rect 385868 396652 385920 396704
rect 257804 396584 257856 396636
rect 343640 396584 343692 396636
rect 363420 396584 363472 396636
rect 363880 396584 363932 396636
rect 336004 396516 336056 396568
rect 352012 396516 352064 396568
rect 382648 396516 382700 396568
rect 383384 396516 383436 396568
rect 355876 396448 355928 396500
rect 361580 396448 361632 396500
rect 383936 396448 383988 396500
rect 384672 396448 384724 396500
rect 360844 396312 360896 396364
rect 362960 396312 363012 396364
rect 351184 396176 351236 396228
rect 355324 396176 355376 396228
rect 372712 396176 372764 396228
rect 373264 396176 373316 396228
rect 341800 396108 341852 396160
rect 354772 396108 354824 396160
rect 385500 396108 385552 396160
rect 386236 396108 386288 396160
rect 346492 396040 346544 396092
rect 346860 396040 346912 396092
rect 335084 395972 335136 396024
rect 361856 396040 361908 396092
rect 360108 395972 360160 396024
rect 363696 395972 363748 396024
rect 379520 395972 379572 396024
rect 379796 395972 379848 396024
rect 341708 395904 341760 395956
rect 368940 395904 368992 395956
rect 381452 395904 381504 395956
rect 382004 395904 382056 395956
rect 340144 395836 340196 395888
rect 368020 395836 368072 395888
rect 336372 395768 336424 395820
rect 369676 395768 369728 395820
rect 330576 395700 330628 395752
rect 365444 395700 365496 395752
rect 281632 395632 281684 395684
rect 303620 395632 303672 395684
rect 329288 395632 329340 395684
rect 368204 395632 368256 395684
rect 369032 395632 369084 395684
rect 369768 395632 369820 395684
rect 372528 395632 372580 395684
rect 374552 395632 374604 395684
rect 383660 395632 383712 395684
rect 384396 395632 384448 395684
rect 281540 395564 281592 395616
rect 305092 395564 305144 395616
rect 339316 395564 339368 395616
rect 381636 395564 381688 395616
rect 385408 395564 385460 395616
rect 386328 395564 386380 395616
rect 278412 395496 278464 395548
rect 347964 395496 348016 395548
rect 350908 395496 350960 395548
rect 351736 395496 351788 395548
rect 356980 395496 357032 395548
rect 361028 395496 361080 395548
rect 366364 395496 366416 395548
rect 370596 395496 370648 395548
rect 275560 395428 275612 395480
rect 353668 395428 353720 395480
rect 378140 395428 378192 395480
rect 379980 395428 380032 395480
rect 346860 395360 346912 395412
rect 347412 395360 347464 395412
rect 354864 395360 354916 395412
rect 356060 395360 356112 395412
rect 361028 395360 361080 395412
rect 374644 395360 374696 395412
rect 275744 395292 275796 395344
rect 341800 395292 341852 395344
rect 337660 395224 337712 395276
rect 352748 395292 352800 395344
rect 355968 395292 356020 395344
rect 343640 395224 343692 395276
rect 350816 395224 350868 395276
rect 353484 395224 353536 395276
rect 354312 395224 354364 395276
rect 367744 395224 367796 395276
rect 368572 395224 368624 395276
rect 369768 395292 369820 395344
rect 371608 395292 371660 395344
rect 371792 395292 371844 395344
rect 372160 395292 372212 395344
rect 374276 395292 374328 395344
rect 375288 395292 375340 395344
rect 369952 395224 370004 395276
rect 374644 395224 374696 395276
rect 375564 395224 375616 395276
rect 375840 395224 375892 395276
rect 376392 395224 376444 395276
rect 328000 395156 328052 395208
rect 343548 395156 343600 395208
rect 374184 395156 374236 395208
rect 375104 395156 375156 395208
rect 267648 395088 267700 395140
rect 345020 395088 345072 395140
rect 364892 395088 364944 395140
rect 365076 395088 365128 395140
rect 370044 395088 370096 395140
rect 371608 395088 371660 395140
rect 378232 395088 378284 395140
rect 390744 395088 390796 395140
rect 361764 395020 361816 395072
rect 362224 395020 362276 395072
rect 345020 394952 345072 395004
rect 350632 394952 350684 395004
rect 353024 394952 353076 395004
rect 354220 394952 354272 395004
rect 361856 394680 361908 394732
rect 362592 394680 362644 394732
rect 341616 394612 341668 394664
rect 360016 394612 360068 394664
rect 334900 394544 334952 394596
rect 359188 394544 359240 394596
rect 336556 394476 336608 394528
rect 368940 394476 368992 394528
rect 339224 394408 339276 394460
rect 378968 394408 379020 394460
rect 322848 394340 322900 394392
rect 382280 394340 382332 394392
rect 272984 394272 273036 394324
rect 345756 394272 345808 394324
rect 276756 394204 276808 394256
rect 339868 394204 339920 394256
rect 279700 394136 279752 394188
rect 358912 394272 358964 394324
rect 359004 394272 359056 394324
rect 359740 394272 359792 394324
rect 352748 394204 352800 394256
rect 374828 394204 374880 394256
rect 375564 394204 375616 394256
rect 376484 394204 376536 394256
rect 380072 394204 380124 394256
rect 380348 394204 380400 394256
rect 354128 394136 354180 394188
rect 264796 394068 264848 394120
rect 342444 394068 342496 394120
rect 385132 394136 385184 394188
rect 385776 394136 385828 394188
rect 272616 394000 272668 394052
rect 342996 394000 343048 394052
rect 347044 394000 347096 394052
rect 352380 394000 352432 394052
rect 352656 394000 352708 394052
rect 376852 394068 376904 394120
rect 386052 394068 386104 394120
rect 389640 394068 389692 394120
rect 355232 394000 355284 394052
rect 356244 394000 356296 394052
rect 357256 394000 357308 394052
rect 273996 393932 274048 393984
rect 342536 393864 342588 393916
rect 343272 393864 343324 393916
rect 342444 393796 342496 393848
rect 344376 393796 344428 393848
rect 357164 393932 357216 393984
rect 359464 393932 359516 393984
rect 376024 393932 376076 393984
rect 376300 393932 376352 393984
rect 350632 393796 350684 393848
rect 351368 393796 351420 393848
rect 352104 393796 352156 393848
rect 352564 393796 352616 393848
rect 376024 393796 376076 393848
rect 376576 393796 376628 393848
rect 377220 393796 377272 393848
rect 377772 393796 377824 393848
rect 364892 393728 364944 393780
rect 374828 393728 374880 393780
rect 377496 393728 377548 393780
rect 378876 393592 378928 393644
rect 379244 393592 379296 393644
rect 345664 393524 345716 393576
rect 347504 393524 347556 393576
rect 348700 393524 348752 393576
rect 349252 393524 349304 393576
rect 363420 393524 363472 393576
rect 364248 393524 364300 393576
rect 345296 393456 345348 393508
rect 346676 393456 346728 393508
rect 351368 393456 351420 393508
rect 353852 393456 353904 393508
rect 363144 393456 363196 393508
rect 364156 393456 364208 393508
rect 364524 393456 364576 393508
rect 364892 393456 364944 393508
rect 367468 393456 367520 393508
rect 368848 393456 368900 393508
rect 339040 393388 339092 393440
rect 346584 393388 346636 393440
rect 347964 393388 348016 393440
rect 349068 393388 349120 393440
rect 349528 393388 349580 393440
rect 349804 393388 349856 393440
rect 360476 393388 360528 393440
rect 361488 393388 361540 393440
rect 362224 393388 362276 393440
rect 370228 393388 370280 393440
rect 321376 393320 321428 393372
rect 378140 393320 378192 393372
rect 282920 393252 282972 393304
rect 344376 393252 344428 393304
rect 346768 393252 346820 393304
rect 347320 393252 347372 393304
rect 348792 393252 348844 393304
rect 349068 393252 349120 393304
rect 349252 393252 349304 393304
rect 350540 393252 350592 393304
rect 350724 393252 350776 393304
rect 351000 393252 351052 393304
rect 353392 393252 353444 393304
rect 354312 393252 354364 393304
rect 359740 393252 359792 393304
rect 360200 393252 360252 393304
rect 364524 393252 364576 393304
rect 364800 393252 364852 393304
rect 365996 393252 366048 393304
rect 366916 393252 366968 393304
rect 367836 393252 367888 393304
rect 370228 393252 370280 393304
rect 341800 393184 341852 393236
rect 386512 393184 386564 393236
rect 341432 393116 341484 393168
rect 366456 393116 366508 393168
rect 373172 393116 373224 393168
rect 373724 393116 373776 393168
rect 336648 393048 336700 393100
rect 364248 393048 364300 393100
rect 364432 393048 364484 393100
rect 364708 393048 364760 393100
rect 364800 393048 364852 393100
rect 365720 393048 365772 393100
rect 315856 392980 315908 393032
rect 375104 392980 375156 393032
rect 282368 392912 282420 392964
rect 342720 392912 342772 392964
rect 343456 392912 343508 392964
rect 345480 392912 345532 392964
rect 346124 392912 346176 392964
rect 350264 392912 350316 392964
rect 358268 392912 358320 392964
rect 358728 392912 358780 392964
rect 359464 392912 359516 392964
rect 364984 392912 365036 392964
rect 279792 392844 279844 392896
rect 345204 392844 345256 392896
rect 349160 392844 349212 392896
rect 349344 392844 349396 392896
rect 363604 392844 363656 392896
rect 366732 392844 366784 392896
rect 276296 392776 276348 392828
rect 350080 392776 350132 392828
rect 370596 392776 370648 392828
rect 370964 392776 371016 392828
rect 347044 392708 347096 392760
rect 348884 392708 348936 392760
rect 352748 392708 352800 392760
rect 381728 392708 381780 392760
rect 274088 392640 274140 392692
rect 353208 392640 353260 392692
rect 271420 392572 271472 392624
rect 363328 392572 363380 392624
rect 371884 392572 371936 392624
rect 382372 392572 382424 392624
rect 330484 392504 330536 392556
rect 343548 392504 343600 392556
rect 359556 392504 359608 392556
rect 360108 392504 360160 392556
rect 271604 392436 271656 392488
rect 361672 392436 361724 392488
rect 344284 392368 344336 392420
rect 353576 392368 353628 392420
rect 375748 392368 375800 392420
rect 376116 392368 376168 392420
rect 365076 392300 365128 392352
rect 369860 392300 369912 392352
rect 367836 392232 367888 392284
rect 368480 392232 368532 392284
rect 355508 392028 355560 392080
rect 364340 392028 364392 392080
rect 364984 391960 365036 392012
rect 370412 391960 370464 392012
rect 360752 391824 360804 391876
rect 361120 391824 361172 391876
rect 367192 391756 367244 391808
rect 369860 391756 369912 391808
rect 311808 391416 311860 391468
rect 371700 391416 371752 391468
rect 281724 391348 281776 391400
rect 342260 391348 342312 391400
rect 270316 391280 270368 391332
rect 344652 391348 344704 391400
rect 343364 391280 343416 391332
rect 381084 391348 381136 391400
rect 368664 391280 368716 391332
rect 369308 391280 369360 391332
rect 369400 391280 369452 391332
rect 371700 391280 371752 391332
rect 267556 391212 267608 391264
rect 348240 391212 348292 391264
rect 359188 391212 359240 391264
rect 359832 391212 359884 391264
rect 363696 391212 363748 391264
rect 383108 391212 383160 391264
rect 374460 391076 374512 391128
rect 374920 391076 374972 391128
rect 341800 391008 341852 391060
rect 354956 391008 355008 391060
rect 313188 390600 313240 390652
rect 372620 390600 372672 390652
rect 314384 390532 314436 390584
rect 374000 390532 374052 390584
rect 345940 390464 345992 390516
rect 375472 390464 375524 390516
rect 356704 390328 356756 390380
rect 360568 390328 360620 390380
rect 337568 390192 337620 390244
rect 345572 390192 345624 390244
rect 319168 390124 319220 390176
rect 379336 390124 379388 390176
rect 319812 390056 319864 390108
rect 378140 390056 378192 390108
rect 319904 389988 319956 390040
rect 380164 389988 380216 390040
rect 281816 389920 281868 389972
rect 342628 389920 342680 389972
rect 343088 389920 343140 389972
rect 367008 389920 367060 389972
rect 269856 389852 269908 389904
rect 342444 389852 342496 389904
rect 259276 389784 259328 389836
rect 347136 389784 347188 389836
rect 351276 389716 351328 389768
rect 361764 389716 361816 389768
rect 347136 389512 347188 389564
rect 354496 389512 354548 389564
rect 349804 389308 349856 389360
rect 355140 389308 355192 389360
rect 318708 389172 318760 389224
rect 378140 389172 378192 389224
rect 351000 388968 351052 389020
rect 351460 388968 351512 389020
rect 333520 388696 333572 388748
rect 365168 388696 365220 388748
rect 343548 388628 343600 388680
rect 383660 388628 383712 388680
rect 276664 388560 276716 388612
rect 343180 388560 343232 388612
rect 262128 388492 262180 388544
rect 348056 388492 348108 388544
rect 349896 388492 349948 388544
rect 381452 388492 381504 388544
rect 257896 388424 257948 388476
rect 347596 388424 347648 388476
rect 354220 388424 354272 388476
rect 386420 388424 386472 388476
rect 356704 388016 356756 388068
rect 356980 388016 357032 388068
rect 352564 387880 352616 387932
rect 354864 387880 354916 387932
rect 321744 387744 321796 387796
rect 322480 387744 322532 387796
rect 348516 387744 348568 387796
rect 355692 387744 355744 387796
rect 348608 387608 348660 387660
rect 357164 387608 357216 387660
rect 331036 387540 331088 387592
rect 355232 387540 355284 387592
rect 305092 387472 305144 387524
rect 305644 387472 305696 387524
rect 329380 387472 329432 387524
rect 365352 387472 365404 387524
rect 333612 387404 333664 387456
rect 373448 387404 373500 387456
rect 332416 387336 332468 387388
rect 374828 387336 374880 387388
rect 329472 387268 329524 387320
rect 371976 387268 372028 387320
rect 275468 387200 275520 387252
rect 341248 387200 341300 387252
rect 347320 387200 347372 387252
rect 359372 387200 359424 387252
rect 263416 387132 263468 387184
rect 342812 387132 342864 387184
rect 344560 387132 344612 387184
rect 357716 387132 357768 387184
rect 275376 387064 275428 387116
rect 363512 387064 363564 387116
rect 262864 386452 262916 386504
rect 321744 386452 321796 386504
rect 279148 386384 279200 386436
rect 292580 386384 292632 386436
rect 293868 386384 293920 386436
rect 580264 386384 580316 386436
rect 320456 386316 320508 386368
rect 320916 386316 320968 386368
rect 277860 385976 277912 386028
rect 349988 385976 350040 386028
rect 280712 385908 280764 385960
rect 358360 385908 358412 385960
rect 279516 385840 279568 385892
rect 360752 385840 360804 385892
rect 268936 385772 268988 385824
rect 353024 385772 353076 385824
rect 279608 385704 279660 385756
rect 368112 385704 368164 385756
rect 3424 385636 3476 385688
rect 255320 385636 255372 385688
rect 278228 385636 278280 385688
rect 366364 385636 366416 385688
rect 269948 385160 270000 385212
rect 320456 385160 320508 385212
rect 264520 385092 264572 385144
rect 323768 385092 323820 385144
rect 255320 385024 255372 385076
rect 316224 385024 316276 385076
rect 316684 385024 316736 385076
rect 319076 384956 319128 385008
rect 319720 384956 319772 385008
rect 325700 384956 325752 385008
rect 326344 384956 326396 385008
rect 344468 384956 344520 385008
rect 358268 384956 358320 385008
rect 345940 384888 345992 384940
rect 361212 384888 361264 384940
rect 348700 384820 348752 384872
rect 363236 384820 363288 384872
rect 346216 384752 346268 384804
rect 361856 384752 361908 384804
rect 344836 384684 344888 384736
rect 362408 384684 362460 384736
rect 343180 384616 343232 384668
rect 363144 384616 363196 384668
rect 345848 384548 345900 384600
rect 366088 384548 366140 384600
rect 347412 384480 347464 384532
rect 370688 384480 370740 384532
rect 338672 384412 338724 384464
rect 364708 384412 364760 384464
rect 329196 384344 329248 384396
rect 379980 384344 380032 384396
rect 283564 384276 283616 384328
rect 352840 384276 352892 384328
rect 262956 383800 263008 383852
rect 322296 383800 322348 383852
rect 265900 383732 265952 383784
rect 325700 383732 325752 383784
rect 257344 383664 257396 383716
rect 319076 383664 319128 383716
rect 313924 383596 313976 383648
rect 314200 383596 314252 383648
rect 314844 383052 314896 383104
rect 315488 383052 315540 383104
rect 318892 382984 318944 383036
rect 319628 382984 319680 383036
rect 318984 382576 319036 382628
rect 319536 382576 319588 382628
rect 272524 382508 272576 382560
rect 321652 382508 321704 382560
rect 322388 382508 322440 382560
rect 265716 382440 265768 382492
rect 318892 382440 318944 382492
rect 253204 382372 253256 382424
rect 313464 382372 313516 382424
rect 258724 382304 258776 382356
rect 318984 382304 319036 382356
rect 254584 382236 254636 382288
rect 314844 382236 314896 382288
rect 324412 381964 324464 382016
rect 324964 381964 325016 382016
rect 343272 381624 343324 381676
rect 359004 381624 359056 381676
rect 345756 381556 345808 381608
rect 368756 381556 368808 381608
rect 350172 381488 350224 381540
rect 374276 381488 374328 381540
rect 279424 381148 279476 381200
rect 317512 381148 317564 381200
rect 318248 381148 318300 381200
rect 261484 381080 261536 381132
rect 311256 381080 311308 381132
rect 268384 381012 268436 381064
rect 246304 380944 246356 380996
rect 305092 380944 305144 380996
rect 264336 380876 264388 380928
rect 324412 380876 324464 380928
rect 324596 380876 324648 380928
rect 325056 380876 325108 380928
rect 250536 379856 250588 379908
rect 309140 379856 309192 379908
rect 309324 379856 309376 379908
rect 254768 379788 254820 379840
rect 314752 379788 314804 379840
rect 246396 379720 246448 379772
rect 306380 379720 306432 379772
rect 306564 379720 306616 379772
rect 255964 379652 256016 379704
rect 316132 379652 316184 379704
rect 243544 379584 243596 379636
rect 303620 379584 303672 379636
rect 259828 379516 259880 379568
rect 320364 379516 320416 379568
rect 321008 379516 321060 379568
rect 317604 378972 317656 379024
rect 318156 378972 318208 379024
rect 286784 378836 286836 378888
rect 341984 378972 342036 379024
rect 307668 378768 307720 378820
rect 345296 378836 345348 378888
rect 342076 378700 342128 378752
rect 367376 378768 367428 378820
rect 317512 378360 317564 378412
rect 317972 378360 318024 378412
rect 259184 378292 259236 378344
rect 317604 378292 317656 378344
rect 253848 378224 253900 378276
rect 314108 378224 314160 378276
rect 262220 378156 262272 378208
rect 322940 378156 322992 378208
rect 323676 378156 323728 378208
rect 301964 377408 302016 377460
rect 337292 377408 337344 377460
rect 351460 377408 351512 377460
rect 359280 377408 359332 377460
rect 250444 376864 250496 376916
rect 302608 376864 302660 376916
rect 302884 376864 302936 376916
rect 263048 376796 263100 376848
rect 323584 376796 323636 376848
rect 323860 376796 323912 376848
rect 254676 376728 254728 376780
rect 315396 376728 315448 376780
rect 261576 376048 261628 376100
rect 300308 376048 300360 376100
rect 267188 375980 267240 376032
rect 310888 375980 310940 376032
rect 267096 375912 267148 375964
rect 312176 375912 312228 375964
rect 264244 375844 264296 375896
rect 312820 375844 312872 375896
rect 232504 375776 232556 375828
rect 291844 375776 291896 375828
rect 292304 375776 292356 375828
rect 235264 375708 235316 375760
rect 294420 375708 294472 375760
rect 294696 375708 294748 375760
rect 237380 375640 237432 375692
rect 297456 375640 297508 375692
rect 240140 375572 240192 375624
rect 300400 375572 300452 375624
rect 261668 375504 261720 375556
rect 321836 375504 321888 375556
rect 322204 375504 322256 375556
rect 236644 375436 236696 375488
rect 297548 375436 297600 375488
rect 220728 375368 220780 375420
rect 291752 375368 291804 375420
rect 291936 375368 291988 375420
rect 297456 375368 297508 375420
rect 297732 375368 297784 375420
rect 281172 375300 281224 375352
rect 281448 375300 281500 375352
rect 258816 374960 258868 375012
rect 298376 374960 298428 375012
rect 259552 374892 259604 374944
rect 319536 374892 319588 374944
rect 281172 374756 281224 374808
rect 307300 374756 307352 374808
rect 275652 374688 275704 374740
rect 300860 374688 300912 374740
rect 301596 374688 301648 374740
rect 220084 374620 220136 374672
rect 282000 374620 282052 374672
rect 314752 374620 314804 374672
rect 315396 374620 315448 374672
rect 321652 374620 321704 374672
rect 322388 374620 322440 374672
rect 324412 374620 324464 374672
rect 324964 374620 325016 374672
rect 273168 374552 273220 374604
rect 301964 374552 302016 374604
rect 264612 374484 264664 374536
rect 294788 374484 294840 374536
rect 305552 374484 305604 374536
rect 305736 374484 305788 374536
rect 272800 374416 272852 374468
rect 304356 374416 304408 374468
rect 264428 374348 264480 374400
rect 297088 374348 297140 374400
rect 274548 374280 274600 374332
rect 308404 374280 308456 374332
rect 272708 374212 272760 374264
rect 307024 374212 307076 374264
rect 267280 374144 267332 374196
rect 305552 374144 305604 374196
rect 290188 374076 290240 374128
rect 295524 374076 295576 374128
rect 300124 374076 300176 374128
rect 277308 374008 277360 374060
rect 278504 374008 278556 374060
rect 283564 374008 283616 374060
rect 153200 373940 153252 373992
rect 282276 373940 282328 373992
rect 304816 373940 304868 373992
rect 309784 373940 309836 373992
rect 277952 373464 278004 373516
rect 281448 373464 281500 373516
rect 294328 373464 294380 373516
rect 294788 373464 294840 373516
rect 278780 373396 278832 373448
rect 278320 373328 278372 373380
rect 287428 373328 287480 373380
rect 226984 373260 227036 373312
rect 278596 373260 278648 373312
rect 288532 373260 288584 373312
rect 298468 373396 298520 373448
rect 337936 373396 337988 373448
rect 295616 373328 295668 373380
rect 297548 373328 297600 373380
rect 340696 373328 340748 373380
rect 296628 373260 296680 373312
rect 340052 373260 340104 373312
rect 220360 373192 220412 373244
rect 282184 373192 282236 373244
rect 286508 373192 286560 373244
rect 278596 373124 278648 373176
rect 278780 373124 278832 373176
rect 278136 373056 278188 373108
rect 295524 373124 295576 373176
rect 281448 373056 281500 373108
rect 298468 373056 298520 373108
rect 275836 372988 275888 373040
rect 295616 372988 295668 373040
rect 275192 372920 275244 372972
rect 300216 372920 300268 372972
rect 267464 372852 267516 372904
rect 301320 372852 301372 372904
rect 244924 372784 244976 372836
rect 304816 372784 304868 372836
rect 238116 372716 238168 372768
rect 299204 372716 299256 372768
rect 273076 372648 273128 372700
rect 303436 372648 303488 372700
rect 306932 372648 306984 372700
rect 308496 372648 308548 372700
rect 219900 372580 219952 372632
rect 293224 372580 293276 372632
rect 342076 372580 342128 372632
rect 3240 372512 3292 372564
rect 259184 372512 259236 372564
rect 303436 372512 303488 372564
rect 337384 372512 337436 372564
rect 309508 372444 309560 372496
rect 309968 372444 310020 372496
rect 315212 372444 315264 372496
rect 315764 372444 315816 372496
rect 323768 372444 323820 372496
rect 324320 372444 324372 372496
rect 279240 372376 279292 372428
rect 320824 372376 320876 372428
rect 321468 372376 321520 372428
rect 291752 372308 291804 372360
rect 327724 372308 327776 372360
rect 239404 372240 239456 372292
rect 295248 372240 295300 372292
rect 316040 372240 316092 372292
rect 316868 372240 316920 372292
rect 238024 372172 238076 372224
rect 293040 372172 293092 372224
rect 293868 372104 293920 372156
rect 329656 372104 329708 372156
rect 288256 372036 288308 372088
rect 328368 372036 328420 372088
rect 332692 372036 332744 372088
rect 333428 372036 333480 372088
rect 282000 371968 282052 372020
rect 306932 371968 306984 372020
rect 331220 371968 331272 372020
rect 347504 371968 347556 372020
rect 280620 371900 280672 371952
rect 285220 371900 285272 371952
rect 304724 371900 304776 371952
rect 332232 371900 332284 371952
rect 332600 371900 332652 371952
rect 345572 371900 345624 371952
rect 275284 371832 275336 371884
rect 290464 371832 290516 371884
rect 295248 371832 295300 371884
rect 336464 371832 336516 371884
rect 282276 371764 282328 371816
rect 282460 371764 282512 371816
rect 308312 371764 308364 371816
rect 280620 371696 280672 371748
rect 302884 371696 302936 371748
rect 280528 371628 280580 371680
rect 315764 371628 315816 371680
rect 280896 371560 280948 371612
rect 316040 371560 316092 371612
rect 273812 371492 273864 371544
rect 309508 371492 309560 371544
rect 276572 371424 276624 371476
rect 302884 371424 302936 371476
rect 314016 371424 314068 371476
rect 293868 371356 293920 371408
rect 303528 371356 303580 371408
rect 303988 371356 304040 371408
rect 320272 371356 320324 371408
rect 332692 371356 332744 371408
rect 325424 371288 325476 371340
rect 332600 371288 332652 371340
rect 332968 371288 333020 371340
rect 259184 371220 259236 371272
rect 259736 371220 259788 371272
rect 287796 371220 287848 371272
rect 290740 371220 290792 371272
rect 281356 371152 281408 371204
rect 291844 371220 291896 371272
rect 323584 371220 323636 371272
rect 331220 371220 331272 371272
rect 331680 371220 331732 371272
rect 299204 371152 299256 371204
rect 332048 371152 332100 371204
rect 318892 371084 318944 371136
rect 319168 371084 319220 371136
rect 279884 370948 279936 371000
rect 307760 370948 307812 371000
rect 301412 370880 301464 370932
rect 333336 370880 333388 370932
rect 234620 370812 234672 370864
rect 233148 370676 233200 370728
rect 281356 370676 281408 370728
rect 231768 370608 231820 370660
rect 280068 370608 280120 370660
rect 303436 370812 303488 370864
rect 335176 370812 335228 370864
rect 296352 370744 296404 370796
rect 332140 370744 332192 370796
rect 298836 370676 298888 370728
rect 335268 370676 335320 370728
rect 295984 370608 296036 370660
rect 334624 370608 334676 370660
rect 339408 370608 339460 370660
rect 523684 370608 523736 370660
rect 258908 370540 258960 370592
rect 318064 370540 318116 370592
rect 318708 370540 318760 370592
rect 342076 370540 342128 370592
rect 580724 370540 580776 370592
rect 228364 370472 228416 370524
rect 278320 370472 278372 370524
rect 290464 370472 290516 370524
rect 294604 370472 294656 370524
rect 580356 370472 580408 370524
rect 271328 370404 271380 370456
rect 301412 370404 301464 370456
rect 282276 370336 282328 370388
rect 312084 370336 312136 370388
rect 265992 370268 266044 370320
rect 298836 370268 298888 370320
rect 281448 370200 281500 370252
rect 314200 370200 314252 370252
rect 235356 370132 235408 370184
rect 296352 370132 296404 370184
rect 242164 370064 242216 370116
rect 302378 370064 302430 370116
rect 303436 370064 303488 370116
rect 306426 370064 306478 370116
rect 307024 370064 307076 370116
rect 312084 370064 312136 370116
rect 312682 370064 312734 370116
rect 314200 370064 314252 370116
rect 314522 370064 314574 370116
rect 318984 370064 319036 370116
rect 320042 370064 320094 370116
rect 322296 370064 322348 370116
rect 323354 370064 323406 370116
rect 280804 369996 280856 370048
rect 317696 369996 317748 370048
rect 279332 369928 279384 369980
rect 279884 369928 279936 369980
rect 293040 369928 293092 369980
rect 339408 369928 339460 369980
rect 245016 369860 245068 369912
rect 304356 369860 304408 369912
rect 340880 369792 340932 369844
rect 291568 369724 291620 369776
rect 233884 369180 233936 369232
rect 279148 369180 279200 369232
rect 231124 369112 231176 369164
rect 291108 369384 291160 369436
rect 292304 369384 292356 369436
rect 245660 368636 245712 368688
rect 305092 369452 305144 369504
rect 305460 369452 305512 369504
rect 243268 368568 243320 368620
rect 303988 369384 304040 369436
rect 228456 368500 228508 368552
rect 276020 368500 276072 368552
rect 340880 369112 340932 369164
rect 341984 369112 342036 369164
rect 580632 369112 580684 369164
rect 333888 368976 333940 369028
rect 334624 368976 334676 369028
rect 388444 368500 388496 368552
rect 329748 367752 329800 367804
rect 384304 367752 384356 367804
rect 329656 365644 329708 365696
rect 342168 365644 342220 365696
rect 580172 365644 580224 365696
rect 249064 363604 249116 363656
rect 274548 363604 274600 363656
rect 329104 363604 329156 363656
rect 382648 363604 382700 363656
rect 256056 362176 256108 362228
rect 280528 362176 280580 362228
rect 224224 361564 224276 361616
rect 279884 361564 279936 361616
rect 280068 361564 280120 361616
rect 253296 359456 253348 359508
rect 280620 359456 280672 359508
rect 331128 359456 331180 359508
rect 375840 359456 375892 359508
rect 268568 358028 268620 358080
rect 279424 358028 279476 358080
rect 333336 358028 333388 358080
rect 352196 358028 352248 358080
rect 3148 357416 3200 357468
rect 268568 357416 268620 357468
rect 335176 356668 335228 356720
rect 345388 356668 345440 356720
rect 333428 355308 333480 355360
rect 350632 355308 350684 355360
rect 229836 353948 229888 354000
rect 276020 353948 276072 354000
rect 330392 353948 330444 354000
rect 375748 353948 375800 354000
rect 276020 353268 276072 353320
rect 277308 353268 277360 353320
rect 278044 353268 278096 353320
rect 257436 351160 257488 351212
rect 280896 351160 280948 351212
rect 261760 349800 261812 349852
rect 279240 349800 279292 349852
rect 332048 349800 332100 349852
rect 351644 349800 351696 349852
rect 332140 348372 332192 348424
rect 349252 348372 349304 348424
rect 256700 345652 256752 345704
rect 280804 345652 280856 345704
rect 3332 345040 3384 345092
rect 256700 345040 256752 345092
rect 332232 342864 332284 342916
rect 349620 342864 349672 342916
rect 329564 334568 329616 334620
rect 385684 334568 385736 334620
rect 380164 333956 380216 334008
rect 380808 333956 380860 334008
rect 498200 333956 498252 334008
rect 333704 333208 333756 333260
rect 389640 333208 389692 333260
rect 379888 332596 379940 332648
rect 484400 332596 484452 332648
rect 335912 331848 335964 331900
rect 379888 331848 379940 331900
rect 385316 330488 385368 330540
rect 385776 330488 385828 330540
rect 386972 329808 387024 329860
rect 569960 329808 570012 329860
rect 329012 329060 329064 329112
rect 384212 329060 384264 329112
rect 385316 327020 385368 327072
rect 385592 327020 385644 327072
rect 280988 326544 281040 326596
rect 337292 326408 337344 326460
rect 378600 326408 378652 326460
rect 233976 326340 234028 326392
rect 276572 326340 276624 326392
rect 280988 326340 281040 326392
rect 329656 326340 329708 326392
rect 372988 326340 373040 326392
rect 385316 325728 385368 325780
rect 547880 325728 547932 325780
rect 385684 325660 385736 325712
rect 563060 325660 563112 325712
rect 388444 325592 388496 325644
rect 579988 325592 580040 325644
rect 333980 325048 334032 325100
rect 378508 325048 378560 325100
rect 337200 324980 337252 325032
rect 377220 324980 377272 325032
rect 231216 324912 231268 324964
rect 275284 324912 275336 324964
rect 372620 324912 372672 324964
rect 384488 324912 384540 324964
rect 396080 324912 396132 324964
rect 340788 323688 340840 323740
rect 372620 323688 372672 323740
rect 342260 323620 342312 323672
rect 385408 323620 385460 323672
rect 331220 323552 331272 323604
rect 331772 323552 331824 323604
rect 384120 323552 384172 323604
rect 263324 322940 263376 322992
rect 280988 322940 281040 322992
rect 330392 322872 330444 322924
rect 384028 322872 384080 322924
rect 331312 322804 331364 322856
rect 338028 322804 338080 322856
rect 209688 322260 209740 322312
rect 260472 322260 260524 322312
rect 212448 322192 212500 322244
rect 263324 322192 263376 322244
rect 332692 322192 332744 322244
rect 385776 322260 385828 322312
rect 327448 321852 327500 321904
rect 327632 321852 327684 321904
rect 216588 321648 216640 321700
rect 265808 321648 265860 321700
rect 204076 321580 204128 321632
rect 273904 321580 273956 321632
rect 378048 321580 378100 321632
rect 378416 321580 378468 321632
rect 327816 321512 327868 321564
rect 328092 321512 328144 321564
rect 275284 321376 275336 321428
rect 279516 321376 279568 321428
rect 282000 321376 282052 321428
rect 249156 321104 249208 321156
rect 273812 321104 273864 321156
rect 208308 320900 208360 320952
rect 268660 321036 268712 321088
rect 277860 320968 277912 321020
rect 209504 320832 209556 320884
rect 280896 320832 280948 320884
rect 282092 320696 282144 320748
rect 285910 320696 285962 320748
rect 290234 320696 290286 320748
rect 274364 320628 274416 320680
rect 280620 320628 280672 320680
rect 273536 320356 273588 320408
rect 280712 320492 280764 320544
rect 281356 320492 281408 320544
rect 271052 320288 271104 320340
rect 282184 320288 282236 320340
rect 216404 320152 216456 320204
rect 272432 320084 272484 320136
rect 272616 320084 272668 320136
rect 282184 320084 282236 320136
rect 282000 320016 282052 320068
rect 281908 319948 281960 320000
rect 273996 319880 274048 319932
rect 216496 319812 216548 319864
rect 276940 319812 276992 319864
rect 282598 319812 282650 319864
rect 284852 319880 284904 319932
rect 286094 319880 286146 319932
rect 289958 319880 290010 319932
rect 290142 319880 290194 319932
rect 290280 319880 290332 319932
rect 289268 319812 289320 319864
rect 213092 319744 213144 319796
rect 269488 319744 269540 319796
rect 217968 319608 218020 319660
rect 281724 319744 281776 319796
rect 282828 319744 282880 319796
rect 284852 319744 284904 319796
rect 280896 319676 280948 319728
rect 290878 319880 290930 319932
rect 290188 319744 290240 319796
rect 279976 319608 280028 319660
rect 280528 319608 280580 319660
rect 216312 319540 216364 319592
rect 277124 319540 277176 319592
rect 213736 319472 213788 319524
rect 274180 319472 274232 319524
rect 282828 319472 282880 319524
rect 3424 319404 3476 319456
rect 258356 319404 258408 319456
rect 258908 319404 258960 319456
rect 276940 319404 276992 319456
rect 282000 319404 282052 319456
rect 283288 319336 283340 319388
rect 283564 319472 283616 319524
rect 286600 319540 286652 319592
rect 287612 319540 287664 319592
rect 289084 319540 289136 319592
rect 290694 319812 290746 319864
rect 290786 319812 290838 319864
rect 327908 321376 327960 321428
rect 328276 321376 328328 321428
rect 332692 321240 332744 321292
rect 370596 321240 370648 321292
rect 327724 321172 327776 321224
rect 361028 321172 361080 321224
rect 344744 321104 344796 321156
rect 291154 319880 291206 319932
rect 292166 319880 292218 319932
rect 290556 319540 290608 319592
rect 287612 319404 287664 319456
rect 283564 319336 283616 319388
rect 283748 319336 283800 319388
rect 290004 319472 290056 319524
rect 291844 319744 291896 319796
rect 294144 319744 294196 319796
rect 291200 319608 291252 319660
rect 295432 319676 295484 319728
rect 295662 319676 295714 319728
rect 296352 319676 296404 319728
rect 293960 319608 294012 319660
rect 295800 319608 295852 319660
rect 357992 321036 358044 321088
rect 358176 320968 358228 321020
rect 368020 320900 368072 320952
rect 307622 320560 307674 320612
rect 354312 320832 354364 320884
rect 314798 320696 314850 320748
rect 327724 320696 327776 320748
rect 298744 319812 298796 319864
rect 299894 319880 299946 319932
rect 301182 319880 301234 319932
rect 301642 319880 301694 319932
rect 302194 319880 302246 319932
rect 299020 319744 299072 319796
rect 298744 319676 298796 319728
rect 298836 319676 298888 319728
rect 302148 319676 302200 319728
rect 302654 319880 302706 319932
rect 302792 319880 302844 319932
rect 327816 320220 327868 320272
rect 303206 319880 303258 319932
rect 303298 319880 303350 319932
rect 303482 319880 303534 319932
rect 298652 319608 298704 319660
rect 301136 319608 301188 319660
rect 301320 319608 301372 319660
rect 302700 319608 302752 319660
rect 291568 319540 291620 319592
rect 291936 319540 291988 319592
rect 292580 319540 292632 319592
rect 294972 319540 295024 319592
rect 295708 319540 295760 319592
rect 291384 319472 291436 319524
rect 294236 319472 294288 319524
rect 295616 319472 295668 319524
rect 296444 319472 296496 319524
rect 297272 319540 297324 319592
rect 297456 319540 297508 319592
rect 299480 319540 299532 319592
rect 299664 319540 299716 319592
rect 303068 319540 303120 319592
rect 304126 319880 304178 319932
rect 304310 319812 304362 319864
rect 304080 319744 304132 319796
rect 303436 319676 303488 319728
rect 303896 319676 303948 319728
rect 304678 319880 304730 319932
rect 305690 319880 305742 319932
rect 306518 319880 306570 319932
rect 306794 319880 306846 319932
rect 307024 319880 307076 319932
rect 304632 319744 304684 319796
rect 307484 319676 307536 319728
rect 327724 320084 327776 320136
rect 327540 320016 327592 320068
rect 328368 320152 328420 320204
rect 332692 320152 332744 320204
rect 308910 319880 308962 319932
rect 309278 319880 309330 319932
rect 306104 319608 306156 319660
rect 307944 319608 307996 319660
rect 310106 319880 310158 319932
rect 310750 319880 310802 319932
rect 312314 319880 312366 319932
rect 309508 319812 309560 319864
rect 310658 319812 310710 319864
rect 311946 319812 311998 319864
rect 310796 319744 310848 319796
rect 308864 319676 308916 319728
rect 309416 319676 309468 319728
rect 310704 319676 310756 319728
rect 307116 319540 307168 319592
rect 307300 319540 307352 319592
rect 307668 319540 307720 319592
rect 307852 319540 307904 319592
rect 308680 319540 308732 319592
rect 308956 319540 309008 319592
rect 310888 319608 310940 319660
rect 311348 319608 311400 319660
rect 311900 319608 311952 319660
rect 313050 319880 313102 319932
rect 314246 319880 314298 319932
rect 314522 319880 314574 319932
rect 315258 319880 315310 319932
rect 313556 319676 313608 319728
rect 313832 319676 313884 319728
rect 314614 319812 314666 319864
rect 312452 319608 312504 319660
rect 312912 319608 312964 319660
rect 314384 319608 314436 319660
rect 316086 319880 316138 319932
rect 317374 319880 317426 319932
rect 317558 319880 317610 319932
rect 315672 319608 315724 319660
rect 316868 319608 316920 319660
rect 317236 319608 317288 319660
rect 318662 319880 318714 319932
rect 319214 319880 319266 319932
rect 319398 319880 319450 319932
rect 320318 319880 320370 319932
rect 320548 319880 320600 319932
rect 321146 319880 321198 319932
rect 318846 319812 318898 319864
rect 319950 319812 320002 319864
rect 320548 319744 320600 319796
rect 320364 319676 320416 319728
rect 324044 319880 324096 319932
rect 325102 319880 325154 319932
rect 325654 319880 325706 319932
rect 327126 319880 327178 319932
rect 322158 319812 322210 319864
rect 322204 319676 322256 319728
rect 323032 319676 323084 319728
rect 323216 319676 323268 319728
rect 323952 319676 324004 319728
rect 324550 319812 324602 319864
rect 324320 319744 324372 319796
rect 325746 319812 325798 319864
rect 327632 319812 327684 319864
rect 346584 319744 346636 319796
rect 325148 319676 325200 319728
rect 317696 319608 317748 319660
rect 318708 319608 318760 319660
rect 318800 319608 318852 319660
rect 319260 319608 319312 319660
rect 319352 319608 319404 319660
rect 319904 319608 319956 319660
rect 321284 319608 321336 319660
rect 322848 319608 322900 319660
rect 328368 319676 328420 319728
rect 326528 319608 326580 319660
rect 326712 319608 326764 319660
rect 327816 319608 327868 319660
rect 359188 319608 359240 319660
rect 330760 319540 330812 319592
rect 304540 319472 304592 319524
rect 304724 319472 304776 319524
rect 306472 319472 306524 319524
rect 330852 319472 330904 319524
rect 288256 319404 288308 319456
rect 288532 319404 288584 319456
rect 289268 319404 289320 319456
rect 294972 319404 295024 319456
rect 295432 319404 295484 319456
rect 343640 319404 343692 319456
rect 291200 319336 291252 319388
rect 291568 319336 291620 319388
rect 292304 319336 292356 319388
rect 293684 319336 293736 319388
rect 352472 319336 352524 319388
rect 278504 319268 278556 319320
rect 292120 319268 292172 319320
rect 295248 319268 295300 319320
rect 295800 319268 295852 319320
rect 354404 319268 354456 319320
rect 269764 319200 269816 319252
rect 271512 319200 271564 319252
rect 292948 319200 293000 319252
rect 294328 319200 294380 319252
rect 353392 319200 353444 319252
rect 282920 319132 282972 319184
rect 284208 319132 284260 319184
rect 284760 319132 284812 319184
rect 344100 319132 344152 319184
rect 272432 318996 272484 319048
rect 295892 319064 295944 319116
rect 295984 319064 296036 319116
rect 352104 319064 352156 319116
rect 275468 318996 275520 319048
rect 282920 318996 282972 319048
rect 283748 318996 283800 319048
rect 299572 318996 299624 319048
rect 300216 318996 300268 319048
rect 308956 318996 309008 319048
rect 309692 318996 309744 319048
rect 359740 318996 359792 319048
rect 208216 318860 208268 318912
rect 287060 318928 287112 318980
rect 288348 318928 288400 318980
rect 288532 318928 288584 318980
rect 289452 318928 289504 318980
rect 348792 318928 348844 318980
rect 274272 318860 274324 318912
rect 280528 318860 280580 318912
rect 280896 318860 280948 318912
rect 294328 318860 294380 318912
rect 294972 318860 295024 318912
rect 301688 318860 301740 318912
rect 276664 318792 276716 318844
rect 278504 318792 278556 318844
rect 280712 318792 280764 318844
rect 283748 318792 283800 318844
rect 283840 318792 283892 318844
rect 289452 318792 289504 318844
rect 290188 318792 290240 318844
rect 295432 318792 295484 318844
rect 296444 318792 296496 318844
rect 296628 318792 296680 318844
rect 298928 318792 298980 318844
rect 299112 318792 299164 318844
rect 299664 318792 299716 318844
rect 306472 318860 306524 318912
rect 307852 318860 307904 318912
rect 308496 318860 308548 318912
rect 308956 318860 309008 318912
rect 361488 318860 361540 318912
rect 310888 318792 310940 318844
rect 311256 318792 311308 318844
rect 320180 318792 320232 318844
rect 320548 318792 320600 318844
rect 324228 318792 324280 318844
rect 330944 318792 330996 318844
rect 253756 318724 253808 318776
rect 256608 318724 256660 318776
rect 283380 318724 283432 318776
rect 284852 318724 284904 318776
rect 280988 318656 281040 318708
rect 285772 318656 285824 318708
rect 272616 318588 272668 318640
rect 272984 318588 273036 318640
rect 285864 318588 285916 318640
rect 287060 318724 287112 318776
rect 287244 318724 287296 318776
rect 287704 318724 287756 318776
rect 287888 318724 287940 318776
rect 290372 318724 290424 318776
rect 287612 318656 287664 318708
rect 291844 318656 291896 318708
rect 292580 318724 292632 318776
rect 295984 318724 296036 318776
rect 296996 318724 297048 318776
rect 302332 318724 302384 318776
rect 306656 318724 306708 318776
rect 310704 318724 310756 318776
rect 310980 318724 311032 318776
rect 297272 318656 297324 318708
rect 298008 318656 298060 318708
rect 298928 318656 298980 318708
rect 304448 318656 304500 318708
rect 307668 318656 307720 318708
rect 316132 318724 316184 318776
rect 322848 318656 322900 318708
rect 291384 318588 291436 318640
rect 292212 318588 292264 318640
rect 269028 318520 269080 318572
rect 280804 318520 280856 318572
rect 286600 318520 286652 318572
rect 287704 318520 287756 318572
rect 296260 318520 296312 318572
rect 299664 318520 299716 318572
rect 300216 318520 300268 318572
rect 311164 318588 311216 318640
rect 324228 318656 324280 318708
rect 323216 318588 323268 318640
rect 324412 318588 324464 318640
rect 324596 318724 324648 318776
rect 329012 318724 329064 318776
rect 329840 318724 329892 318776
rect 330208 318724 330260 318776
rect 331220 318724 331272 318776
rect 324688 318656 324740 318708
rect 329748 318656 329800 318708
rect 331496 318656 331548 318708
rect 329840 318588 329892 318640
rect 330024 318588 330076 318640
rect 331128 318588 331180 318640
rect 333060 318588 333112 318640
rect 333336 318520 333388 318572
rect 277216 318452 277268 318504
rect 296536 318452 296588 318504
rect 298008 318452 298060 318504
rect 305644 318452 305696 318504
rect 309140 318452 309192 318504
rect 317512 318452 317564 318504
rect 320548 318452 320600 318504
rect 320732 318452 320784 318504
rect 323860 318452 323912 318504
rect 324044 318452 324096 318504
rect 288440 318384 288492 318436
rect 290740 318384 290792 318436
rect 291016 318384 291068 318436
rect 292488 318384 292540 318436
rect 332048 318384 332100 318436
rect 256792 318316 256844 318368
rect 257804 318316 257856 318368
rect 283656 318316 283708 318368
rect 284208 318316 284260 318368
rect 290464 318316 290516 318368
rect 290924 318316 290976 318368
rect 327908 318316 327960 318368
rect 328736 318316 328788 318368
rect 365996 318316 366048 318368
rect 244280 318248 244332 318300
rect 281540 318248 281592 318300
rect 282736 318248 282788 318300
rect 283196 318248 283248 318300
rect 284024 318248 284076 318300
rect 285864 318248 285916 318300
rect 286692 318248 286744 318300
rect 288440 318248 288492 318300
rect 297088 318248 297140 318300
rect 315028 318248 315080 318300
rect 328552 318248 328604 318300
rect 365904 318248 365956 318300
rect 247040 318180 247092 318232
rect 256792 318180 256844 318232
rect 272432 318180 272484 318232
rect 272616 318180 272668 318232
rect 281356 318180 281408 318232
rect 242440 318112 242492 318164
rect 281632 318112 281684 318164
rect 282184 318180 282236 318232
rect 291476 318180 291528 318232
rect 291844 318180 291896 318232
rect 293960 318180 294012 318232
rect 294144 318180 294196 318232
rect 295340 318180 295392 318232
rect 313464 318180 313516 318232
rect 324228 318180 324280 318232
rect 327540 318180 327592 318232
rect 328276 318180 328328 318232
rect 328460 318180 328512 318232
rect 368664 318180 368716 318232
rect 206836 318044 206888 318096
rect 269028 318044 269080 318096
rect 271236 318044 271288 318096
rect 283196 318044 283248 318096
rect 283932 318044 283984 318096
rect 285312 318112 285364 318164
rect 299940 318112 299992 318164
rect 316500 318112 316552 318164
rect 286600 318044 286652 318096
rect 286692 318044 286744 318096
rect 298008 318044 298060 318096
rect 328644 318112 328696 318164
rect 371516 318112 371568 318164
rect 330024 318044 330076 318096
rect 330760 318044 330812 318096
rect 381268 318044 381320 318096
rect 277032 317976 277084 318028
rect 287704 317976 287756 318028
rect 289452 317976 289504 318028
rect 281264 317908 281316 317960
rect 289820 317908 289872 317960
rect 292764 317976 292816 318028
rect 293040 317976 293092 318028
rect 297456 317976 297508 318028
rect 303344 317976 303396 318028
rect 303988 317976 304040 318028
rect 331404 317976 331456 318028
rect 354220 317976 354272 318028
rect 293684 317908 293736 317960
rect 346032 317908 346084 317960
rect 257068 317840 257120 317892
rect 257988 317840 258040 317892
rect 285128 317840 285180 317892
rect 286600 317840 286652 317892
rect 296996 317840 297048 317892
rect 297272 317840 297324 317892
rect 332140 317840 332192 317892
rect 265808 317772 265860 317824
rect 283012 317772 283064 317824
rect 290280 317772 290332 317824
rect 332232 317772 332284 317824
rect 270040 317704 270092 317756
rect 275560 317704 275612 317756
rect 293868 317704 293920 317756
rect 299572 317704 299624 317756
rect 300952 317704 301004 317756
rect 303988 317704 304040 317756
rect 307484 317704 307536 317756
rect 311256 317704 311308 317756
rect 324596 317704 324648 317756
rect 324964 317704 325016 317756
rect 284852 317636 284904 317688
rect 285036 317636 285088 317688
rect 286048 317636 286100 317688
rect 287336 317636 287388 317688
rect 291936 317636 291988 317688
rect 292304 317636 292356 317688
rect 333428 317636 333480 317688
rect 282828 317568 282880 317620
rect 288808 317568 288860 317620
rect 279884 317500 279936 317552
rect 296260 317568 296312 317620
rect 296720 317568 296772 317620
rect 299848 317568 299900 317620
rect 300584 317568 300636 317620
rect 300952 317568 301004 317620
rect 302148 317568 302200 317620
rect 314108 317568 314160 317620
rect 314568 317568 314620 317620
rect 325792 317568 325844 317620
rect 326528 317568 326580 317620
rect 327448 317568 327500 317620
rect 329104 317568 329156 317620
rect 295984 317500 296036 317552
rect 299664 317500 299716 317552
rect 314016 317500 314068 317552
rect 317328 317500 317380 317552
rect 321928 317500 321980 317552
rect 328828 317500 328880 317552
rect 276848 317432 276900 317484
rect 277216 317432 277268 317484
rect 280620 317432 280672 317484
rect 268844 317364 268896 317416
rect 269580 317364 269632 317416
rect 281080 317364 281132 317416
rect 283380 317364 283432 317416
rect 284208 317364 284260 317416
rect 285404 317432 285456 317484
rect 286876 317432 286928 317484
rect 287152 317364 287204 317416
rect 288348 317364 288400 317416
rect 290280 317432 290332 317484
rect 290464 317432 290516 317484
rect 297916 317432 297968 317484
rect 298376 317432 298428 317484
rect 302148 317432 302200 317484
rect 304724 317432 304776 317484
rect 307576 317432 307628 317484
rect 307944 317432 307996 317484
rect 313188 317432 313240 317484
rect 314108 317432 314160 317484
rect 320640 317432 320692 317484
rect 327816 317432 327868 317484
rect 298836 317364 298888 317416
rect 325608 317364 325660 317416
rect 394884 317364 394936 317416
rect 395988 317364 396040 317416
rect 270132 317296 270184 317348
rect 297548 317296 297600 317348
rect 322480 317296 322532 317348
rect 322664 317296 322716 317348
rect 329104 317296 329156 317348
rect 330116 317296 330168 317348
rect 389548 317296 389600 317348
rect 278688 317228 278740 317280
rect 298192 317228 298244 317280
rect 323584 317228 323636 317280
rect 324136 317228 324188 317280
rect 326160 317228 326212 317280
rect 332876 317228 332928 317280
rect 333704 317228 333756 317280
rect 340880 317228 340932 317280
rect 341984 317228 342036 317280
rect 279608 317160 279660 317212
rect 299020 317160 299072 317212
rect 309140 317160 309192 317212
rect 309416 317160 309468 317212
rect 328460 317160 328512 317212
rect 291292 317092 291344 317144
rect 292212 317092 292264 317144
rect 293684 317092 293736 317144
rect 299480 317092 299532 317144
rect 307024 317092 307076 317144
rect 328552 317092 328604 317144
rect 328828 317092 328880 317144
rect 329748 317092 329800 317144
rect 339316 317092 339368 317144
rect 277032 317024 277084 317076
rect 303344 317024 303396 317076
rect 317328 317024 317380 317076
rect 340972 317024 341024 317076
rect 277768 316956 277820 317008
rect 278688 316956 278740 317008
rect 279240 316956 279292 317008
rect 309140 316956 309192 317008
rect 317512 316956 317564 317008
rect 340880 316956 340932 317008
rect 275376 316888 275428 316940
rect 309416 316888 309468 316940
rect 321100 316888 321152 316940
rect 321284 316888 321336 316940
rect 324228 316888 324280 316940
rect 328552 316888 328604 316940
rect 329656 316888 329708 316940
rect 213552 316820 213604 316872
rect 270132 316820 270184 316872
rect 273904 316820 273956 316872
rect 311992 316820 312044 316872
rect 324136 316820 324188 316872
rect 328276 316820 328328 316872
rect 341340 316820 341392 316872
rect 347504 316820 347556 316872
rect 362316 316820 362368 316872
rect 212172 316752 212224 316804
rect 280160 316752 280212 316804
rect 309416 316752 309468 316804
rect 309600 316752 309652 316804
rect 324228 316752 324280 316804
rect 325976 316752 326028 316804
rect 212356 316684 212408 316736
rect 296076 316684 296128 316736
rect 296536 316684 296588 316736
rect 312728 316684 312780 316736
rect 347504 316684 347556 316736
rect 348792 316684 348844 316736
rect 385224 316684 385276 316736
rect 395988 316684 396040 316736
rect 527824 316684 527876 316736
rect 275744 316616 275796 316668
rect 276388 316616 276440 316668
rect 295064 316616 295116 316668
rect 298284 316616 298336 316668
rect 299296 316616 299348 316668
rect 304724 316616 304776 316668
rect 336648 316616 336700 316668
rect 272892 316548 272944 316600
rect 276296 316548 276348 316600
rect 304448 316548 304500 316600
rect 317512 316548 317564 316600
rect 317696 316548 317748 316600
rect 319444 316548 319496 316600
rect 320088 316548 320140 316600
rect 378324 316548 378376 316600
rect 296536 316480 296588 316532
rect 355048 316480 355100 316532
rect 303344 316412 303396 316464
rect 305276 316412 305328 316464
rect 329380 316412 329432 316464
rect 278504 316344 278556 316396
rect 303712 316344 303764 316396
rect 304724 316344 304776 316396
rect 316684 316344 316736 316396
rect 329472 316344 329524 316396
rect 294512 316208 294564 316260
rect 294972 316208 295024 316260
rect 298836 316208 298888 316260
rect 304448 316276 304500 316328
rect 313004 316276 313056 316328
rect 313188 316276 313240 316328
rect 321284 316276 321336 316328
rect 321468 316276 321520 316328
rect 324872 316276 324924 316328
rect 325608 316276 325660 316328
rect 272984 316140 273036 316192
rect 300860 316208 300912 316260
rect 301136 316208 301188 316260
rect 304172 316208 304224 316260
rect 304724 316208 304776 316260
rect 306656 316208 306708 316260
rect 307116 316208 307168 316260
rect 311440 316208 311492 316260
rect 311624 316208 311676 316260
rect 313740 316208 313792 316260
rect 316132 316208 316184 316260
rect 316408 316208 316460 316260
rect 311992 316140 312044 316192
rect 312176 316140 312228 316192
rect 313004 316140 313056 316192
rect 313556 316140 313608 316192
rect 314292 316140 314344 316192
rect 315028 316140 315080 316192
rect 315488 316140 315540 316192
rect 320456 316140 320508 316192
rect 321468 316140 321520 316192
rect 321836 316140 321888 316192
rect 322572 316140 322624 316192
rect 285680 316072 285732 316124
rect 286140 316072 286192 316124
rect 282552 316004 282604 316056
rect 294788 316004 294840 316056
rect 295064 316004 295116 316056
rect 303988 316072 304040 316124
rect 304448 316072 304500 316124
rect 323492 316072 323544 316124
rect 323676 316072 323728 316124
rect 299940 316004 299992 316056
rect 300676 316004 300728 316056
rect 302792 316004 302844 316056
rect 303436 316004 303488 316056
rect 304172 316004 304224 316056
rect 304816 316004 304868 316056
rect 305276 316004 305328 316056
rect 305920 316004 305972 316056
rect 306840 316004 306892 316056
rect 307300 316004 307352 316056
rect 308312 316004 308364 316056
rect 309048 316004 309100 316056
rect 310704 316004 310756 316056
rect 311716 316004 311768 316056
rect 312084 316004 312136 316056
rect 312912 316004 312964 316056
rect 313372 316004 313424 316056
rect 314292 316004 314344 316056
rect 314844 316004 314896 316056
rect 315856 316004 315908 316056
rect 316224 316004 316276 316056
rect 316960 316004 317012 316056
rect 324596 316004 324648 316056
rect 325148 316004 325200 316056
rect 264796 315936 264848 315988
rect 283472 315936 283524 315988
rect 284484 315936 284536 315988
rect 285588 315936 285640 315988
rect 285956 315936 286008 315988
rect 286968 315936 287020 315988
rect 287152 315936 287204 315988
rect 287796 315936 287848 315988
rect 288808 315936 288860 315988
rect 289360 315936 289412 315988
rect 291384 315936 291436 315988
rect 292396 315936 292448 315988
rect 292856 315936 292908 315988
rect 293500 315936 293552 315988
rect 294512 315936 294564 315988
rect 295156 315936 295208 315988
rect 295524 315936 295576 315988
rect 296168 315936 296220 315988
rect 296812 315936 296864 315988
rect 297548 315936 297600 315988
rect 299848 315936 299900 315988
rect 300400 315936 300452 315988
rect 302516 315936 302568 315988
rect 302884 315936 302936 315988
rect 303988 315936 304040 315988
rect 304356 315936 304408 315988
rect 307116 315936 307168 315988
rect 307392 315936 307444 315988
rect 308588 315936 308640 315988
rect 308864 315936 308916 315988
rect 309416 315936 309468 315988
rect 310428 315936 310480 315988
rect 310796 315936 310848 315988
rect 311072 315936 311124 315988
rect 312176 315936 312228 315988
rect 312820 315936 312872 315988
rect 314936 315936 314988 315988
rect 315948 315936 316000 315988
rect 316316 315936 316368 315988
rect 316776 315936 316828 315988
rect 317696 315936 317748 315988
rect 318432 315936 318484 315988
rect 320456 315936 320508 315988
rect 321376 315936 321428 315988
rect 323032 315936 323084 315988
rect 323400 315936 323452 315988
rect 324412 315936 324464 315988
rect 324780 315936 324832 315988
rect 288532 315868 288584 315920
rect 288900 315868 288952 315920
rect 288992 315868 289044 315920
rect 289636 315868 289688 315920
rect 299664 315868 299716 315920
rect 300768 315868 300820 315920
rect 303804 315868 303856 315920
rect 304908 315868 304960 315920
rect 309600 315868 309652 315920
rect 310336 315868 310388 315920
rect 310612 315868 310664 315920
rect 311716 315868 311768 315920
rect 312360 315868 312412 315920
rect 313096 315868 313148 315920
rect 314752 315868 314804 315920
rect 315580 315868 315632 315920
rect 318064 315868 318116 315920
rect 318524 315868 318576 315920
rect 324136 315868 324188 315920
rect 328644 315868 328696 315920
rect 285404 315800 285456 315852
rect 285588 315800 285640 315852
rect 287244 315800 287296 315852
rect 288256 315800 288308 315852
rect 288624 315800 288676 315852
rect 289360 315800 289412 315852
rect 278228 315664 278280 315716
rect 310520 315800 310572 315852
rect 310796 315800 310848 315852
rect 311808 315800 311860 315852
rect 312084 315800 312136 315852
rect 312544 315800 312596 315852
rect 296812 315732 296864 315784
rect 297732 315732 297784 315784
rect 302424 315732 302476 315784
rect 302976 315732 303028 315784
rect 309140 315732 309192 315784
rect 310244 315732 310296 315784
rect 319812 315800 319864 315852
rect 328184 315800 328236 315852
rect 302332 315664 302384 315716
rect 303068 315664 303120 315716
rect 281356 315596 281408 315648
rect 315764 315732 315816 315784
rect 375656 315732 375708 315784
rect 314384 315664 314436 315716
rect 375012 315664 375064 315716
rect 281264 315528 281316 315580
rect 319720 315596 319772 315648
rect 316408 315528 316460 315580
rect 317328 315528 317380 315580
rect 337752 315528 337804 315580
rect 213644 315460 213696 315512
rect 272616 315460 272668 315512
rect 275560 315460 275612 315512
rect 320732 315460 320784 315512
rect 246948 315392 247000 315444
rect 302240 315392 302292 315444
rect 302516 315392 302568 315444
rect 303528 315392 303580 315444
rect 307024 315392 307076 315444
rect 307484 315392 307536 315444
rect 213460 315324 213512 315376
rect 283840 315324 283892 315376
rect 285128 315324 285180 315376
rect 312452 315392 312504 315444
rect 336556 315392 336608 315444
rect 321008 315324 321060 315376
rect 331588 315324 331640 315376
rect 334992 315324 335044 315376
rect 219716 315256 219768 315308
rect 313648 315256 313700 315308
rect 328460 315256 328512 315308
rect 328828 315256 328880 315308
rect 385040 315256 385092 315308
rect 291936 315188 291988 315240
rect 317512 315188 317564 315240
rect 291660 315120 291712 315172
rect 292212 315120 292264 315172
rect 308772 315120 308824 315172
rect 327724 315120 327776 315172
rect 327816 315120 327868 315172
rect 328644 315120 328696 315172
rect 337844 315120 337896 315172
rect 314568 315052 314620 315104
rect 382740 315052 382792 315104
rect 317236 314984 317288 315036
rect 377128 314984 377180 315036
rect 313188 314916 313240 314968
rect 372896 314916 372948 314968
rect 287336 314848 287388 314900
rect 288164 314848 288216 314900
rect 292948 314848 293000 314900
rect 293592 314848 293644 314900
rect 317512 314848 317564 314900
rect 332416 314848 332468 314900
rect 317328 314780 317380 314832
rect 352656 314780 352708 314832
rect 302240 314712 302292 314764
rect 306472 314712 306524 314764
rect 328736 314712 328788 314764
rect 248144 314644 248196 314696
rect 307024 314644 307076 314696
rect 327816 314644 327868 314696
rect 328276 314644 328328 314696
rect 274548 314576 274600 314628
rect 306380 314576 306432 314628
rect 308404 314576 308456 314628
rect 329288 314576 329340 314628
rect 275928 314508 275980 314560
rect 305000 314508 305052 314560
rect 317880 314508 317932 314560
rect 318432 314508 318484 314560
rect 284300 314440 284352 314492
rect 285220 314440 285272 314492
rect 297640 314440 297692 314492
rect 298008 314440 298060 314492
rect 311992 314440 312044 314492
rect 333612 314508 333664 314560
rect 318616 314440 318668 314492
rect 379152 314440 379204 314492
rect 296260 314372 296312 314424
rect 356152 314372 356204 314424
rect 299480 314304 299532 314356
rect 300860 314304 300912 314356
rect 360660 314304 360712 314356
rect 270224 314236 270276 314288
rect 300308 314236 300360 314288
rect 318432 314236 318484 314288
rect 376944 314236 376996 314288
rect 260472 314168 260524 314220
rect 260656 314168 260708 314220
rect 297640 314168 297692 314220
rect 341892 314168 341944 314220
rect 298008 314100 298060 314152
rect 300584 314100 300636 314152
rect 332324 314100 332376 314152
rect 222200 314032 222252 314084
rect 242440 314032 242492 314084
rect 248052 314032 248104 314084
rect 308496 314032 308548 314084
rect 311256 314032 311308 314084
rect 341432 314032 341484 314084
rect 210976 313964 211028 314016
rect 271420 313964 271472 314016
rect 211896 313896 211948 313948
rect 273720 313896 273772 313948
rect 274548 313896 274600 313948
rect 282460 313896 282512 313948
rect 321100 313964 321152 314016
rect 330024 313964 330076 314016
rect 390836 313964 390888 314016
rect 336280 313896 336332 313948
rect 379244 313896 379296 313948
rect 466460 313896 466512 313948
rect 310520 313828 310572 313880
rect 311348 313828 311400 313880
rect 329840 313828 329892 313880
rect 317880 313760 317932 313812
rect 318708 313760 318760 313812
rect 379244 313760 379296 313812
rect 319444 313692 319496 313744
rect 319812 313692 319864 313744
rect 379704 313692 379756 313744
rect 298744 313624 298796 313676
rect 330668 313624 330720 313676
rect 279792 313556 279844 313608
rect 284300 313556 284352 313608
rect 279424 313420 279476 313472
rect 286048 313420 286100 313472
rect 292672 313420 292724 313472
rect 293408 313420 293460 313472
rect 275744 313352 275796 313404
rect 287704 313352 287756 313404
rect 270224 313284 270276 313336
rect 270684 313284 270736 313336
rect 272616 313284 272668 313336
rect 312452 313284 312504 313336
rect 260564 313216 260616 313268
rect 260748 313216 260800 313268
rect 287060 313216 287112 313268
rect 309876 313216 309928 313268
rect 310428 313216 310480 313268
rect 322112 313216 322164 313268
rect 389272 313216 389324 313268
rect 523684 313216 523736 313268
rect 579620 313216 579672 313268
rect 305644 313148 305696 313200
rect 330576 313148 330628 313200
rect 313096 313080 313148 313132
rect 372804 313080 372856 313132
rect 309692 313012 309744 313064
rect 310060 313012 310112 313064
rect 329932 313012 329984 313064
rect 294880 312944 294932 312996
rect 341800 312944 341852 312996
rect 295432 312876 295484 312928
rect 331036 312876 331088 312928
rect 315212 312808 315264 312860
rect 350172 312808 350224 312860
rect 202696 312740 202748 312792
rect 260748 312740 260800 312792
rect 253664 312672 253716 312724
rect 313096 312672 313148 312724
rect 252468 312604 252520 312656
rect 312820 312604 312872 312656
rect 210608 312536 210660 312588
rect 278412 312536 278464 312588
rect 278688 312536 278740 312588
rect 322848 312740 322900 312792
rect 329840 312740 329892 312792
rect 330944 312740 330996 312792
rect 317144 312672 317196 312724
rect 343364 312740 343416 312792
rect 328368 312604 328420 312656
rect 333152 312604 333204 312656
rect 387892 312604 387944 312656
rect 322848 312536 322900 312588
rect 336188 312536 336240 312588
rect 301504 312468 301556 312520
rect 301872 312468 301924 312520
rect 335084 312468 335136 312520
rect 305000 312400 305052 312452
rect 305644 312400 305696 312452
rect 321008 312400 321060 312452
rect 321284 312400 321336 312452
rect 381360 312400 381412 312452
rect 502340 312536 502392 312588
rect 277860 312332 277912 312384
rect 322112 312332 322164 312384
rect 322756 312332 322808 312384
rect 371884 312332 371936 312384
rect 310428 312196 310480 312248
rect 336372 312264 336424 312316
rect 312820 312128 312872 312180
rect 321560 312128 321612 312180
rect 262036 311788 262088 311840
rect 287244 311788 287296 311840
rect 295340 311788 295392 311840
rect 297916 311788 297968 311840
rect 333244 311788 333296 311840
rect 266360 311720 266412 311772
rect 267556 311720 267608 311772
rect 287428 311720 287480 311772
rect 299112 311720 299164 311772
rect 358084 311720 358136 311772
rect 293040 311652 293092 311704
rect 293408 311652 293460 311704
rect 352380 311652 352432 311704
rect 287796 311448 287848 311500
rect 301596 311516 301648 311568
rect 313740 311584 313792 311636
rect 369768 311584 369820 311636
rect 374092 311584 374144 311636
rect 355600 311516 355652 311568
rect 304356 311448 304408 311500
rect 306012 311448 306064 311500
rect 311532 311448 311584 311500
rect 313740 311448 313792 311500
rect 321560 311448 321612 311500
rect 371424 311448 371476 311500
rect 289176 311380 289228 311432
rect 298008 311380 298060 311432
rect 300768 311380 300820 311432
rect 346216 311380 346268 311432
rect 287980 311312 288032 311364
rect 288900 311244 288952 311296
rect 289084 311244 289136 311296
rect 293224 311312 293276 311364
rect 336096 311312 336148 311364
rect 299848 311244 299900 311296
rect 300676 311244 300728 311296
rect 219164 311176 219216 311228
rect 262036 311176 262088 311228
rect 282736 311176 282788 311228
rect 298284 311176 298336 311228
rect 299112 311176 299164 311228
rect 299940 311176 299992 311228
rect 342904 311244 342956 311296
rect 209412 311108 209464 311160
rect 266360 311108 266412 311160
rect 285036 311108 285088 311160
rect 300216 311108 300268 311160
rect 300768 311108 300820 311160
rect 300676 310972 300728 311024
rect 339132 311176 339184 311228
rect 310888 311108 310940 311160
rect 311256 311108 311308 311160
rect 315948 311108 316000 311160
rect 351552 311108 351604 311160
rect 311072 311040 311124 311092
rect 311808 311040 311860 311092
rect 347412 311040 347464 311092
rect 308312 310972 308364 311024
rect 342352 310972 342404 311024
rect 311256 310904 311308 310956
rect 371240 310904 371292 310956
rect 271696 310496 271748 310548
rect 291108 310496 291160 310548
rect 315028 310496 315080 310548
rect 315948 310496 316000 310548
rect 259368 310428 259420 310480
rect 284484 310428 284536 310480
rect 299112 310428 299164 310480
rect 305092 310428 305144 310480
rect 333520 310428 333572 310480
rect 283288 310360 283340 310412
rect 283564 310360 283616 310412
rect 297364 310360 297416 310412
rect 305000 310360 305052 310412
rect 317512 310360 317564 310412
rect 327724 310360 327776 310412
rect 341708 310360 341760 310412
rect 381176 310292 381228 310344
rect 313556 310224 313608 310276
rect 374920 310224 374972 310276
rect 330392 310156 330444 310208
rect 383752 310156 383804 310208
rect 297824 310088 297876 310140
rect 298928 310088 298980 310140
rect 356796 310088 356848 310140
rect 286508 310020 286560 310072
rect 295432 310020 295484 310072
rect 313924 310020 313976 310072
rect 373264 310020 373316 310072
rect 286876 309952 286928 310004
rect 297180 309952 297232 310004
rect 355324 309952 355376 310004
rect 226064 309884 226116 309936
rect 259368 309884 259420 309936
rect 219072 309816 219124 309868
rect 295708 309816 295760 309868
rect 340512 309884 340564 309936
rect 342352 309884 342404 309936
rect 342904 309884 342956 309936
rect 369216 309884 369268 309936
rect 302884 309816 302936 309868
rect 344836 309816 344888 309868
rect 217784 309748 217836 309800
rect 294512 309748 294564 309800
rect 338948 309748 339000 309800
rect 316960 309680 317012 309732
rect 354128 309680 354180 309732
rect 316224 309612 316276 309664
rect 390744 309612 390796 309664
rect 310980 309544 311032 309596
rect 311532 309544 311584 309596
rect 319996 309544 320048 309596
rect 387800 309544 387852 309596
rect 283564 309476 283616 309528
rect 328000 309476 328052 309528
rect 323676 309408 323728 309460
rect 330392 309408 330444 309460
rect 275928 309204 275980 309256
rect 285680 309204 285732 309256
rect 316316 309204 316368 309256
rect 316960 309204 317012 309256
rect 327172 309204 327224 309256
rect 327540 309204 327592 309256
rect 274548 309136 274600 309188
rect 288256 309136 288308 309188
rect 260472 309068 260524 309120
rect 260748 309068 260800 309120
rect 285956 309068 286008 309120
rect 300308 309068 300360 309120
rect 302148 309068 302200 309120
rect 302792 309068 302844 309120
rect 302976 309068 303028 309120
rect 316224 309136 316276 309188
rect 316684 309136 316736 309188
rect 317512 309136 317564 309188
rect 318524 309136 318576 309188
rect 364616 309068 364668 309120
rect 270408 309000 270460 309052
rect 288072 309000 288124 309052
rect 302608 309000 302660 309052
rect 303160 309000 303212 309052
rect 310796 309000 310848 309052
rect 311348 309000 311400 309052
rect 371332 309000 371384 309052
rect 301688 308932 301740 308984
rect 304172 308932 304224 308984
rect 364524 308932 364576 308984
rect 302976 308864 303028 308916
rect 360936 308864 360988 308916
rect 303160 308796 303212 308848
rect 359648 308796 359700 308848
rect 293960 308728 294012 308780
rect 294420 308728 294472 308780
rect 350080 308728 350132 308780
rect 294052 308660 294104 308712
rect 294328 308660 294380 308712
rect 348884 308660 348936 308712
rect 207940 308592 207992 308644
rect 270408 308592 270460 308644
rect 304080 308592 304132 308644
rect 304448 308592 304500 308644
rect 355508 308592 355560 308644
rect 219808 308524 219860 308576
rect 260748 308524 260800 308576
rect 264888 308524 264940 308576
rect 332968 308524 333020 308576
rect 259644 308456 259696 308508
rect 332600 308456 332652 308508
rect 217416 308388 217468 308440
rect 293960 308388 294012 308440
rect 300216 308388 300268 308440
rect 302700 308388 302752 308440
rect 340604 308388 340656 308440
rect 371332 308388 371384 308440
rect 372160 308388 372212 308440
rect 378140 308388 378192 308440
rect 305276 308320 305328 308372
rect 305828 308320 305880 308372
rect 340420 308320 340472 308372
rect 292948 308252 293000 308304
rect 298284 308252 298336 308304
rect 331956 308252 332008 308304
rect 319628 308184 319680 308236
rect 339224 308184 339276 308236
rect 216128 307844 216180 307896
rect 292948 307844 293000 307896
rect 216220 307776 216272 307828
rect 293960 307776 294012 307828
rect 263140 307708 263192 307760
rect 263416 307708 263468 307760
rect 283196 307708 283248 307760
rect 287704 307640 287756 307692
rect 303988 307640 304040 307692
rect 338672 307708 338724 307760
rect 310704 307640 310756 307692
rect 311440 307640 311492 307692
rect 323768 307640 323820 307692
rect 334072 307640 334124 307692
rect 335268 307640 335320 307692
rect 292948 307572 293000 307624
rect 293316 307572 293368 307624
rect 351368 307572 351420 307624
rect 291108 307504 291160 307556
rect 348424 307504 348476 307556
rect 281908 307436 281960 307488
rect 299480 307436 299532 307488
rect 356704 307436 356756 307488
rect 280712 307368 280764 307420
rect 290832 307368 290884 307420
rect 291108 307368 291160 307420
rect 294236 307368 294288 307420
rect 347136 307368 347188 307420
rect 285220 307300 285272 307352
rect 298100 307300 298152 307352
rect 344560 307300 344612 307352
rect 285496 307232 285548 307284
rect 331864 307232 331916 307284
rect 213368 307164 213420 307216
rect 263140 307164 263192 307216
rect 283840 307164 283892 307216
rect 217508 307096 217560 307148
rect 293224 307096 293276 307148
rect 293960 307164 294012 307216
rect 294972 307164 295024 307216
rect 337660 307164 337712 307216
rect 294052 307096 294104 307148
rect 314476 307096 314528 307148
rect 355416 307096 355468 307148
rect 217600 307028 217652 307080
rect 299940 307028 299992 307080
rect 314936 307028 314988 307080
rect 315580 307028 315632 307080
rect 376300 307028 376352 307080
rect 431960 307028 432012 307080
rect 311440 306960 311492 307012
rect 370504 306960 370556 307012
rect 313556 306892 313608 306944
rect 314476 306892 314528 306944
rect 209228 306348 209280 306400
rect 267004 306348 267056 306400
rect 266360 306280 266412 306332
rect 267648 306280 267700 306332
rect 286416 306280 286468 306332
rect 305184 306280 305236 306332
rect 365812 306280 365864 306332
rect 308220 306212 308272 306264
rect 367928 306212 367980 306264
rect 308128 306144 308180 306196
rect 367836 306144 367888 306196
rect 293224 306076 293276 306128
rect 309784 306076 309836 306128
rect 365076 306076 365128 306128
rect 285864 306008 285916 306060
rect 339040 306008 339092 306060
rect 296076 305940 296128 305992
rect 308128 305940 308180 305992
rect 309600 305940 309652 305992
rect 362224 305940 362276 305992
rect 292856 305872 292908 305924
rect 344284 305872 344336 305924
rect 286324 305804 286376 305856
rect 302516 305804 302568 305856
rect 348700 305804 348752 305856
rect 291476 305736 291528 305788
rect 336004 305736 336056 305788
rect 210700 305668 210752 305720
rect 266360 305668 266412 305720
rect 214840 305600 214892 305652
rect 292856 305600 292908 305652
rect 290096 305532 290148 305584
rect 291016 305532 291068 305584
rect 330484 305668 330536 305720
rect 307392 305600 307444 305652
rect 343088 305600 343140 305652
rect 299756 305396 299808 305448
rect 300584 305396 300636 305448
rect 334900 305532 334952 305584
rect 322756 305464 322808 305516
rect 349896 305464 349948 305516
rect 306748 305396 306800 305448
rect 307392 305396 307444 305448
rect 314108 305396 314160 305448
rect 339592 305396 339644 305448
rect 321652 305124 321704 305176
rect 322756 305124 322808 305176
rect 216036 305056 216088 305108
rect 259644 305056 259696 305108
rect 206284 304988 206336 305040
rect 265900 304988 265952 305040
rect 288164 304988 288216 305040
rect 291476 304988 291528 305040
rect 305184 304988 305236 305040
rect 305644 304988 305696 305040
rect 308220 304988 308272 305040
rect 308588 304988 308640 305040
rect 339592 304988 339644 305040
rect 340788 304988 340840 305040
rect 282644 304920 282696 304972
rect 359556 304920 359608 304972
rect 264980 304852 265032 304904
rect 266176 304852 266228 304904
rect 288992 304852 289044 304904
rect 295340 304852 295392 304904
rect 295616 304852 295668 304904
rect 357072 304852 357124 304904
rect 271788 304784 271840 304836
rect 291384 304784 291436 304836
rect 302424 304784 302476 304836
rect 360844 304784 360896 304836
rect 267004 304716 267056 304768
rect 283104 304716 283156 304768
rect 300952 304716 301004 304768
rect 351276 304716 351328 304768
rect 299664 304648 299716 304700
rect 349804 304648 349856 304700
rect 261300 304580 261352 304632
rect 261760 304580 261812 304632
rect 298652 304580 298704 304632
rect 347320 304580 347372 304632
rect 220636 304512 220688 304564
rect 271788 304512 271840 304564
rect 286692 304512 286744 304564
rect 301228 304512 301280 304564
rect 348516 304512 348568 304564
rect 208124 304444 208176 304496
rect 264980 304444 265032 304496
rect 293316 304444 293368 304496
rect 300952 304444 301004 304496
rect 301136 304444 301188 304496
rect 345940 304444 345992 304496
rect 218888 304376 218940 304428
rect 208032 304308 208084 304360
rect 285864 304308 285916 304360
rect 301044 304376 301096 304428
rect 344468 304376 344520 304428
rect 296904 304308 296956 304360
rect 340328 304308 340380 304360
rect 213276 304240 213328 304292
rect 295340 304240 295392 304292
rect 299572 304240 299624 304292
rect 348608 304240 348660 304292
rect 300492 304172 300544 304224
rect 341616 304172 341668 304224
rect 299112 304104 299164 304156
rect 334716 304104 334768 304156
rect 284116 304036 284168 304088
rect 302424 304036 302476 304088
rect 307024 304036 307076 304088
rect 313188 304036 313240 304088
rect 334808 304036 334860 304088
rect 298560 303968 298612 304020
rect 299572 303968 299624 304020
rect 204536 303696 204588 303748
rect 264060 303764 264112 303816
rect 264520 303764 264572 303816
rect 297456 303696 297508 303748
rect 301136 303696 301188 303748
rect 201408 303628 201460 303680
rect 261300 303628 261352 303680
rect 298652 303628 298704 303680
rect 299020 303628 299072 303680
rect 299664 303628 299716 303680
rect 300124 303628 300176 303680
rect 301044 303628 301096 303680
rect 301596 303628 301648 303680
rect 317512 303560 317564 303612
rect 390560 303560 390612 303612
rect 320732 303492 320784 303544
rect 320916 303492 320968 303544
rect 390652 303492 390704 303544
rect 301780 303424 301832 303476
rect 362132 303424 362184 303476
rect 320916 303356 320968 303408
rect 321100 303356 321152 303408
rect 321192 303356 321244 303408
rect 380164 303356 380216 303408
rect 320180 303288 320232 303340
rect 321468 303288 321520 303340
rect 380072 303288 380124 303340
rect 321100 303220 321152 303272
rect 321284 303220 321336 303272
rect 321376 303220 321428 303272
rect 380348 303220 380400 303272
rect 295340 303152 295392 303204
rect 296444 303152 296496 303204
rect 354036 303152 354088 303204
rect 292028 303084 292080 303136
rect 294144 303084 294196 303136
rect 351184 303084 351236 303136
rect 288256 303016 288308 303068
rect 295524 303016 295576 303068
rect 352564 303016 352616 303068
rect 213828 302948 213880 303000
rect 291752 302948 291804 303000
rect 340236 302948 340288 303000
rect 215944 302880 215996 302932
rect 295340 302880 295392 302932
rect 298008 302880 298060 302932
rect 337476 302880 337528 302932
rect 305368 302812 305420 302864
rect 329196 302812 329248 302864
rect 301964 302744 302016 302796
rect 303896 302744 303948 302796
rect 343180 302744 343232 302796
rect 300032 302676 300084 302728
rect 343272 302676 343324 302728
rect 204352 302268 204404 302320
rect 200120 302200 200172 302252
rect 260932 302200 260984 302252
rect 264520 302200 264572 302252
rect 264888 302200 264940 302252
rect 296812 302200 296864 302252
rect 298008 302200 298060 302252
rect 269948 302132 270000 302184
rect 297548 302132 297600 302184
rect 360568 302132 360620 302184
rect 289360 302064 289412 302116
rect 296352 302064 296404 302116
rect 357808 302064 357860 302116
rect 312912 301996 312964 302048
rect 374460 301996 374512 302048
rect 309784 301928 309836 301980
rect 371700 301928 371752 301980
rect 307208 301860 307260 301912
rect 307668 301860 307720 301912
rect 368848 301860 368900 301912
rect 300768 301792 300820 301844
rect 361948 301792 362000 301844
rect 297548 301724 297600 301776
rect 297916 301724 297968 301776
rect 309232 301724 309284 301776
rect 310152 301724 310204 301776
rect 309324 301656 309376 301708
rect 309784 301656 309836 301708
rect 370320 301724 370372 301776
rect 312084 301656 312136 301708
rect 312360 301656 312412 301708
rect 372252 301656 372304 301708
rect 309416 301588 309468 301640
rect 310244 301588 310296 301640
rect 310336 301588 310388 301640
rect 369032 301588 369084 301640
rect 287520 301520 287572 301572
rect 287888 301520 287940 301572
rect 345664 301520 345716 301572
rect 224316 301452 224368 301504
rect 293408 301452 293460 301504
rect 298376 301452 298428 301504
rect 351460 301452 351512 301504
rect 305920 301384 305972 301436
rect 344376 301384 344428 301436
rect 256700 301316 256752 301368
rect 257252 301316 257304 301368
rect 262312 301316 262364 301368
rect 262956 301316 263008 301368
rect 320732 301316 320784 301368
rect 321284 301316 321336 301368
rect 197360 300908 197412 300960
rect 256700 300908 256752 300960
rect 202788 300840 202840 300892
rect 262312 300840 262364 300892
rect 255320 300772 255372 300824
rect 256148 300772 256200 300824
rect 262404 300772 262456 300824
rect 262864 300772 262916 300824
rect 308036 300772 308088 300824
rect 308680 300772 308732 300824
rect 307484 300704 307536 300756
rect 369860 300772 369912 300824
rect 312636 300704 312688 300756
rect 313004 300704 313056 300756
rect 374368 300704 374420 300756
rect 300400 300636 300452 300688
rect 306012 300636 306064 300688
rect 367652 300636 367704 300688
rect 304632 300568 304684 300620
rect 364892 300568 364944 300620
rect 302332 300500 302384 300552
rect 302976 300500 303028 300552
rect 363880 300500 363932 300552
rect 307668 300432 307720 300484
rect 366548 300432 366600 300484
rect 318708 300364 318760 300416
rect 377956 300364 378008 300416
rect 306932 300296 306984 300348
rect 363604 300296 363656 300348
rect 289084 300092 289136 300144
rect 303804 300228 303856 300280
rect 359464 300228 359516 300280
rect 305736 300160 305788 300212
rect 306564 300160 306616 300212
rect 307668 300160 307720 300212
rect 307760 300160 307812 300212
rect 349988 300160 350040 300212
rect 304356 300092 304408 300144
rect 345848 300092 345900 300144
rect 230756 300024 230808 300076
rect 231768 300024 231820 300076
rect 307208 300024 307260 300076
rect 307668 300024 307720 300076
rect 308680 300024 308732 300076
rect 340144 300024 340196 300076
rect 209044 299684 209096 299736
rect 253204 299684 253256 299736
rect 195980 299616 196032 299668
rect 256148 299616 256200 299668
rect 201684 299548 201736 299600
rect 262404 299548 262456 299600
rect 231768 299480 231820 299532
rect 577504 299480 577556 299532
rect 310336 299412 310388 299464
rect 371608 299412 371660 299464
rect 316132 299344 316184 299396
rect 316776 299344 316828 299396
rect 317420 299344 317472 299396
rect 318064 299344 318116 299396
rect 318708 299344 318760 299396
rect 378692 299344 378744 299396
rect 295064 299276 295116 299328
rect 353944 299276 353996 299328
rect 310152 299208 310204 299260
rect 310336 299208 310388 299260
rect 310060 299140 310112 299192
rect 314292 299140 314344 299192
rect 372712 299208 372764 299260
rect 318064 299140 318116 299192
rect 377680 299140 377732 299192
rect 316776 299072 316828 299124
rect 376208 299072 376260 299124
rect 311716 299004 311768 299056
rect 364984 299004 365036 299056
rect 285588 298936 285640 298988
rect 337568 298936 337620 298988
rect 4160 298800 4212 298852
rect 221924 298800 221976 298852
rect 233148 298732 233200 298784
rect 580172 298732 580224 298784
rect 207848 298256 207900 298308
rect 265624 298256 265676 298308
rect 202880 298188 202932 298240
rect 263048 298188 263100 298240
rect 194600 298120 194652 298172
rect 254768 298120 254820 298172
rect 233700 298052 233752 298104
rect 233976 298052 234028 298104
rect 255964 298052 256016 298104
rect 256332 298052 256384 298104
rect 259276 298052 259328 298104
rect 265716 298052 265768 298104
rect 282828 298052 282880 298104
rect 349068 298052 349120 298104
rect 287152 297984 287204 298036
rect 303252 297984 303304 298036
rect 366180 297984 366232 298036
rect 307944 297916 307996 297968
rect 308496 297916 308548 297968
rect 309048 297916 309100 297968
rect 370228 297916 370280 297968
rect 304724 297848 304776 297900
rect 363420 297848 363472 297900
rect 305460 297780 305512 297832
rect 306104 297780 306156 297832
rect 364800 297780 364852 297832
rect 308496 297712 308548 297764
rect 368204 297712 368256 297764
rect 309048 297644 309100 297696
rect 347228 297644 347280 297696
rect 308956 297576 309008 297628
rect 345756 297576 345808 297628
rect 264060 297440 264112 297492
rect 264244 297440 264296 297492
rect 209136 297372 209188 297424
rect 236644 297372 236696 297424
rect 218796 297304 218848 297356
rect 258724 297304 258776 297356
rect 211804 297236 211856 297288
rect 256332 297236 256384 297288
rect 179420 297168 179472 297220
rect 238116 297168 238168 297220
rect 248604 297168 248656 297220
rect 249064 297168 249116 297220
rect 282092 297168 282144 297220
rect 282828 297168 282880 297220
rect 204444 297100 204496 297152
rect 264336 297100 264388 297152
rect 173900 297032 173952 297084
rect 233700 297032 233752 297084
rect 186320 296964 186372 297016
rect 246396 296964 246448 297016
rect 175280 296896 175332 296948
rect 235356 296896 235408 296948
rect 187700 296828 187752 296880
rect 248604 296828 248656 296880
rect 183560 296760 183612 296812
rect 244556 296760 244608 296812
rect 245016 296760 245068 296812
rect 206652 296692 206704 296744
rect 284576 296692 284628 296744
rect 288716 296624 288768 296676
rect 348976 296624 349028 296676
rect 288348 296556 288400 296608
rect 342996 296556 343048 296608
rect 230572 296148 230624 296200
rect 231216 296148 231268 296200
rect 240048 296080 240100 296132
rect 265992 296080 266044 296132
rect 242808 296012 242860 296064
rect 273168 296012 273220 296064
rect 222292 295944 222344 295996
rect 283564 295944 283616 295996
rect 169760 295876 169812 295928
rect 230572 295876 230624 295928
rect 214748 295808 214800 295860
rect 243360 295808 243412 295860
rect 186964 295740 187016 295792
rect 234896 295740 234948 295792
rect 202144 295672 202196 295724
rect 261668 295672 261720 295724
rect 182180 295604 182232 295656
rect 242164 295604 242216 295656
rect 178040 295536 178092 295588
rect 239036 295536 239088 295588
rect 240048 295536 240100 295588
rect 172520 295468 172572 295520
rect 233516 295468 233568 295520
rect 233884 295468 233936 295520
rect 234988 295468 235040 295520
rect 239404 295468 239456 295520
rect 214656 295400 214708 295452
rect 241980 295400 242032 295452
rect 242808 295400 242860 295452
rect 189080 295332 189132 295384
rect 250536 295332 250588 295384
rect 243084 295264 243136 295316
rect 243360 295264 243412 295316
rect 273076 295264 273128 295316
rect 284024 295264 284076 295316
rect 341524 295264 341576 295316
rect 288624 295196 288676 295248
rect 347044 295196 347096 295248
rect 284576 295128 284628 295180
rect 338856 295128 338908 295180
rect 193220 294788 193272 294840
rect 254492 294788 254544 294840
rect 234252 294720 234304 294772
rect 264612 294720 264664 294772
rect 167000 294652 167052 294704
rect 227996 294652 228048 294704
rect 228456 294652 228508 294704
rect 240048 294652 240100 294704
rect 275192 294652 275244 294704
rect 164516 294584 164568 294636
rect 222016 294584 222068 294636
rect 238392 294584 238444 294636
rect 277952 294584 278004 294636
rect 165896 294516 165948 294568
rect 227076 294516 227128 294568
rect 170404 294448 170456 294500
rect 225696 294448 225748 294500
rect 169852 294380 169904 294432
rect 229836 294380 229888 294432
rect 230204 294380 230256 294432
rect 180800 294312 180852 294364
rect 241612 294312 241664 294364
rect 171140 294244 171192 294296
rect 232412 294244 232464 294296
rect 168380 294176 168432 294228
rect 229100 294176 229152 294228
rect 229376 294176 229428 294228
rect 212080 294108 212132 294160
rect 234252 294108 234304 294160
rect 215024 294040 215076 294092
rect 247040 294040 247092 294092
rect 222016 293972 222068 294024
rect 225052 293972 225104 294024
rect 225696 293972 225748 294024
rect 225972 293972 226024 294024
rect 178132 293632 178184 293684
rect 237380 293632 237432 293684
rect 178224 293564 178276 293616
rect 238392 293564 238444 293616
rect 199660 293496 199712 293548
rect 256976 293496 257028 293548
rect 257344 293496 257396 293548
rect 237472 293360 237524 293412
rect 275836 293360 275888 293412
rect 231952 293292 232004 293344
rect 236460 293292 236512 293344
rect 278596 293292 278648 293344
rect 162676 293224 162728 293276
rect 220360 293224 220412 293276
rect 226524 293224 226576 293276
rect 235356 293224 235408 293276
rect 278136 293224 278188 293276
rect 212264 293156 212316 293208
rect 232044 293156 232096 293208
rect 217232 293088 217284 293140
rect 241888 293088 241940 293140
rect 200764 293020 200816 293072
rect 231952 293020 232004 293072
rect 232044 293020 232096 293072
rect 233148 293020 233200 293072
rect 259644 293020 259696 293072
rect 260196 293020 260248 293072
rect 262312 293020 262364 293072
rect 263140 293020 263192 293072
rect 189724 292952 189776 293004
rect 240048 292952 240100 293004
rect 178684 292884 178736 292936
rect 237472 292884 237524 292936
rect 172612 292816 172664 292868
rect 232780 292816 232832 292868
rect 238024 292816 238076 292868
rect 171232 292748 171284 292800
rect 231124 292748 231176 292800
rect 231308 292748 231360 292800
rect 218520 292680 218572 292732
rect 226984 292680 227036 292732
rect 219256 292612 219308 292664
rect 227720 292612 227772 292664
rect 3424 292544 3476 292596
rect 198740 292544 198792 292596
rect 199660 292544 199712 292596
rect 217692 292544 217744 292596
rect 235356 292544 235408 292596
rect 226984 292476 227036 292528
rect 228732 292476 228784 292528
rect 241888 292476 241940 292528
rect 275652 292476 275704 292528
rect 307208 292476 307260 292528
rect 314108 292476 314160 292528
rect 372620 292476 372672 292528
rect 373172 292476 373224 292528
rect 227720 292408 227772 292460
rect 228364 292408 228416 292460
rect 229836 292408 229888 292460
rect 247040 292408 247092 292460
rect 247500 292408 247552 292460
rect 281172 292408 281224 292460
rect 241612 292340 241664 292392
rect 271328 292340 271380 292392
rect 219992 292272 220044 292324
rect 237380 292204 237432 292256
rect 238300 292204 238352 292256
rect 189908 292136 189960 292188
rect 246304 292136 246356 292188
rect 227720 292068 227772 292120
rect 233148 292068 233200 292120
rect 256976 292272 257028 292324
rect 249340 292204 249392 292256
rect 258540 292204 258592 292256
rect 258724 292272 258776 292324
rect 260012 292272 260064 292324
rect 263048 292272 263100 292324
rect 264060 292272 264112 292324
rect 264520 292272 264572 292324
rect 265532 292272 265584 292324
rect 258908 292204 258960 292256
rect 264336 292204 264388 292256
rect 265164 292204 265216 292256
rect 257068 292136 257120 292188
rect 257436 292136 257488 292188
rect 258172 292136 258224 292188
rect 268476 292136 268528 292188
rect 271972 292136 272024 292188
rect 249340 292068 249392 292120
rect 252836 292068 252888 292120
rect 263968 292068 264020 292120
rect 245292 292000 245344 292052
rect 267280 292000 267332 292052
rect 218612 291932 218664 291984
rect 222108 291932 222160 291984
rect 227260 291932 227312 291984
rect 242716 291932 242768 291984
rect 250444 291932 250496 291984
rect 252560 291932 252612 291984
rect 282276 291932 282328 291984
rect 308864 291932 308916 291984
rect 336372 291932 336424 291984
rect 214564 291864 214616 291916
rect 234988 291864 235040 291916
rect 247868 291864 247920 291916
rect 279332 291864 279384 291916
rect 309140 291864 309192 291916
rect 310520 291864 310572 291916
rect 355968 291864 356020 291916
rect 357440 291864 357492 291916
rect 166908 291796 166960 291848
rect 220452 291796 220504 291848
rect 220728 291796 220780 291848
rect 220820 291796 220872 291848
rect 215852 291728 215904 291780
rect 231676 291796 231728 291848
rect 236828 291796 236880 291848
rect 264428 291796 264480 291848
rect 272432 291796 272484 291848
rect 331680 291796 331732 291848
rect 372620 291796 372672 291848
rect 402980 291796 403032 291848
rect 221004 291728 221056 291780
rect 243636 291728 243688 291780
rect 256148 291728 256200 291780
rect 256700 291728 256752 291780
rect 256792 291728 256844 291780
rect 259736 291728 259788 291780
rect 222016 291660 222068 291712
rect 244188 291660 244240 291712
rect 254492 291660 254544 291712
rect 220360 291592 220412 291644
rect 247776 291592 247828 291644
rect 254768 291592 254820 291644
rect 255596 291592 255648 291644
rect 271880 291660 271932 291712
rect 272524 291660 272576 291712
rect 281448 291592 281500 291644
rect 220084 291524 220136 291576
rect 247408 291524 247460 291576
rect 220820 291456 220872 291508
rect 253296 291456 253348 291508
rect 253756 291456 253808 291508
rect 220912 291388 220964 291440
rect 254584 291388 254636 291440
rect 221280 291320 221332 291372
rect 255964 291320 256016 291372
rect 264796 291320 264848 291372
rect 268384 291320 268436 291372
rect 269028 291320 269080 291372
rect 217324 291252 217376 291304
rect 228548 291252 228600 291304
rect 221372 291184 221424 291236
rect 235448 291184 235500 291236
rect 236092 291184 236144 291236
rect 238116 291184 238168 291236
rect 239404 291184 239456 291236
rect 240876 291252 240928 291304
rect 241888 291252 241940 291304
rect 263692 291252 263744 291304
rect 272432 291252 272484 291304
rect 242716 291184 242768 291236
rect 244280 291184 244332 291236
rect 244924 291184 244976 291236
rect 247776 291184 247828 291236
rect 248236 291184 248288 291236
rect 248328 291184 248380 291236
rect 250812 291184 250864 291236
rect 262588 291184 262640 291236
rect 271880 291184 271932 291236
rect 269028 291116 269080 291168
rect 272248 291116 272300 291168
rect 336004 291116 336056 291168
rect 336372 291116 336424 291168
rect 367744 291116 367796 291168
rect 262220 290776 262272 290828
rect 262956 290776 263008 290828
rect 172704 290708 172756 290760
rect 219900 290708 219952 290760
rect 227720 290708 227772 290760
rect 240140 290708 240192 290760
rect 261576 290708 261628 290760
rect 197544 290640 197596 290692
rect 256516 290640 256568 290692
rect 256792 290640 256844 290692
rect 194692 290572 194744 290624
rect 254676 290572 254728 290624
rect 193312 290504 193364 290556
rect 253848 290504 253900 290556
rect 179512 290436 179564 290488
rect 240140 290436 240192 290488
rect 244188 290436 244240 290488
rect 272800 290436 272852 290488
rect 221740 290368 221792 290420
rect 240508 290368 240560 290420
rect 168288 290300 168340 290352
rect 220728 290300 220780 290352
rect 221924 290300 221976 290352
rect 259276 290300 259328 290352
rect 219900 290232 219952 290284
rect 260564 290232 260616 290284
rect 202972 290164 203024 290216
rect 262220 290164 262272 290216
rect 176660 290096 176712 290148
rect 236828 290096 236880 290148
rect 199384 290028 199436 290080
rect 259552 290028 259604 290080
rect 169944 289960 169996 290012
rect 230756 289960 230808 290012
rect 256516 289960 256568 290012
rect 257252 289960 257304 290012
rect 197452 289892 197504 289944
rect 258356 289892 258408 289944
rect 182272 289824 182324 289876
rect 243268 289824 243320 289876
rect 220544 289756 220596 289808
rect 223580 289756 223632 289808
rect 180064 289212 180116 289264
rect 234528 289348 234580 289400
rect 235540 289348 235592 289400
rect 184940 289144 184992 289196
rect 244004 289348 244056 289400
rect 245200 289416 245252 289468
rect 245476 289348 245528 289400
rect 185032 289076 185084 289128
rect 183652 288396 183704 288448
rect 323492 289076 323544 289128
rect 328828 289076 328880 289128
rect 389180 289076 389232 289128
rect 538220 289076 538272 289128
rect 306012 288396 306064 288448
rect 307484 288396 307536 288448
rect 268384 287648 268436 287700
rect 325424 287648 325476 287700
rect 194784 286356 194836 286408
rect 220912 286356 220964 286408
rect 183744 286288 183796 286340
rect 268936 286288 268988 286340
rect 321192 286288 321244 286340
rect 220912 286220 220964 286272
rect 219348 285132 219400 285184
rect 220912 285132 220964 285184
rect 193404 284928 193456 284980
rect 220820 285064 220872 285116
rect 269028 284928 269080 284980
rect 325240 284928 325292 284980
rect 196072 283568 196124 283620
rect 220912 283568 220964 283620
rect 271328 283568 271380 283620
rect 290924 283568 290976 283620
rect 271420 282140 271472 282192
rect 292488 282140 292540 282192
rect 196164 280780 196216 280832
rect 219992 280780 220044 280832
rect 271512 280780 271564 280832
rect 292396 280780 292448 280832
rect 182364 279420 182416 279472
rect 220912 279420 220964 279472
rect 271604 279420 271656 279472
rect 292304 279420 292356 279472
rect 323952 277380 324004 277432
rect 327264 277380 327316 277432
rect 531320 277380 531372 277432
rect 185124 276632 185176 276684
rect 220912 276632 220964 276684
rect 322664 276020 322716 276072
rect 322940 276020 322992 276072
rect 516140 276020 516192 276072
rect 187884 273912 187936 273964
rect 220360 273912 220412 273964
rect 321284 273232 321336 273284
rect 321652 273232 321704 273284
rect 495440 273232 495492 273284
rect 3056 266364 3108 266416
rect 14464 266364 14516 266416
rect 325148 266364 325200 266416
rect 325608 266364 325660 266416
rect 543004 266364 543056 266416
rect 317052 264596 317104 264648
rect 317420 264596 317472 264648
rect 314108 263644 314160 263696
rect 314384 263644 314436 263696
rect 414020 263644 414072 263696
rect 317420 263576 317472 263628
rect 445760 263576 445812 263628
rect 312452 262828 312504 262880
rect 347504 262828 347556 262880
rect 389180 262828 389232 262880
rect 318248 262692 318300 262744
rect 318524 262692 318576 262744
rect 318248 262216 318300 262268
rect 452660 262216 452712 262268
rect 295064 260108 295116 260160
rect 322296 260108 322348 260160
rect 310244 259428 310296 259480
rect 360200 259428 360252 259480
rect 316960 258068 317012 258120
rect 441620 258068 441672 258120
rect 269948 257320 270000 257372
rect 313096 257320 313148 257372
rect 391940 257320 391992 257372
rect 319720 256708 319772 256760
rect 470600 256708 470652 256760
rect 315580 255280 315632 255332
rect 315856 255280 315908 255332
rect 427820 255280 427872 255332
rect 268936 254532 268988 254584
rect 290372 254532 290424 254584
rect 311532 253988 311584 254040
rect 364340 253988 364392 254040
rect 3424 253920 3476 253972
rect 323768 253920 323820 253972
rect 527180 253920 527232 253972
rect 200212 253852 200264 253904
rect 216036 253852 216088 253904
rect 275652 253172 275704 253224
rect 321100 253172 321152 253224
rect 316776 253036 316828 253088
rect 317236 253036 317288 253088
rect 310336 252696 310388 252748
rect 349252 252696 349304 252748
rect 317236 252628 317288 252680
rect 448612 252628 448664 252680
rect 323860 252560 323912 252612
rect 324136 252560 324188 252612
rect 523132 252560 523184 252612
rect 268936 251812 268988 251864
rect 290648 251812 290700 251864
rect 214932 251608 214984 251660
rect 215668 251608 215720 251660
rect 315672 251268 315724 251320
rect 315948 251268 316000 251320
rect 423772 251268 423824 251320
rect 321376 251200 321428 251252
rect 491300 251200 491352 251252
rect 271788 250452 271840 250504
rect 317144 250452 317196 250504
rect 438860 250452 438912 250504
rect 323032 249772 323084 249824
rect 324228 249772 324280 249824
rect 534080 249772 534132 249824
rect 307484 249704 307536 249756
rect 308680 249704 308732 249756
rect 314200 249704 314252 249756
rect 314568 249704 314620 249756
rect 292304 249092 292356 249144
rect 316684 249092 316736 249144
rect 171324 249024 171376 249076
rect 215852 249024 215904 249076
rect 273076 249024 273128 249076
rect 323032 249024 323084 249076
rect 312912 248480 312964 248532
rect 382280 248480 382332 248532
rect 314200 248412 314252 248464
rect 407120 248412 407172 248464
rect 168472 247664 168524 247716
rect 217140 247664 217192 247716
rect 282000 247664 282052 247716
rect 307392 247664 307444 247716
rect 314292 247120 314344 247172
rect 409880 247120 409932 247172
rect 318156 247052 318208 247104
rect 318616 247052 318668 247104
rect 459560 247052 459612 247104
rect 168564 246304 168616 246356
rect 217324 246304 217376 246356
rect 269304 246304 269356 246356
rect 292120 246304 292172 246356
rect 310428 245828 310480 245880
rect 353300 245692 353352 245744
rect 310060 245624 310112 245676
rect 310428 245624 310480 245676
rect 316684 245624 316736 245676
rect 317328 245624 317380 245676
rect 434720 245624 434772 245676
rect 577504 245556 577556 245608
rect 579620 245556 579672 245608
rect 287612 244944 287664 244996
rect 312728 244944 312780 244996
rect 167092 244876 167144 244928
rect 218612 244876 218664 244928
rect 285864 244876 285916 244928
rect 314016 244876 314068 244928
rect 312360 244400 312412 244452
rect 312912 244400 312964 244452
rect 385040 244400 385092 244452
rect 318340 244332 318392 244384
rect 456800 244332 456852 244384
rect 321560 244264 321612 244316
rect 322756 244264 322808 244316
rect 507124 244264 507176 244316
rect 288532 243720 288584 243772
rect 270592 243652 270644 243704
rect 288900 243652 288952 243704
rect 313924 243652 313976 243704
rect 273352 243584 273404 243636
rect 315488 243584 315540 243636
rect 191932 243516 191984 243568
rect 218704 243516 218756 243568
rect 274916 243516 274968 243568
rect 321560 243516 321612 243568
rect 210516 243448 210568 243500
rect 213828 243448 213880 243500
rect 320088 242972 320140 243024
rect 471244 242972 471296 243024
rect 321560 242904 321612 242956
rect 322848 242904 322900 242956
rect 520280 242904 520332 242956
rect 313924 242496 313976 242548
rect 315396 242496 315448 242548
rect 268936 242360 268988 242412
rect 271236 242360 271288 242412
rect 284852 242292 284904 242344
rect 309876 242292 309928 242344
rect 271236 242224 271288 242276
rect 277492 242224 277544 242276
rect 321560 242224 321612 242276
rect 173992 242156 174044 242208
rect 214564 242156 214616 242208
rect 269212 242156 269264 242208
rect 276112 242156 276164 242208
rect 324964 242156 325016 242208
rect 268292 242020 268344 242072
rect 271604 242020 271656 242072
rect 274548 241884 274600 241936
rect 275928 241884 275980 241936
rect 160008 241612 160060 241664
rect 204904 241612 204956 241664
rect 221188 241612 221240 241664
rect 269396 241612 269448 241664
rect 271328 241612 271380 241664
rect 157248 241544 157300 241596
rect 206376 241544 206428 241596
rect 207664 241544 207716 241596
rect 222292 241544 222344 241596
rect 269488 241544 269540 241596
rect 271512 241544 271564 241596
rect 274640 241544 274692 241596
rect 275652 241544 275704 241596
rect 320088 241544 320140 241596
rect 481640 241544 481692 241596
rect 154304 241476 154356 241528
rect 209228 241476 209280 241528
rect 215668 241476 215720 241528
rect 14464 241408 14516 241460
rect 198832 241408 198884 241460
rect 199384 241408 199436 241460
rect 219992 241408 220044 241460
rect 220176 241408 220228 241460
rect 221372 241408 221424 241460
rect 216128 241272 216180 241324
rect 221372 241272 221424 241324
rect 214840 241136 214892 241188
rect 219072 241068 219124 241120
rect 220820 241068 220872 241120
rect 213920 241000 213972 241052
rect 220268 240864 220320 240916
rect 218888 240796 218940 240848
rect 189172 240728 189224 240780
rect 220176 240728 220228 240780
rect 220360 240728 220412 240780
rect 206652 240660 206704 240712
rect 222016 240660 222068 240712
rect 219532 240592 219584 240644
rect 215852 240524 215904 240576
rect 216404 240524 216456 240576
rect 213736 240456 213788 240508
rect 214472 240320 214524 240372
rect 216128 240320 216180 240372
rect 206376 240252 206428 240304
rect 213184 240184 213236 240236
rect 214840 240184 214892 240236
rect 216036 240184 216088 240236
rect 219072 240184 219124 240236
rect 219348 240184 219400 240236
rect 217876 240048 217928 240100
rect 219532 240048 219584 240100
rect 222292 240048 222344 240100
rect 217968 239980 218020 240032
rect 222108 239980 222160 240032
rect 215208 239912 215260 239964
rect 222522 239912 222574 239964
rect 222614 239912 222666 239964
rect 222706 239912 222758 239964
rect 210424 239844 210476 239896
rect 221280 239844 221332 239896
rect 221556 239844 221608 239896
rect 222384 239844 222436 239896
rect 216680 239776 216732 239828
rect 223074 239912 223126 239964
rect 223166 239912 223218 239964
rect 222890 239844 222942 239896
rect 163504 239708 163556 239760
rect 222844 239708 222896 239760
rect 198924 239640 198976 239692
rect 218796 239640 218848 239692
rect 218980 239640 219032 239692
rect 222200 239640 222252 239692
rect 223120 239776 223172 239828
rect 186504 239572 186556 239624
rect 220084 239572 220136 239624
rect 221096 239572 221148 239624
rect 223350 239912 223402 239964
rect 223442 239912 223494 239964
rect 223534 239912 223586 239964
rect 223626 239912 223678 239964
rect 223718 239912 223770 239964
rect 223902 239912 223954 239964
rect 223672 239776 223724 239828
rect 223396 239708 223448 239760
rect 223488 239708 223540 239760
rect 223672 239640 223724 239692
rect 159732 239504 159784 239556
rect 205088 239504 205140 239556
rect 205456 239504 205508 239556
rect 215116 239504 215168 239556
rect 224178 239912 224230 239964
rect 224270 239912 224322 239964
rect 224362 239912 224414 239964
rect 224638 239912 224690 239964
rect 224822 239912 224874 239964
rect 224914 239912 224966 239964
rect 225006 239912 225058 239964
rect 224086 239844 224138 239896
rect 224224 239776 224276 239828
rect 224316 239776 224368 239828
rect 224132 239572 224184 239624
rect 224546 239844 224598 239896
rect 224730 239844 224782 239896
rect 224868 239776 224920 239828
rect 224592 239708 224644 239760
rect 224684 239708 224736 239760
rect 224776 239640 224828 239692
rect 224960 239640 225012 239692
rect 225558 239912 225610 239964
rect 225742 239912 225794 239964
rect 225834 239912 225886 239964
rect 226110 239912 226162 239964
rect 226386 239912 226438 239964
rect 226478 239912 226530 239964
rect 226846 239912 226898 239964
rect 227030 239912 227082 239964
rect 227306 239912 227358 239964
rect 225190 239844 225242 239896
rect 225466 239844 225518 239896
rect 225236 239708 225288 239760
rect 224500 239572 224552 239624
rect 158536 239436 158588 239488
rect 220544 239436 220596 239488
rect 221280 239436 221332 239488
rect 221372 239436 221424 239488
rect 223488 239436 223540 239488
rect 224408 239436 224460 239488
rect 3332 239368 3384 239420
rect 198924 239368 198976 239420
rect 212172 239300 212224 239352
rect 223304 239368 223356 239420
rect 224684 239368 224736 239420
rect 225420 239572 225472 239624
rect 225788 239776 225840 239828
rect 225972 239640 226024 239692
rect 226754 239844 226806 239896
rect 226524 239708 226576 239760
rect 226800 239708 226852 239760
rect 226432 239640 226484 239692
rect 227214 239844 227266 239896
rect 227168 239708 227220 239760
rect 227076 239640 227128 239692
rect 227674 239912 227726 239964
rect 227950 239912 228002 239964
rect 228042 239912 228094 239964
rect 228502 239912 228554 239964
rect 227628 239708 227680 239760
rect 227812 239708 227864 239760
rect 227352 239572 227404 239624
rect 227444 239572 227496 239624
rect 228226 239844 228278 239896
rect 228318 239844 228370 239896
rect 227996 239776 228048 239828
rect 228870 239912 228922 239964
rect 229146 239912 229198 239964
rect 229238 239912 229290 239964
rect 229330 239912 229382 239964
rect 229422 239912 229474 239964
rect 229882 239912 229934 239964
rect 228686 239844 228738 239896
rect 229376 239776 229428 239828
rect 228180 239572 228232 239624
rect 228456 239572 228508 239624
rect 228548 239572 228600 239624
rect 228732 239572 228784 239624
rect 228824 239572 228876 239624
rect 229284 239572 229336 239624
rect 229100 239504 229152 239556
rect 229790 239844 229842 239896
rect 229836 239708 229888 239760
rect 230066 239912 230118 239964
rect 230020 239708 230072 239760
rect 229652 239572 229704 239624
rect 225144 239436 225196 239488
rect 225236 239436 225288 239488
rect 225512 239436 225564 239488
rect 226064 239436 226116 239488
rect 226616 239436 226668 239488
rect 229744 239436 229796 239488
rect 270224 241476 270276 241528
rect 273352 241476 273404 241528
rect 321008 241476 321060 241528
rect 321468 241476 321520 241528
rect 488540 241476 488592 241528
rect 271420 241340 271472 241392
rect 271328 241272 271380 241324
rect 273260 241272 273312 241324
rect 273904 241272 273956 241324
rect 230526 239912 230578 239964
rect 230986 239912 231038 239964
rect 231262 239912 231314 239964
rect 230802 239844 230854 239896
rect 230664 239572 230716 239624
rect 230756 239572 230808 239624
rect 231446 239844 231498 239896
rect 231124 239708 231176 239760
rect 231400 239640 231452 239692
rect 231722 239912 231774 239964
rect 232274 239912 232326 239964
rect 232458 239912 232510 239964
rect 232642 239912 232694 239964
rect 232918 239912 232970 239964
rect 233378 239912 233430 239964
rect 233470 239912 233522 239964
rect 233562 239912 233614 239964
rect 233654 239912 233706 239964
rect 233746 239912 233798 239964
rect 233838 239912 233890 239964
rect 233930 239912 233982 239964
rect 234206 239912 234258 239964
rect 234298 239912 234350 239964
rect 234758 239912 234810 239964
rect 234850 239912 234902 239964
rect 231906 239844 231958 239896
rect 231860 239708 231912 239760
rect 232412 239640 232464 239692
rect 232596 239640 232648 239692
rect 233286 239844 233338 239896
rect 233424 239776 233476 239828
rect 233516 239776 233568 239828
rect 234574 239844 234626 239896
rect 233792 239776 233844 239828
rect 233884 239776 233936 239828
rect 234252 239776 234304 239828
rect 233332 239708 233384 239760
rect 233700 239708 233752 239760
rect 234620 239708 234672 239760
rect 233240 239640 233292 239692
rect 231124 239572 231176 239624
rect 231952 239504 232004 239556
rect 233240 239504 233292 239556
rect 233424 239504 233476 239556
rect 232780 239436 232832 239488
rect 232872 239436 232924 239488
rect 233056 239436 233108 239488
rect 233148 239436 233200 239488
rect 234252 239572 234304 239624
rect 234436 239572 234488 239624
rect 234620 239572 234672 239624
rect 235034 239912 235086 239964
rect 235402 239912 235454 239964
rect 235586 239912 235638 239964
rect 235678 239912 235730 239964
rect 236046 239912 236098 239964
rect 234344 239436 234396 239488
rect 234528 239436 234580 239488
rect 235862 239844 235914 239896
rect 235448 239708 235500 239760
rect 235632 239708 235684 239760
rect 235264 239572 235316 239624
rect 236322 239912 236374 239964
rect 236414 239912 236466 239964
rect 236598 239912 236650 239964
rect 236966 239912 237018 239964
rect 237058 239912 237110 239964
rect 235908 239708 235960 239760
rect 236184 239708 236236 239760
rect 236276 239708 236328 239760
rect 235816 239436 235868 239488
rect 217784 239300 217836 239352
rect 224500 239300 224552 239352
rect 225144 239300 225196 239352
rect 225696 239368 225748 239420
rect 227996 239368 228048 239420
rect 230112 239368 230164 239420
rect 230664 239368 230716 239420
rect 236460 239640 236512 239692
rect 236874 239844 236926 239896
rect 236966 239776 237018 239828
rect 236828 239708 236880 239760
rect 236920 239640 236972 239692
rect 236184 239572 236236 239624
rect 237334 239912 237386 239964
rect 237518 239912 237570 239964
rect 237104 239504 237156 239556
rect 237702 239912 237754 239964
rect 237564 239708 237616 239760
rect 237472 239572 237524 239624
rect 237886 239912 237938 239964
rect 238254 239912 238306 239964
rect 238346 239912 238398 239964
rect 238438 239912 238490 239964
rect 271052 241136 271104 241188
rect 268108 240864 268160 240916
rect 283564 241204 283616 241256
rect 308588 241204 308640 241256
rect 282276 241136 282328 241188
rect 307300 241136 307352 241188
rect 271512 241068 271564 241120
rect 303160 241068 303212 241120
rect 272064 241000 272116 241052
rect 320088 241000 320140 241052
rect 271696 240932 271748 240984
rect 321008 240932 321060 240984
rect 271420 240864 271472 240916
rect 294972 240864 295024 240916
rect 271328 240796 271380 240848
rect 299112 240796 299164 240848
rect 239082 239912 239134 239964
rect 238070 239844 238122 239896
rect 238530 239844 238582 239896
rect 238622 239844 238674 239896
rect 238806 239844 238858 239896
rect 238898 239844 238950 239896
rect 238300 239776 238352 239828
rect 238484 239708 238536 239760
rect 238576 239708 238628 239760
rect 238760 239708 238812 239760
rect 238116 239640 238168 239692
rect 238208 239572 238260 239624
rect 237932 239504 237984 239556
rect 238024 239436 238076 239488
rect 238760 239436 238812 239488
rect 236736 239368 236788 239420
rect 237012 239368 237064 239420
rect 238852 239368 238904 239420
rect 239542 239912 239594 239964
rect 239910 239912 239962 239964
rect 240094 239912 240146 239964
rect 240370 239912 240422 239964
rect 240830 239912 240882 239964
rect 240922 239912 240974 239964
rect 241014 239912 241066 239964
rect 239726 239844 239778 239896
rect 239588 239708 239640 239760
rect 239496 239436 239548 239488
rect 239864 239572 239916 239624
rect 240554 239844 240606 239896
rect 240140 239572 240192 239624
rect 240508 239640 240560 239692
rect 240692 239572 240744 239624
rect 240876 239504 240928 239556
rect 240784 239436 240836 239488
rect 241198 239912 241250 239964
rect 241474 239912 241526 239964
rect 241934 239912 241986 239964
rect 242026 239912 242078 239964
rect 242394 239912 242446 239964
rect 242762 239912 242814 239964
rect 242854 239912 242906 239964
rect 242946 239912 242998 239964
rect 243130 239912 243182 239964
rect 243314 239912 243366 239964
rect 243406 239912 243458 239964
rect 243682 239912 243734 239964
rect 243866 239912 243918 239964
rect 241060 239640 241112 239692
rect 241290 239844 241342 239896
rect 241842 239844 241894 239896
rect 241520 239640 241572 239692
rect 241888 239708 241940 239760
rect 242072 239708 242124 239760
rect 241980 239640 242032 239692
rect 241244 239572 241296 239624
rect 239404 239368 239456 239420
rect 241336 239436 241388 239488
rect 241796 239436 241848 239488
rect 242716 239640 242768 239692
rect 242808 239640 242860 239692
rect 243038 239844 243090 239896
rect 242992 239640 243044 239692
rect 243084 239640 243136 239692
rect 243268 239640 243320 239692
rect 243452 239572 243504 239624
rect 243360 239504 243412 239556
rect 243820 239708 243872 239760
rect 271052 240728 271104 240780
rect 292764 240728 292816 240780
rect 244418 239912 244470 239964
rect 244694 239912 244746 239964
rect 244970 239912 245022 239964
rect 244142 239844 244194 239896
rect 244234 239844 244286 239896
rect 244096 239708 244148 239760
rect 244510 239844 244562 239896
rect 244004 239640 244056 239692
rect 244188 239640 244240 239692
rect 244556 239640 244608 239692
rect 244464 239572 244516 239624
rect 244740 239708 244792 239760
rect 244004 239504 244056 239556
rect 244372 239504 244424 239556
rect 244372 239368 244424 239420
rect 245016 239708 245068 239760
rect 244924 239572 244976 239624
rect 245338 239912 245390 239964
rect 245522 239912 245574 239964
rect 245614 239912 245666 239964
rect 245982 239912 246034 239964
rect 246534 239912 246586 239964
rect 246626 239912 246678 239964
rect 246810 239912 246862 239964
rect 246994 239912 247046 239964
rect 247086 239912 247138 239964
rect 247270 239912 247322 239964
rect 247362 239912 247414 239964
rect 245706 239844 245758 239896
rect 245200 239572 245252 239624
rect 245476 239572 245528 239624
rect 245568 239572 245620 239624
rect 245016 239368 245068 239420
rect 246074 239844 246126 239896
rect 246166 239844 246218 239896
rect 246258 239844 246310 239896
rect 246350 239844 246402 239896
rect 246028 239708 246080 239760
rect 246120 239708 246172 239760
rect 246304 239640 246356 239692
rect 246672 239708 246724 239760
rect 246856 239708 246908 239760
rect 247546 239844 247598 239896
rect 247132 239708 247184 239760
rect 247224 239708 247276 239760
rect 246488 239640 246540 239692
rect 247040 239640 247092 239692
rect 247500 239572 247552 239624
rect 246580 239504 246632 239556
rect 247316 239436 247368 239488
rect 247684 239436 247736 239488
rect 246304 239368 246356 239420
rect 247040 239368 247092 239420
rect 247408 239368 247460 239420
rect 248006 239912 248058 239964
rect 247868 239572 247920 239624
rect 248466 239912 248518 239964
rect 248650 239912 248702 239964
rect 248742 239912 248794 239964
rect 248834 239912 248886 239964
rect 248926 239912 248978 239964
rect 249018 239912 249070 239964
rect 249202 239912 249254 239964
rect 249386 239912 249438 239964
rect 249478 239912 249530 239964
rect 249938 239912 249990 239964
rect 250122 239912 250174 239964
rect 250306 239912 250358 239964
rect 250490 239912 250542 239964
rect 250582 239912 250634 239964
rect 250766 239912 250818 239964
rect 248512 239708 248564 239760
rect 248696 239708 248748 239760
rect 248788 239708 248840 239760
rect 248880 239640 248932 239692
rect 249294 239844 249346 239896
rect 249156 239708 249208 239760
rect 249248 239708 249300 239760
rect 248880 239504 248932 239556
rect 249340 239640 249392 239692
rect 249662 239844 249714 239896
rect 249846 239844 249898 239896
rect 249616 239708 249668 239760
rect 249708 239572 249760 239624
rect 249800 239572 249852 239624
rect 250950 239912 251002 239964
rect 250260 239708 250312 239760
rect 250444 239708 250496 239760
rect 250628 239708 250680 239760
rect 250812 239708 250864 239760
rect 250536 239640 250588 239692
rect 251134 239912 251186 239964
rect 251226 239844 251278 239896
rect 251502 239844 251554 239896
rect 251594 239844 251646 239896
rect 251180 239640 251232 239692
rect 251088 239572 251140 239624
rect 251456 239572 251508 239624
rect 251870 239912 251922 239964
rect 251640 239572 251692 239624
rect 251824 239572 251876 239624
rect 249892 239504 249944 239556
rect 250076 239504 250128 239556
rect 251364 239504 251416 239556
rect 252514 239912 252566 239964
rect 252974 239912 253026 239964
rect 252146 239844 252198 239896
rect 252330 239844 252382 239896
rect 252008 239572 252060 239624
rect 252376 239708 252428 239760
rect 252100 239504 252152 239556
rect 252698 239844 252750 239896
rect 253158 239844 253210 239896
rect 253434 239912 253486 239964
rect 253526 239912 253578 239964
rect 253618 239912 253670 239964
rect 253894 239912 253946 239964
rect 253986 239912 254038 239964
rect 254262 239912 254314 239964
rect 254446 239912 254498 239964
rect 254814 239912 254866 239964
rect 252652 239640 252704 239692
rect 253020 239640 253072 239692
rect 253204 239640 253256 239692
rect 253296 239640 253348 239692
rect 253664 239640 253716 239692
rect 253756 239640 253808 239692
rect 254308 239708 254360 239760
rect 254630 239844 254682 239896
rect 253572 239572 253624 239624
rect 253940 239572 253992 239624
rect 252836 239504 252888 239556
rect 254216 239572 254268 239624
rect 254998 239912 255050 239964
rect 255090 239912 255142 239964
rect 254768 239640 254820 239692
rect 255274 239912 255326 239964
rect 255458 239912 255510 239964
rect 256010 239912 256062 239964
rect 256102 239912 256154 239964
rect 256378 239912 256430 239964
rect 254952 239708 255004 239760
rect 255136 239708 255188 239760
rect 255734 239844 255786 239896
rect 255826 239844 255878 239896
rect 255504 239708 255556 239760
rect 255228 239572 255280 239624
rect 255872 239640 255924 239692
rect 255780 239572 255832 239624
rect 255964 239572 256016 239624
rect 256286 239844 256338 239896
rect 256240 239640 256292 239692
rect 256332 239640 256384 239692
rect 256562 239912 256614 239964
rect 256654 239912 256706 239964
rect 256148 239572 256200 239624
rect 254492 239504 254544 239556
rect 255136 239504 255188 239556
rect 255412 239504 255464 239556
rect 255596 239504 255648 239556
rect 256516 239504 256568 239556
rect 256930 239912 256982 239964
rect 257114 239912 257166 239964
rect 257298 239912 257350 239964
rect 257482 239912 257534 239964
rect 257574 239912 257626 239964
rect 257758 239912 257810 239964
rect 257850 239912 257902 239964
rect 258402 239912 258454 239964
rect 258494 239912 258546 239964
rect 258678 239912 258730 239964
rect 258862 239912 258914 239964
rect 259138 239912 259190 239964
rect 257206 239844 257258 239896
rect 257160 239708 257212 239760
rect 257620 239640 257672 239692
rect 257712 239640 257764 239692
rect 256884 239572 256936 239624
rect 257528 239572 257580 239624
rect 258218 239844 258270 239896
rect 258448 239776 258500 239828
rect 258356 239708 258408 239760
rect 258540 239640 258592 239692
rect 258264 239572 258316 239624
rect 257068 239504 257120 239556
rect 257804 239504 257856 239556
rect 257988 239504 258040 239556
rect 258816 239708 258868 239760
rect 259322 239912 259374 239964
rect 259690 239912 259742 239964
rect 260058 239912 260110 239964
rect 260426 239912 260478 239964
rect 260518 239912 260570 239964
rect 260610 239912 260662 239964
rect 260702 239912 260754 239964
rect 259184 239708 259236 239760
rect 259460 239640 259512 239692
rect 259092 239572 259144 239624
rect 259644 239572 259696 239624
rect 259920 239572 259972 239624
rect 260472 239776 260524 239828
rect 260564 239776 260616 239828
rect 260656 239708 260708 239760
rect 278136 240524 278188 240576
rect 267924 240456 267976 240508
rect 271236 240320 271288 240372
rect 267740 240252 267792 240304
rect 268108 240184 268160 240236
rect 273076 240184 273128 240236
rect 269212 240116 269264 240168
rect 276020 240116 276072 240168
rect 267924 240048 267976 240100
rect 260978 239912 261030 239964
rect 261438 239912 261490 239964
rect 260840 239640 260892 239692
rect 260196 239572 260248 239624
rect 260840 239504 260892 239556
rect 261254 239844 261306 239896
rect 261346 239844 261398 239896
rect 261300 239640 261352 239692
rect 261898 239912 261950 239964
rect 261990 239912 262042 239964
rect 262082 239912 262134 239964
rect 262174 239912 262226 239964
rect 261622 239844 261674 239896
rect 261714 239844 261766 239896
rect 261484 239708 261536 239760
rect 261576 239708 261628 239760
rect 261668 239708 261720 239760
rect 261944 239776 261996 239828
rect 262128 239776 262180 239828
rect 262036 239708 262088 239760
rect 262358 239912 262410 239964
rect 262450 239912 262502 239964
rect 262818 239912 262870 239964
rect 262910 239912 262962 239964
rect 263002 239912 263054 239964
rect 263278 239912 263330 239964
rect 263370 239912 263422 239964
rect 263830 239912 263882 239964
rect 264014 239912 264066 239964
rect 262220 239640 262272 239692
rect 262404 239776 262456 239828
rect 263186 239844 263238 239896
rect 262956 239776 263008 239828
rect 263048 239708 263100 239760
rect 262864 239640 262916 239692
rect 263232 239640 263284 239692
rect 270500 239980 270552 240032
rect 264290 239912 264342 239964
rect 264382 239912 264434 239964
rect 264658 239912 264710 239964
rect 264336 239776 264388 239828
rect 264520 239708 264572 239760
rect 264842 239844 264894 239896
rect 263508 239640 263560 239692
rect 263876 239640 263928 239692
rect 264428 239640 264480 239692
rect 264796 239640 264848 239692
rect 265026 239912 265078 239964
rect 265578 239912 265630 239964
rect 265762 239912 265814 239964
rect 266130 239912 266182 239964
rect 266314 239912 266366 239964
rect 266682 239912 266734 239964
rect 266958 239912 267010 239964
rect 267050 239912 267102 239964
rect 268016 239912 268068 239964
rect 268476 239912 268528 239964
rect 269212 239912 269264 239964
rect 265118 239844 265170 239896
rect 265210 239844 265262 239896
rect 265302 239844 265354 239896
rect 265072 239640 265124 239692
rect 263140 239572 263192 239624
rect 264888 239572 264940 239624
rect 261392 239504 261444 239556
rect 262680 239504 262732 239556
rect 265946 239844 265998 239896
rect 266406 239844 266458 239896
rect 266498 239844 266550 239896
rect 265900 239708 265952 239760
rect 265992 239708 266044 239760
rect 266268 239708 266320 239760
rect 266360 239708 266412 239760
rect 267142 239844 267194 239896
rect 267832 239844 267884 239896
rect 267004 239776 267056 239828
rect 266544 239708 266596 239760
rect 266636 239708 266688 239760
rect 266820 239708 266872 239760
rect 270960 239708 271012 239760
rect 266912 239640 266964 239692
rect 269120 239640 269172 239692
rect 266176 239572 266228 239624
rect 267372 239572 267424 239624
rect 269304 239572 269356 239624
rect 278412 239708 278464 239760
rect 299296 239708 299348 239760
rect 278136 239640 278188 239692
rect 292212 239640 292264 239692
rect 278412 239572 278464 239624
rect 265808 239504 265860 239556
rect 266084 239504 266136 239556
rect 268200 239504 268252 239556
rect 286968 239504 287020 239556
rect 311440 239504 311492 239556
rect 248328 239436 248380 239488
rect 260748 239436 260800 239488
rect 263600 239436 263652 239488
rect 264980 239436 265032 239488
rect 265256 239436 265308 239488
rect 266636 239436 266688 239488
rect 273260 239436 273312 239488
rect 278136 239436 278188 239488
rect 305828 239436 305880 239488
rect 249064 239368 249116 239420
rect 285312 239368 285364 239420
rect 302148 239368 302200 239420
rect 348792 239368 348844 239420
rect 558920 239368 558972 239420
rect 152924 239232 152976 239284
rect 154120 239164 154172 239216
rect 224224 239164 224276 239216
rect 224408 239164 224460 239216
rect 224960 239232 225012 239284
rect 225236 239232 225288 239284
rect 227444 239300 227496 239352
rect 232228 239300 232280 239352
rect 280712 239300 280764 239352
rect 226616 239232 226668 239284
rect 227168 239232 227220 239284
rect 228548 239232 228600 239284
rect 229284 239232 229336 239284
rect 231308 239232 231360 239284
rect 231676 239232 231728 239284
rect 248052 239232 248104 239284
rect 250536 239232 250588 239284
rect 282092 239232 282144 239284
rect 213000 239028 213052 239080
rect 216220 239028 216272 239080
rect 224684 239096 224736 239148
rect 225880 239096 225932 239148
rect 227996 239164 228048 239216
rect 282920 239164 282972 239216
rect 228824 239096 228876 239148
rect 231676 239096 231728 239148
rect 233056 239096 233108 239148
rect 234712 239028 234764 239080
rect 234988 239096 235040 239148
rect 248328 239096 248380 239148
rect 248512 239096 248564 239148
rect 292672 239096 292724 239148
rect 237012 239028 237064 239080
rect 237840 239028 237892 239080
rect 297824 239028 297876 239080
rect 215852 238960 215904 239012
rect 225144 238960 225196 239012
rect 226064 238960 226116 239012
rect 228088 238960 228140 239012
rect 229744 238960 229796 239012
rect 220268 238892 220320 238944
rect 230664 238892 230716 238944
rect 230848 238892 230900 238944
rect 231492 238892 231544 238944
rect 232412 238892 232464 238944
rect 234988 238892 235040 238944
rect 237564 238960 237616 239012
rect 297640 238960 297692 239012
rect 238760 238892 238812 238944
rect 240600 238892 240652 238944
rect 217600 238824 217652 238876
rect 220728 238824 220780 238876
rect 222108 238824 222160 238876
rect 240232 238824 240284 238876
rect 220360 238756 220412 238808
rect 233056 238756 233108 238808
rect 233240 238756 233292 238808
rect 248512 238892 248564 238944
rect 249248 238892 249300 238944
rect 305920 238892 305972 238944
rect 246488 238824 246540 238876
rect 262772 238824 262824 238876
rect 245292 238756 245344 238808
rect 245844 238756 245896 238808
rect 247316 238756 247368 238808
rect 262956 238756 263008 238808
rect 209228 238688 209280 238740
rect 223764 238688 223816 238740
rect 224224 238688 224276 238740
rect 226708 238688 226760 238740
rect 230020 238688 230072 238740
rect 222844 238620 222896 238672
rect 232412 238620 232464 238672
rect 233516 238688 233568 238740
rect 233792 238688 233844 238740
rect 236184 238688 236236 238740
rect 234988 238620 235040 238672
rect 240968 238688 241020 238740
rect 245200 238688 245252 238740
rect 249248 238688 249300 238740
rect 250904 238688 250956 238740
rect 251180 238688 251232 238740
rect 257160 238688 257212 238740
rect 257896 238688 257948 238740
rect 260472 238688 260524 238740
rect 269580 238824 269632 238876
rect 296628 238824 296680 238876
rect 506480 238824 506532 238876
rect 264980 238756 265032 238808
rect 278136 238756 278188 238808
rect 296536 238756 296588 238808
rect 540980 238756 541032 238808
rect 264428 238688 264480 238740
rect 269212 238688 269264 238740
rect 240232 238620 240284 238672
rect 249064 238620 249116 238672
rect 249432 238620 249484 238672
rect 251456 238620 251508 238672
rect 251824 238620 251876 238672
rect 258816 238620 258868 238672
rect 207756 238552 207808 238604
rect 231860 238552 231912 238604
rect 232780 238552 232832 238604
rect 239588 238552 239640 238604
rect 250168 238552 250220 238604
rect 251272 238552 251324 238604
rect 252008 238552 252060 238604
rect 270960 238620 271012 238672
rect 271052 238620 271104 238672
rect 312452 238620 312504 238672
rect 261300 238552 261352 238604
rect 264428 238552 264480 238604
rect 265992 238552 266044 238604
rect 270868 238552 270920 238604
rect 210332 238484 210384 238536
rect 226524 238484 226576 238536
rect 228824 238484 228876 238536
rect 231216 238484 231268 238536
rect 232136 238484 232188 238536
rect 233056 238484 233108 238536
rect 233240 238484 233292 238536
rect 268568 238484 268620 238536
rect 209320 238416 209372 238468
rect 222568 238416 222620 238468
rect 222844 238416 222896 238468
rect 230204 238416 230256 238468
rect 230664 238416 230716 238468
rect 267280 238416 267332 238468
rect 269304 238416 269356 238468
rect 271512 238416 271564 238468
rect 192484 238348 192536 238400
rect 223580 238348 223632 238400
rect 225328 238348 225380 238400
rect 225788 238348 225840 238400
rect 226524 238348 226576 238400
rect 227352 238348 227404 238400
rect 228456 238348 228508 238400
rect 229100 238348 229152 238400
rect 231952 238348 232004 238400
rect 237104 238348 237156 238400
rect 239220 238348 239272 238400
rect 239588 238348 239640 238400
rect 191656 238280 191708 238332
rect 222752 238280 222804 238332
rect 194324 238212 194376 238264
rect 225420 238280 225472 238332
rect 227444 238280 227496 238332
rect 229836 238280 229888 238332
rect 230388 238280 230440 238332
rect 233240 238280 233292 238332
rect 233424 238280 233476 238332
rect 270776 238348 270828 238400
rect 225328 238212 225380 238264
rect 227904 238212 227956 238264
rect 229192 238212 229244 238264
rect 229652 238212 229704 238264
rect 231492 238212 231544 238264
rect 268844 238280 268896 238332
rect 182916 238144 182968 238196
rect 218980 238144 219032 238196
rect 222568 238144 222620 238196
rect 225696 238144 225748 238196
rect 225880 238144 225932 238196
rect 226984 238144 227036 238196
rect 227812 238144 227864 238196
rect 231952 238144 232004 238196
rect 233056 238144 233108 238196
rect 259828 238144 259880 238196
rect 263876 238144 263928 238196
rect 161296 238076 161348 238128
rect 215944 238076 215996 238128
rect 216588 238076 216640 238128
rect 225604 238076 225656 238128
rect 231676 238076 231728 238128
rect 231768 238076 231820 238128
rect 247684 238076 247736 238128
rect 267372 238212 267424 238264
rect 267740 238212 267792 238264
rect 268384 238212 268436 238264
rect 268476 238144 268528 238196
rect 319628 238144 319680 238196
rect 265808 238076 265860 238128
rect 322940 238076 322992 238128
rect 161204 238008 161256 238060
rect 238484 238008 238536 238060
rect 239220 238008 239272 238060
rect 239404 238008 239456 238060
rect 242900 238008 242952 238060
rect 245016 238008 245068 238060
rect 246580 238008 246632 238060
rect 268016 238008 268068 238060
rect 335544 238008 335596 238060
rect 221464 237940 221516 237992
rect 232320 237940 232372 237992
rect 236276 237940 236328 237992
rect 236920 237940 236972 237992
rect 246396 237940 246448 237992
rect 247132 237940 247184 237992
rect 262036 237940 262088 237992
rect 266636 237940 266688 237992
rect 266820 237940 266872 237992
rect 267556 237940 267608 237992
rect 268568 237940 268620 237992
rect 268752 237940 268804 237992
rect 304724 237940 304776 237992
rect 225144 237872 225196 237924
rect 238944 237872 238996 237924
rect 239864 237872 239916 237924
rect 241612 237872 241664 237924
rect 243728 237872 243780 237924
rect 258908 237872 258960 237924
rect 259736 237872 259788 237924
rect 269120 237872 269172 237924
rect 270316 237872 270368 237924
rect 275744 237872 275796 237924
rect 216588 237804 216640 237856
rect 229100 237804 229152 237856
rect 216312 237736 216364 237788
rect 235724 237804 235776 237856
rect 236276 237804 236328 237856
rect 236460 237804 236512 237856
rect 254308 237804 254360 237856
rect 260472 237804 260524 237856
rect 263876 237804 263928 237856
rect 270592 237804 270644 237856
rect 272064 237804 272116 237856
rect 229928 237736 229980 237788
rect 233424 237736 233476 237788
rect 253940 237736 253992 237788
rect 271236 237736 271288 237788
rect 231860 237668 231912 237720
rect 224500 237600 224552 237652
rect 235172 237600 235224 237652
rect 257988 237668 258040 237720
rect 259920 237668 259972 237720
rect 264060 237668 264112 237720
rect 270316 237668 270368 237720
rect 271604 237600 271656 237652
rect 162308 237396 162360 237448
rect 231584 237532 231636 237584
rect 231676 237532 231728 237584
rect 269488 237532 269540 237584
rect 230572 237464 230624 237516
rect 269396 237464 269448 237516
rect 229376 237396 229428 237448
rect 229560 237396 229612 237448
rect 229928 237396 229980 237448
rect 231308 237396 231360 237448
rect 231492 237396 231544 237448
rect 231584 237396 231636 237448
rect 236920 237396 236972 237448
rect 252284 237396 252336 237448
rect 252652 237396 252704 237448
rect 271052 237396 271104 237448
rect 281540 237396 281592 237448
rect 284484 237396 284536 237448
rect 231952 237328 232004 237380
rect 232228 237328 232280 237380
rect 267556 237328 267608 237380
rect 267832 237328 267884 237380
rect 269120 237328 269172 237380
rect 270408 237328 270460 237380
rect 281356 237328 281408 237380
rect 213460 237260 213512 237312
rect 221648 237260 221700 237312
rect 255688 237260 255740 237312
rect 261484 237260 261536 237312
rect 274640 237260 274692 237312
rect 276296 237260 276348 237312
rect 277124 237260 277176 237312
rect 277400 237260 277452 237312
rect 278504 237260 278556 237312
rect 205548 237192 205600 237244
rect 224316 237192 224368 237244
rect 234896 237192 234948 237244
rect 253296 237192 253348 237244
rect 254400 237192 254452 237244
rect 294788 237192 294840 237244
rect 239864 237124 239916 237176
rect 240048 237124 240100 237176
rect 252652 237124 252704 237176
rect 253664 237124 253716 237176
rect 234804 237056 234856 237108
rect 235632 237056 235684 237108
rect 237288 237056 237340 237108
rect 241152 237056 241204 237108
rect 245660 237056 245712 237108
rect 253296 237056 253348 237108
rect 214840 236920 214892 236972
rect 235908 236988 235960 237040
rect 239864 236988 239916 237040
rect 240692 236988 240744 237040
rect 240784 236988 240836 237040
rect 241060 236988 241112 237040
rect 246580 236988 246632 237040
rect 254400 236988 254452 237040
rect 254860 236988 254912 237040
rect 286600 237124 286652 237176
rect 232504 236920 232556 236972
rect 232688 236920 232740 236972
rect 235632 236920 235684 236972
rect 252284 236920 252336 236972
rect 253296 236920 253348 236972
rect 277032 237056 277084 237108
rect 259552 236988 259604 237040
rect 260288 236988 260340 237040
rect 260472 236988 260524 237040
rect 285864 236988 285916 237040
rect 258908 236920 258960 236972
rect 268384 236920 268436 236972
rect 212172 236852 212224 236904
rect 238116 236852 238168 236904
rect 240692 236852 240744 236904
rect 241428 236852 241480 236904
rect 244556 236852 244608 236904
rect 267832 236852 267884 236904
rect 287704 236852 287756 236904
rect 161388 236784 161440 236836
rect 213276 236784 213328 236836
rect 214932 236784 214984 236836
rect 253020 236784 253072 236836
rect 255872 236784 255924 236836
rect 276020 236784 276072 236836
rect 296076 236784 296128 236836
rect 150348 236716 150400 236768
rect 215116 236716 215168 236768
rect 221556 236716 221608 236768
rect 244096 236716 244148 236768
rect 278780 236716 278832 236768
rect 332876 236716 332928 236768
rect 159824 236648 159876 236700
rect 231952 236648 232004 236700
rect 242532 236648 242584 236700
rect 243084 236648 243136 236700
rect 245200 236648 245252 236700
rect 299664 236648 299716 236700
rect 307668 236648 307720 236700
rect 321560 236648 321612 236700
rect 213368 236580 213420 236632
rect 223672 236580 223724 236632
rect 241336 236580 241388 236632
rect 242992 236580 243044 236632
rect 244832 236580 244884 236632
rect 245292 236580 245344 236632
rect 247224 236580 247276 236632
rect 247684 236580 247736 236632
rect 248236 236580 248288 236632
rect 248972 236580 249024 236632
rect 266360 236580 266412 236632
rect 330024 236580 330076 236632
rect 217600 236512 217652 236564
rect 219992 236512 220044 236564
rect 254584 236512 254636 236564
rect 255780 236512 255832 236564
rect 256424 236512 256476 236564
rect 259184 236512 259236 236564
rect 276296 236512 276348 236564
rect 244832 236444 244884 236496
rect 245476 236444 245528 236496
rect 253940 236444 253992 236496
rect 255044 236444 255096 236496
rect 268384 236444 268436 236496
rect 277400 236444 277452 236496
rect 244556 236376 244608 236428
rect 249616 236376 249668 236428
rect 310152 236376 310204 236428
rect 252560 236308 252612 236360
rect 261208 236308 261260 236360
rect 263508 236308 263560 236360
rect 270776 236308 270828 236360
rect 233976 236104 234028 236156
rect 244924 236104 244976 236156
rect 245660 236104 245712 236156
rect 237472 236036 237524 236088
rect 238668 236036 238720 236088
rect 242072 236036 242124 236088
rect 212356 235968 212408 236020
rect 214840 235968 214892 236020
rect 217508 235968 217560 236020
rect 246304 235968 246356 236020
rect 246948 235968 247000 236020
rect 247132 235968 247184 236020
rect 248420 235968 248472 236020
rect 214012 235900 214064 235952
rect 224408 235900 224460 235952
rect 224868 235900 224920 235952
rect 236920 235900 236972 235952
rect 242072 235900 242124 235952
rect 207020 235832 207072 235884
rect 208032 235832 208084 235884
rect 224224 235832 224276 235884
rect 242164 235832 242216 235884
rect 243728 235832 243780 235884
rect 256976 236036 257028 236088
rect 267188 236036 267240 236088
rect 256056 235968 256108 236020
rect 261484 235968 261536 236020
rect 265256 235968 265308 236020
rect 265992 235968 266044 236020
rect 266176 235968 266228 236020
rect 269028 235968 269080 236020
rect 272708 235968 272760 236020
rect 299664 235968 299716 236020
rect 300400 235968 300452 236020
rect 288348 235900 288400 235952
rect 329932 235900 329984 235952
rect 276940 235832 276992 235884
rect 278780 235832 278832 235884
rect 301964 235832 302016 235884
rect 242808 235764 242860 235816
rect 244924 235764 244976 235816
rect 250352 235764 250404 235816
rect 284852 235764 284904 235816
rect 210608 235696 210660 235748
rect 245200 235696 245252 235748
rect 263324 235696 263376 235748
rect 268936 235696 268988 235748
rect 269028 235696 269080 235748
rect 277860 235696 277912 235748
rect 211620 235628 211672 235680
rect 244556 235628 244608 235680
rect 266176 235628 266228 235680
rect 267464 235628 267516 235680
rect 209228 235560 209280 235612
rect 239404 235560 239456 235612
rect 252284 235560 252336 235612
rect 252928 235560 252980 235612
rect 260196 235560 260248 235612
rect 270224 235560 270276 235612
rect 281264 235560 281316 235612
rect 214840 235492 214892 235544
rect 244740 235492 244792 235544
rect 285680 235492 285732 235544
rect 159640 235424 159692 235476
rect 207020 235424 207072 235476
rect 210700 235424 210752 235476
rect 256424 235424 256476 235476
rect 264704 235424 264756 235476
rect 282460 235424 282512 235476
rect 331496 235424 331548 235476
rect 161020 235356 161072 235408
rect 216680 235356 216732 235408
rect 155776 235288 155828 235340
rect 216496 235288 216548 235340
rect 225972 235356 226024 235408
rect 229744 235356 229796 235408
rect 230388 235356 230440 235408
rect 245476 235356 245528 235408
rect 246488 235356 246540 235408
rect 260564 235356 260616 235408
rect 273904 235356 273956 235408
rect 328644 235356 328696 235408
rect 220176 235288 220228 235340
rect 237104 235288 237156 235340
rect 243452 235288 243504 235340
rect 243912 235288 243964 235340
rect 261668 235288 261720 235340
rect 267924 235288 267976 235340
rect 268936 235288 268988 235340
rect 271236 235288 271288 235340
rect 329104 235288 329156 235340
rect 158444 235220 158496 235272
rect 233148 235220 233200 235272
rect 234712 235220 234764 235272
rect 235724 235220 235776 235272
rect 207020 235152 207072 235204
rect 207848 235152 207900 235204
rect 227720 235152 227772 235204
rect 236644 235152 236696 235204
rect 258356 235220 258408 235272
rect 259460 235220 259512 235272
rect 260932 235220 260984 235272
rect 269120 235220 269172 235272
rect 331588 235220 331640 235272
rect 254032 235152 254084 235204
rect 254676 235152 254728 235204
rect 257620 235152 257672 235204
rect 266452 235152 266504 235204
rect 239404 235084 239456 235136
rect 250812 235084 250864 235136
rect 263876 235084 263928 235136
rect 266360 235084 266412 235136
rect 267004 235084 267056 235136
rect 222568 235016 222620 235068
rect 226156 235016 226208 235068
rect 256884 235016 256936 235068
rect 257252 235016 257304 235068
rect 259460 235016 259512 235068
rect 270132 235016 270184 235068
rect 244648 234948 244700 235000
rect 245200 234948 245252 235000
rect 245660 234948 245712 235000
rect 289084 234948 289136 235000
rect 237196 234880 237248 234932
rect 240416 234880 240468 234932
rect 240876 234880 240928 234932
rect 241060 234880 241112 234932
rect 262312 234880 262364 234932
rect 269028 234880 269080 234932
rect 251916 234812 251968 234864
rect 265808 234812 265860 234864
rect 232872 234744 232924 234796
rect 238300 234744 238352 234796
rect 263048 234744 263100 234796
rect 270132 234744 270184 234796
rect 215944 234608 215996 234660
rect 245476 234676 245528 234728
rect 258356 234676 258408 234728
rect 259276 234676 259328 234728
rect 260840 234676 260892 234728
rect 261576 234676 261628 234728
rect 263508 234676 263560 234728
rect 263784 234676 263836 234728
rect 265164 234676 265216 234728
rect 265716 234676 265768 234728
rect 284300 234676 284352 234728
rect 284852 234676 284904 234728
rect 247316 234608 247368 234660
rect 291844 234608 291896 234660
rect 212540 234540 212592 234592
rect 243360 234540 243412 234592
rect 243544 234540 243596 234592
rect 303068 234540 303120 234592
rect 211896 234472 211948 234524
rect 246672 234472 246724 234524
rect 247040 234472 247092 234524
rect 305644 234472 305696 234524
rect 237656 234404 237708 234456
rect 286876 234404 286928 234456
rect 223764 234336 223816 234388
rect 226064 234336 226116 234388
rect 228180 234336 228232 234388
rect 228456 234336 228508 234388
rect 237012 234336 237064 234388
rect 279884 234336 279936 234388
rect 285680 234336 285732 234388
rect 304632 234336 304684 234388
rect 249800 234268 249852 234320
rect 293224 234268 293276 234320
rect 237564 234200 237616 234252
rect 238300 234200 238352 234252
rect 239588 234200 239640 234252
rect 282736 234200 282788 234252
rect 210792 234132 210844 234184
rect 212540 234132 212592 234184
rect 219992 234132 220044 234184
rect 153108 234064 153160 234116
rect 211988 234064 212040 234116
rect 237104 234132 237156 234184
rect 240784 234132 240836 234184
rect 281908 234132 281960 234184
rect 238208 234064 238260 234116
rect 277768 234064 277820 234116
rect 161112 233996 161164 234048
rect 234896 233996 234948 234048
rect 236276 233996 236328 234048
rect 276848 233996 276900 234048
rect 156972 233928 157024 233980
rect 224868 233928 224920 233980
rect 240600 233928 240652 233980
rect 279700 233928 279752 233980
rect 151636 233860 151688 233912
rect 231216 233860 231268 233912
rect 216128 233588 216180 233640
rect 217784 233588 217836 233640
rect 241428 233588 241480 233640
rect 273536 233860 273588 233912
rect 243544 233792 243596 233844
rect 244188 233792 244240 233844
rect 246120 233792 246172 233844
rect 271788 233792 271840 233844
rect 272524 233792 272576 233844
rect 272892 233792 272944 233844
rect 244924 233724 244976 233776
rect 274364 233724 274416 233776
rect 247960 233520 248012 233572
rect 272524 233656 272576 233708
rect 256700 233588 256752 233640
rect 257436 233588 257488 233640
rect 260012 233588 260064 233640
rect 260472 233588 260524 233640
rect 271788 233588 271840 233640
rect 274824 233588 274876 233640
rect 263692 233520 263744 233572
rect 264520 233520 264572 233572
rect 219532 233316 219584 233368
rect 223856 233316 223908 233368
rect 248328 233316 248380 233368
rect 249800 233316 249852 233368
rect 217416 233248 217468 233300
rect 231860 233248 231912 233300
rect 258264 233248 258316 233300
rect 259368 233248 259420 233300
rect 278044 233248 278096 233300
rect 212448 233180 212500 233232
rect 219808 233180 219860 233232
rect 226432 233180 226484 233232
rect 227168 233180 227220 233232
rect 276204 233180 276256 233232
rect 278320 233180 278372 233232
rect 579620 233180 579672 233232
rect 222568 233112 222620 233164
rect 249432 233112 249484 233164
rect 335452 233112 335504 233164
rect 219164 233044 219216 233096
rect 223764 233044 223816 233096
rect 245200 233044 245252 233096
rect 300308 233044 300360 233096
rect 194416 232840 194468 232892
rect 219716 232976 219768 233028
rect 252560 232976 252612 233028
rect 253204 232976 253256 233028
rect 304540 232976 304592 233028
rect 248880 232908 248932 232960
rect 296260 232908 296312 232960
rect 252284 232840 252336 232892
rect 297732 232840 297784 232892
rect 159548 232772 159600 232824
rect 209412 232772 209464 232824
rect 235540 232772 235592 232824
rect 274272 232772 274324 232824
rect 277860 232772 277912 232824
rect 281080 232772 281132 232824
rect 156880 232704 156932 232756
rect 207020 232704 207072 232756
rect 232504 232704 232556 232756
rect 240968 232704 241020 232756
rect 275284 232704 275336 232756
rect 161480 232636 161532 232688
rect 191656 232636 191708 232688
rect 195888 232636 195940 232688
rect 256056 232636 256108 232688
rect 261208 232636 261260 232688
rect 287152 232636 287204 232688
rect 287612 232636 287664 232688
rect 155684 232568 155736 232620
rect 231676 232568 231728 232620
rect 240324 232568 240376 232620
rect 240968 232568 241020 232620
rect 241704 232568 241756 232620
rect 242716 232568 242768 232620
rect 249156 232568 249208 232620
rect 278412 232568 278464 232620
rect 279240 232568 279292 232620
rect 157064 232500 157116 232552
rect 234620 232500 234672 232552
rect 253572 232500 253624 232552
rect 284024 232500 284076 232552
rect 328552 232500 328604 232552
rect 225696 232432 225748 232484
rect 226800 232432 226852 232484
rect 233700 232432 233752 232484
rect 234252 232432 234304 232484
rect 247500 232432 247552 232484
rect 271144 232432 271196 232484
rect 280252 232432 280304 232484
rect 282552 232432 282604 232484
rect 243176 232364 243228 232416
rect 260196 232364 260248 232416
rect 269304 232364 269356 232416
rect 236736 232296 236788 232348
rect 239680 232296 239732 232348
rect 280620 232296 280672 232348
rect 242072 232160 242124 232212
rect 242440 232160 242492 232212
rect 229468 231888 229520 231940
rect 230388 231888 230440 231940
rect 227996 231820 228048 231872
rect 230756 231820 230808 231872
rect 254768 231820 254820 231872
rect 264520 231820 264572 231872
rect 209504 231752 209556 231804
rect 229652 231752 229704 231804
rect 242624 231752 242676 231804
rect 243636 231752 243688 231804
rect 261576 231752 261628 231804
rect 262404 231752 262456 231804
rect 262496 231752 262548 231804
rect 269672 231752 269724 231804
rect 284392 231752 284444 231804
rect 285128 231752 285180 231804
rect 291292 231752 291344 231804
rect 291936 231752 291988 231804
rect 230756 231684 230808 231736
rect 230940 231684 230992 231736
rect 240968 231684 241020 231736
rect 300492 231684 300544 231736
rect 246764 231616 246816 231668
rect 248788 231616 248840 231668
rect 256792 231616 256844 231668
rect 316868 231616 316920 231668
rect 250076 231548 250128 231600
rect 250812 231548 250864 231600
rect 294880 231548 294932 231600
rect 234528 231480 234580 231532
rect 261760 231480 261812 231532
rect 262404 231480 262456 231532
rect 305184 231480 305236 231532
rect 252376 231412 252428 231464
rect 284392 231412 284444 231464
rect 291200 231412 291252 231464
rect 292304 231412 292356 231464
rect 234068 231344 234120 231396
rect 234436 231344 234488 231396
rect 246856 231344 246908 231396
rect 277584 231344 277636 231396
rect 277860 231344 277912 231396
rect 199844 231276 199896 231328
rect 259092 231276 259144 231328
rect 262496 231276 262548 231328
rect 267188 231276 267240 231328
rect 291200 231276 291252 231328
rect 164148 231208 164200 231260
rect 223120 231208 223172 231260
rect 227352 231208 227404 231260
rect 266176 231208 266228 231260
rect 266452 231208 266504 231260
rect 291292 231208 291344 231260
rect 199936 231140 199988 231192
rect 259644 231140 259696 231192
rect 262312 231140 262364 231192
rect 263232 231140 263284 231192
rect 264520 231140 264572 231192
rect 278964 231140 279016 231192
rect 279516 231140 279568 231192
rect 198648 231072 198700 231124
rect 258540 231072 258592 231124
rect 258816 231072 258868 231124
rect 280160 231072 280212 231124
rect 332692 231072 332744 231124
rect 248144 231004 248196 231056
rect 276204 231004 276256 231056
rect 226616 230936 226668 230988
rect 227536 230936 227588 230988
rect 232596 230936 232648 230988
rect 233608 230936 233660 230988
rect 250904 230936 250956 230988
rect 329840 230936 329892 230988
rect 251732 230868 251784 230920
rect 252284 230868 252336 230920
rect 256792 230868 256844 230920
rect 257068 230868 257120 230920
rect 199752 230528 199804 230580
rect 258264 230664 258316 230716
rect 265440 230596 265492 230648
rect 265900 230596 265952 230648
rect 239312 230528 239364 230580
rect 239588 230528 239640 230580
rect 198464 230460 198516 230512
rect 254492 230528 254544 230580
rect 228916 230392 228968 230444
rect 236000 230392 236052 230444
rect 244096 230392 244148 230444
rect 244832 230392 244884 230444
rect 245292 230392 245344 230444
rect 249248 230460 249300 230512
rect 249064 230392 249116 230444
rect 301504 230392 301556 230444
rect 305644 230392 305696 230444
rect 306012 230392 306064 230444
rect 230020 230324 230072 230376
rect 240968 230324 241020 230376
rect 244004 230324 244056 230376
rect 304448 230324 304500 230376
rect 217784 230256 217836 230308
rect 237104 230256 237156 230308
rect 241336 230256 241388 230308
rect 300216 230256 300268 230308
rect 223212 230188 223264 230240
rect 239128 230188 239180 230240
rect 239404 230188 239456 230240
rect 240048 230188 240100 230240
rect 249064 230188 249116 230240
rect 212448 230120 212500 230172
rect 239864 230120 239916 230172
rect 244740 230120 244792 230172
rect 245292 230120 245344 230172
rect 247408 230120 247460 230172
rect 305644 230188 305696 230240
rect 249248 230120 249300 230172
rect 301688 230120 301740 230172
rect 162216 229780 162268 229832
rect 235908 230052 235960 230104
rect 288256 230052 288308 230104
rect 236000 229984 236052 230036
rect 237196 229984 237248 230036
rect 287980 229984 288032 230036
rect 239128 229916 239180 229968
rect 247408 229916 247460 229968
rect 247592 229916 247644 229968
rect 287796 229916 287848 229968
rect 225420 229848 225472 229900
rect 225788 229848 225840 229900
rect 225972 229848 226024 229900
rect 228364 229780 228416 229832
rect 228732 229780 228784 229832
rect 232964 229848 233016 229900
rect 276664 229848 276716 229900
rect 160928 229712 160980 229764
rect 236092 229712 236144 229764
rect 240876 229780 240928 229832
rect 247592 229780 247644 229832
rect 249248 229780 249300 229832
rect 279608 229780 279660 229832
rect 236552 229712 236604 229764
rect 235264 229644 235316 229696
rect 240876 229644 240928 229696
rect 245292 229644 245344 229696
rect 245568 229644 245620 229696
rect 245752 229644 245804 229696
rect 246672 229644 246724 229696
rect 269856 229712 269908 229764
rect 274732 229712 274784 229764
rect 275376 229712 275428 229764
rect 275928 229712 275980 229764
rect 277032 229712 277084 229764
rect 251272 229576 251324 229628
rect 252468 229576 252520 229628
rect 273996 229644 274048 229696
rect 212356 229508 212408 229560
rect 236736 229508 236788 229560
rect 239864 229508 239916 229560
rect 249248 229508 249300 229560
rect 247500 229440 247552 229492
rect 248328 229440 248380 229492
rect 245016 229372 245068 229424
rect 248604 229304 248656 229356
rect 249248 229304 249300 229356
rect 249524 229304 249576 229356
rect 274732 229576 274784 229628
rect 262864 229508 262916 229560
rect 280252 229508 280304 229560
rect 252744 229236 252796 229288
rect 253756 229236 253808 229288
rect 222936 229168 222988 229220
rect 236460 229168 236512 229220
rect 227536 229100 227588 229152
rect 244096 229100 244148 229152
rect 271144 229100 271196 229152
rect 277400 229100 277452 229152
rect 208308 229032 208360 229084
rect 230296 229032 230348 229084
rect 258448 229032 258500 229084
rect 338212 229032 338264 229084
rect 230572 228964 230624 229016
rect 231308 228964 231360 229016
rect 233332 228964 233384 229016
rect 233792 228964 233844 229016
rect 260104 228964 260156 229016
rect 335360 228964 335412 229016
rect 161572 228896 161624 228948
rect 215208 228896 215260 228948
rect 231124 228896 231176 228948
rect 236828 228896 236880 228948
rect 263508 228896 263560 228948
rect 327264 228896 327316 228948
rect 154028 228828 154080 228880
rect 208308 228828 208360 228880
rect 152740 228760 152792 228812
rect 209504 228760 209556 228812
rect 213736 228760 213788 228812
rect 239036 228760 239088 228812
rect 299020 228828 299072 228880
rect 249156 228760 249208 228812
rect 258448 228760 258500 228812
rect 265624 228760 265676 228812
rect 268200 228760 268252 228812
rect 327908 228760 327960 228812
rect 155592 228624 155644 228676
rect 225604 228624 225656 228676
rect 239680 228624 239732 228676
rect 259920 228692 259972 228744
rect 301872 228692 301924 228744
rect 264704 228624 264756 228676
rect 325148 228624 325200 228676
rect 201224 228556 201276 228608
rect 271880 228556 271932 228608
rect 152832 228488 152884 228540
rect 225236 228488 225288 228540
rect 234436 228488 234488 228540
rect 295248 228488 295300 228540
rect 197912 228420 197964 228472
rect 271972 228420 272024 228472
rect 160836 228352 160888 228404
rect 237840 228352 237892 228404
rect 239772 228352 239824 228404
rect 260104 228352 260156 228404
rect 266544 228352 266596 228404
rect 267188 228352 267240 228404
rect 232688 228284 232740 228336
rect 288164 228284 288216 228336
rect 233700 228216 233752 228268
rect 234160 228216 234212 228268
rect 235540 228216 235592 228268
rect 286508 228216 286560 228268
rect 236460 228148 236512 228200
rect 273628 228148 273680 228200
rect 202604 228080 202656 228132
rect 272432 228080 272484 228132
rect 234804 227740 234856 227792
rect 235540 227740 235592 227792
rect 262864 227740 262916 227792
rect 263508 227740 263560 227792
rect 215116 227536 215168 227588
rect 260564 227672 260616 227724
rect 321008 227672 321060 227724
rect 262956 227604 263008 227656
rect 323860 227604 323912 227656
rect 263232 227536 263284 227588
rect 323768 227536 323820 227588
rect 228180 227468 228232 227520
rect 228640 227468 228692 227520
rect 260932 227468 260984 227520
rect 321652 227468 321704 227520
rect 234712 227400 234764 227452
rect 294604 227400 294656 227452
rect 223028 227264 223080 227316
rect 239312 227332 239364 227384
rect 289176 227332 289228 227384
rect 251088 227264 251140 227316
rect 278228 227264 278280 227316
rect 287520 227264 287572 227316
rect 336832 227264 336884 227316
rect 226984 227196 227036 227248
rect 257068 227196 257120 227248
rect 258356 227196 258408 227248
rect 292672 227196 292724 227248
rect 256608 227128 256660 227180
rect 282368 227128 282420 227180
rect 234344 227060 234396 227112
rect 236000 227060 236052 227112
rect 280896 227060 280948 227112
rect 155408 226992 155460 227044
rect 210976 226992 211028 227044
rect 211712 226992 211764 227044
rect 269396 226992 269448 227044
rect 255780 226924 255832 226976
rect 289268 226924 289320 226976
rect 333060 227060 333112 227112
rect 292672 226992 292724 227044
rect 293224 226992 293276 227044
rect 336924 226992 336976 227044
rect 239864 226856 239916 226908
rect 265532 226856 265584 226908
rect 265808 226856 265860 226908
rect 285772 226856 285824 226908
rect 262036 226788 262088 226840
rect 282000 226788 282052 226840
rect 250628 226720 250680 226772
rect 251088 226720 251140 226772
rect 265716 226652 265768 226704
rect 266268 226652 266320 226704
rect 285772 226652 285824 226704
rect 286968 226652 287020 226704
rect 250812 226584 250864 226636
rect 251088 226584 251140 226636
rect 234712 226516 234764 226568
rect 235448 226516 235500 226568
rect 260104 226312 260156 226364
rect 260932 226312 260984 226364
rect 281540 226312 281592 226364
rect 282000 226312 282052 226364
rect 287520 226312 287572 226364
rect 287796 226312 287848 226364
rect 202696 226244 202748 226296
rect 227076 226244 227128 226296
rect 249892 226244 249944 226296
rect 250536 226244 250588 226296
rect 258264 226244 258316 226296
rect 345020 226244 345072 226296
rect 266268 226176 266320 226228
rect 342260 226176 342312 226228
rect 241152 226108 241204 226160
rect 301780 226108 301832 226160
rect 246304 226040 246356 226092
rect 307024 226040 307076 226092
rect 245476 225972 245528 226024
rect 305736 225972 305788 226024
rect 250444 225904 250496 225956
rect 309968 225904 310020 225956
rect 245200 225836 245252 225888
rect 245476 225836 245528 225888
rect 250536 225836 250588 225888
rect 310060 225836 310112 225888
rect 255596 225768 255648 225820
rect 255964 225768 256016 225820
rect 315672 225768 315724 225820
rect 243912 225700 243964 225752
rect 302976 225700 303028 225752
rect 234252 225632 234304 225684
rect 240508 225632 240560 225684
rect 295984 225632 296036 225684
rect 156788 225564 156840 225616
rect 202696 225564 202748 225616
rect 244096 225564 244148 225616
rect 296720 225564 296772 225616
rect 297364 225564 297416 225616
rect 241704 225496 241756 225548
rect 242716 225496 242768 225548
rect 285036 225496 285088 225548
rect 242532 225428 242584 225480
rect 284116 225428 284168 225480
rect 243820 225360 243872 225412
rect 282644 225360 282696 225412
rect 243544 225020 243596 225072
rect 243820 225020 243872 225072
rect 240876 224952 240928 225004
rect 241152 224952 241204 225004
rect 242164 224952 242216 225004
rect 242532 224952 242584 225004
rect 243636 224952 243688 225004
rect 243912 224952 243964 225004
rect 248972 224952 249024 225004
rect 249340 224952 249392 225004
rect 222016 224884 222068 224936
rect 298008 224884 298060 224936
rect 236736 224816 236788 224868
rect 237288 224816 237340 224868
rect 301596 224816 301648 224868
rect 234160 224748 234212 224800
rect 298284 224748 298336 224800
rect 225880 224680 225932 224732
rect 245108 224680 245160 224732
rect 252008 224680 252060 224732
rect 312820 224680 312872 224732
rect 209412 224272 209464 224324
rect 238576 224612 238628 224664
rect 298744 224612 298796 224664
rect 239588 224544 239640 224596
rect 299572 224544 299624 224596
rect 240968 224476 241020 224528
rect 300124 224476 300176 224528
rect 232872 224408 232924 224460
rect 285220 224408 285272 224460
rect 243728 224340 243780 224392
rect 293316 224340 293368 224392
rect 240692 224272 240744 224324
rect 242900 224272 242952 224324
rect 297456 224272 297508 224324
rect 160744 224204 160796 224256
rect 237656 224204 237708 224256
rect 240784 224204 240836 224256
rect 241244 224204 241296 224256
rect 242072 224204 242124 224256
rect 244280 224204 244332 224256
rect 302884 224204 302936 224256
rect 230204 224136 230256 224188
rect 230664 224136 230716 224188
rect 238208 224136 238260 224188
rect 283748 224136 283800 224188
rect 241244 224068 241296 224120
rect 286692 224068 286744 224120
rect 238024 224000 238076 224052
rect 247224 224000 247276 224052
rect 252836 224000 252888 224052
rect 253296 224000 253348 224052
rect 272616 224000 272668 224052
rect 264336 223932 264388 223984
rect 264612 223932 264664 223984
rect 264152 223864 264204 223916
rect 264428 223864 264480 223916
rect 251456 223524 251508 223576
rect 252192 223524 252244 223576
rect 259000 223524 259052 223576
rect 319720 223524 319772 223576
rect 251364 223456 251416 223508
rect 251916 223456 251968 223508
rect 256884 223456 256936 223508
rect 257344 223456 257396 223508
rect 318340 223456 318392 223508
rect 256700 223388 256752 223440
rect 257436 223388 257488 223440
rect 318248 223388 318300 223440
rect 256056 223320 256108 223372
rect 256424 223320 256476 223372
rect 316684 223320 316736 223372
rect 260472 223252 260524 223304
rect 319444 223252 319496 223304
rect 258908 223184 258960 223236
rect 318156 223184 318208 223236
rect 251916 223116 251968 223168
rect 311256 223116 311308 223168
rect 252192 223048 252244 223100
rect 311164 223048 311216 223100
rect 155500 222844 155552 222896
rect 226616 222980 226668 223032
rect 280804 222980 280856 223032
rect 303620 222980 303672 223032
rect 304356 222980 304408 223032
rect 245844 222844 245896 222896
rect 246304 222844 246356 222896
rect 303620 222844 303672 222896
rect 251272 222096 251324 222148
rect 252100 222096 252152 222148
rect 252744 222096 252796 222148
rect 253388 222096 253440 222148
rect 252652 222028 252704 222080
rect 253572 222028 253624 222080
rect 254400 222096 254452 222148
rect 254768 222096 254820 222148
rect 340972 222096 341024 222148
rect 336740 222028 336792 222080
rect 254308 221960 254360 222012
rect 254860 221960 254912 222012
rect 254952 221960 255004 222012
rect 312912 221960 312964 222012
rect 314292 221892 314344 221944
rect 227076 221824 227128 221876
rect 248512 221824 248564 221876
rect 252100 221824 252152 221876
rect 254952 221824 255004 221876
rect 255044 221824 255096 221876
rect 314108 221824 314160 221876
rect 230112 221756 230164 221808
rect 254032 221756 254084 221808
rect 254216 221756 254268 221808
rect 254676 221756 254728 221808
rect 314200 221756 314252 221808
rect 223120 221688 223172 221740
rect 250260 221688 250312 221740
rect 253388 221688 253440 221740
rect 307208 221688 307260 221740
rect 158260 221484 158312 221536
rect 233700 221620 233752 221672
rect 283840 221620 283892 221672
rect 234988 221552 235040 221604
rect 276388 221552 276440 221604
rect 242624 221484 242676 221536
rect 272432 221484 272484 221536
rect 286324 221484 286376 221536
rect 160652 221416 160704 221468
rect 238300 221416 238352 221468
rect 254032 221416 254084 221468
rect 255044 221416 255096 221468
rect 260840 221416 260892 221468
rect 294604 221416 294656 221468
rect 320824 221416 320876 221468
rect 248972 220736 249024 220788
rect 249340 220736 249392 220788
rect 258724 220736 258776 220788
rect 338120 220736 338172 220788
rect 247040 220668 247092 220720
rect 247684 220668 247736 220720
rect 307116 220668 307168 220720
rect 226064 220600 226116 220652
rect 279424 220600 279476 220652
rect 246672 220532 246724 220584
rect 281172 220532 281224 220584
rect 225512 220260 225564 220312
rect 226064 220260 226116 220312
rect 257620 220124 257672 220176
rect 283748 220124 283800 220176
rect 318064 220124 318116 220176
rect 232780 220056 232832 220108
rect 247040 220056 247092 220108
rect 249340 220056 249392 220108
rect 309784 220056 309836 220108
rect 231860 219376 231912 219428
rect 232320 219376 232372 219428
rect 292580 219376 292632 219428
rect 256424 219308 256476 219360
rect 315304 219308 315356 219360
rect 246580 219240 246632 219292
rect 304264 219240 304316 219292
rect 238392 219172 238444 219224
rect 290464 219172 290516 219224
rect 255136 219104 255188 219156
rect 294696 219104 294748 219156
rect 253756 219036 253808 219088
rect 288072 219036 288124 219088
rect 253940 218900 253992 218952
rect 254952 218900 255004 218952
rect 158168 218696 158220 218748
rect 231860 218696 231912 218748
rect 254952 218696 255004 218748
rect 313924 218696 313976 218748
rect 238116 218084 238168 218136
rect 238392 218084 238444 218136
rect 246580 218084 246632 218136
rect 246856 218084 246908 218136
rect 158076 218016 158128 218068
rect 230572 218016 230624 218068
rect 231492 218016 231544 218068
rect 236920 218016 236972 218068
rect 240968 218016 241020 218068
rect 204076 217948 204128 218000
rect 223580 217948 223632 218000
rect 227168 217948 227220 218000
rect 227720 217948 227772 218000
rect 187516 217336 187568 217388
rect 215024 217336 215076 217388
rect 227720 217336 227772 217388
rect 287888 217336 287940 217388
rect 151544 217268 151596 217320
rect 204076 217268 204128 217320
rect 247132 217268 247184 217320
rect 247684 217268 247736 217320
rect 308404 217268 308456 217320
rect 226800 216588 226852 216640
rect 227168 216588 227220 216640
rect 228456 216588 228508 216640
rect 228640 216588 228692 216640
rect 228732 216588 228784 216640
rect 292856 216588 292908 216640
rect 227996 216452 228048 216504
rect 228640 216452 228692 216504
rect 246488 216520 246540 216572
rect 247868 216520 247920 216572
rect 307116 216520 307168 216572
rect 307484 216520 307536 216572
rect 286416 216452 286468 216504
rect 228456 216384 228508 216436
rect 283656 216384 283708 216436
rect 228640 216316 228692 216368
rect 283932 216316 283984 216368
rect 225328 216248 225380 216300
rect 228732 216248 228784 216300
rect 230572 216248 230624 216300
rect 282184 216248 282236 216300
rect 193404 216044 193456 216096
rect 209044 216044 209096 216096
rect 180892 215976 180944 216028
rect 217232 215976 217284 216028
rect 161664 215908 161716 215960
rect 222292 215908 222344 215960
rect 205732 215228 205784 215280
rect 206836 215228 206888 215280
rect 228180 215228 228232 215280
rect 205640 215160 205692 215212
rect 206928 215160 206980 215212
rect 226892 215160 226944 215212
rect 183100 214752 183152 214804
rect 214748 214752 214800 214804
rect 157984 214684 158036 214736
rect 205640 214684 205692 214736
rect 156696 214616 156748 214668
rect 205732 214616 205784 214668
rect 167000 214548 167052 214600
rect 167736 214548 167788 214600
rect 168380 214548 168432 214600
rect 168840 214548 168892 214600
rect 168472 214480 168524 214532
rect 169208 214480 169260 214532
rect 161756 214412 161808 214464
rect 222200 214548 222252 214600
rect 171140 214480 171192 214532
rect 172152 214480 172204 214532
rect 172520 214480 172572 214532
rect 173256 214480 173308 214532
rect 178040 214480 178092 214532
rect 178776 214480 178828 214532
rect 180800 214480 180852 214532
rect 181352 214480 181404 214532
rect 182272 214480 182324 214532
rect 183192 214480 183244 214532
rect 183560 214480 183612 214532
rect 184296 214480 184348 214532
rect 185032 214480 185084 214532
rect 185400 214480 185452 214532
rect 186320 214480 186372 214532
rect 186504 214480 186556 214532
rect 187700 214480 187752 214532
rect 188344 214480 188396 214532
rect 189080 214480 189132 214532
rect 189816 214480 189868 214532
rect 190460 214480 190512 214532
rect 190920 214480 190972 214532
rect 191932 214480 191984 214532
rect 192392 214480 192444 214532
rect 193312 214480 193364 214532
rect 193864 214480 193916 214532
rect 194600 214480 194652 214532
rect 195336 214480 195388 214532
rect 183652 214412 183704 214464
rect 183928 214412 183980 214464
rect 184940 214412 184992 214464
rect 185216 214412 185268 214464
rect 187792 214412 187844 214464
rect 188712 214412 188764 214464
rect 186044 214208 186096 214260
rect 189908 214208 189960 214260
rect 202880 214004 202932 214056
rect 203156 214004 203208 214056
rect 3148 213936 3200 213988
rect 200672 213868 200724 213920
rect 202880 213868 202932 213920
rect 204168 213868 204220 213920
rect 224408 213868 224460 213920
rect 177212 213392 177264 213444
rect 209136 213392 209188 213444
rect 181996 213324 182048 213376
rect 214656 213324 214708 213376
rect 153936 213256 153988 213308
rect 202880 213256 202932 213308
rect 184848 213188 184900 213240
rect 244004 213188 244056 213240
rect 249248 213188 249300 213240
rect 335360 213188 335412 213240
rect 336004 213188 336056 213240
rect 194692 212712 194744 212764
rect 194968 212712 195020 212764
rect 159272 212508 159324 212560
rect 163504 212508 163556 212560
rect 165620 212440 165672 212492
rect 170404 212440 170456 212492
rect 177580 212440 177632 212492
rect 178684 212440 178736 212492
rect 187884 212440 187936 212492
rect 189724 212440 189776 212492
rect 186320 212372 186372 212424
rect 200580 212440 200632 212492
rect 200672 212440 200724 212492
rect 219900 212440 219952 212492
rect 196348 212372 196400 212424
rect 162032 212304 162084 212356
rect 162768 212304 162820 212356
rect 179788 212236 179840 212288
rect 189632 212236 189684 212288
rect 176476 212168 176528 212220
rect 200764 212304 200816 212356
rect 197452 212236 197504 212288
rect 198556 212236 198608 212288
rect 198924 212236 198976 212288
rect 200028 212236 200080 212288
rect 200580 212236 200632 212288
rect 202696 212304 202748 212356
rect 203708 212304 203760 212356
rect 211804 212304 211856 212356
rect 201224 212236 201276 212288
rect 202604 212236 202656 212288
rect 202788 212236 202840 212288
rect 203340 212236 203392 212288
rect 199292 212168 199344 212220
rect 221924 212236 221976 212288
rect 175740 212100 175792 212152
rect 180064 212100 180116 212152
rect 174636 212032 174688 212084
rect 186964 212100 187016 212152
rect 189724 212100 189776 212152
rect 221832 212100 221884 212152
rect 172060 211964 172112 212016
rect 212264 212032 212316 212084
rect 180524 211964 180576 212016
rect 221740 211964 221792 212016
rect 161940 211896 161992 211948
rect 162676 211896 162728 211948
rect 166540 211896 166592 211948
rect 167644 211896 167696 211948
rect 168288 211896 168340 211948
rect 175372 211896 175424 211948
rect 217692 211896 217744 211948
rect 156604 211828 156656 211880
rect 201500 211828 201552 211880
rect 11704 211760 11756 211812
rect 201224 211760 201276 211812
rect 189080 211692 189132 211744
rect 202788 211692 202840 211744
rect 95884 211488 95936 211540
rect 204812 211488 204864 211540
rect 272248 211760 272300 211812
rect 170128 211420 170180 211472
rect 187608 211420 187660 211472
rect 168748 211352 168800 211404
rect 182548 211352 182600 211404
rect 168288 211284 168340 211336
rect 189540 211284 189592 211336
rect 191748 211284 191800 211336
rect 202144 211284 202196 211336
rect 183468 211216 183520 211268
rect 206284 211216 206336 211268
rect 162032 211148 162084 211200
rect 165436 211148 165488 211200
rect 195980 211012 196032 211064
rect 196440 211012 196492 211064
rect 200120 210740 200172 210792
rect 201132 210740 201184 210792
rect 174268 210672 174320 210724
rect 212080 210672 212132 210724
rect 3424 210604 3476 210656
rect 183468 210604 183520 210656
rect 3608 210536 3660 210588
rect 186320 210536 186372 210588
rect 197360 210536 197412 210588
rect 197636 210536 197688 210588
rect 3516 210468 3568 210520
rect 189080 210468 189132 210520
rect 3700 210400 3752 210452
rect 191748 210400 191800 210452
rect 193220 210264 193272 210316
rect 194508 210264 194560 210316
rect 160560 209924 160612 209976
rect 200948 209924 201000 209976
rect 159364 209856 159416 209908
rect 201684 209856 201736 209908
rect 202420 209924 202472 209976
rect 155224 209788 155276 209840
rect 204628 209788 204680 209840
rect 187700 209720 187752 209772
rect 219256 209720 219308 209772
rect 199200 209584 199252 209636
rect 199844 209584 199896 209636
rect 142804 209176 142856 209228
rect 202880 209380 202932 209432
rect 203156 209380 203208 209432
rect 203892 209380 203944 209432
rect 120724 209108 120776 209160
rect 204352 209380 204404 209432
rect 204996 209380 205048 209432
rect 43444 209040 43496 209092
rect 219256 209040 219308 209092
rect 579988 209040 580040 209092
rect 209136 207748 209188 207800
rect 263232 207748 263284 207800
rect 209504 207680 209556 207732
rect 264336 207680 264388 207732
rect 209044 207612 209096 207664
rect 265808 207612 265860 207664
rect 210792 206252 210844 206304
rect 263324 206252 263376 206304
rect 245660 204212 245712 204264
rect 246764 204212 246816 204264
rect 327724 204212 327776 204264
rect 237012 203532 237064 203584
rect 245660 203532 245712 203584
rect 3332 202784 3384 202836
rect 156604 202784 156656 202836
rect 209596 202104 209648 202156
rect 259092 202104 259144 202156
rect 247040 200064 247092 200116
rect 248144 200064 248196 200116
rect 342260 200064 342312 200116
rect 342260 199452 342312 199504
rect 342904 199452 342956 199504
rect 235816 199384 235868 199436
rect 247040 199384 247092 199436
rect 210884 196596 210936 196648
rect 224132 196596 224184 196648
rect 338764 193128 338816 193180
rect 580172 193128 580224 193180
rect 210976 192448 211028 192500
rect 223396 192448 223448 192500
rect 3332 188980 3384 189032
rect 160560 188980 160612 189032
rect 211068 186940 211120 186992
rect 224040 186940 224092 186992
rect 242716 186940 242768 186992
rect 259460 186940 259512 186992
rect 257528 186328 257580 186380
rect 257804 186328 257856 186380
rect 443000 186328 443052 186380
rect 230204 184152 230256 184204
rect 250720 184152 250772 184204
rect 361580 184152 361632 184204
rect 209688 177284 209740 177336
rect 266360 177284 266412 177336
rect 246580 176672 246632 176724
rect 246856 176672 246908 176724
rect 305000 176672 305052 176724
rect 259368 175244 259420 175296
rect 467840 175244 467892 175296
rect 256240 173952 256292 174004
rect 256516 173952 256568 174004
rect 425060 173952 425112 174004
rect 256148 173884 256200 173936
rect 432052 173884 432104 173936
rect 208952 173136 209004 173188
rect 262312 173136 262364 173188
rect 245292 171096 245344 171148
rect 298100 171096 298152 171148
rect 260380 169736 260432 169788
rect 481732 169736 481784 169788
rect 245384 168376 245436 168428
rect 287060 168376 287112 168428
rect 257620 167016 257672 167068
rect 257988 167016 258040 167068
rect 447140 167016 447192 167068
rect 156972 166336 157024 166388
rect 156880 166132 156932 166184
rect 253756 165588 253808 165640
rect 397460 165588 397512 165640
rect 209780 164840 209832 164892
rect 226064 164840 226116 164892
rect 161572 161508 161624 161560
rect 162400 161508 162452 161560
rect 158628 160624 158680 160676
rect 161848 160624 161900 160676
rect 160008 160488 160060 160540
rect 162308 160420 162360 160472
rect 156972 160352 157024 160404
rect 159180 160284 159232 160336
rect 158076 159944 158128 159996
rect 152464 159876 152516 159928
rect 152832 159876 152884 159928
rect 161756 159876 161808 159928
rect 162584 159876 162636 159928
rect 159180 159808 159232 159860
rect 161664 159808 161716 159860
rect 162676 159808 162728 159860
rect 162492 159740 162544 159792
rect 161204 159672 161256 159724
rect 156512 159604 156564 159656
rect 156972 159604 157024 159656
rect 158352 159604 158404 159656
rect 162676 159604 162728 159656
rect 162952 159672 163004 159724
rect 163412 159808 163464 159860
rect 164792 159876 164844 159928
rect 165804 159876 165856 159928
rect 167736 159876 167788 159928
rect 167828 159876 167880 159928
rect 207480 161236 207532 161288
rect 207664 161100 207716 161152
rect 249340 161100 249392 161152
rect 225604 161032 225656 161084
rect 208400 160964 208452 161016
rect 250628 160964 250680 161016
rect 207480 160896 207532 160948
rect 229744 160896 229796 160948
rect 230756 160828 230808 160880
rect 249064 160760 249116 160812
rect 253204 160692 253256 160744
rect 170404 159876 170456 159928
rect 170496 159808 170548 159860
rect 163688 159740 163740 159792
rect 164792 159740 164844 159792
rect 165436 159740 165488 159792
rect 165620 159740 165672 159792
rect 170864 159876 170916 159928
rect 170956 159876 171008 159928
rect 171416 159876 171468 159928
rect 171876 159876 171928 159928
rect 174360 159876 174412 159928
rect 174452 159876 174504 159928
rect 171048 159672 171100 159724
rect 165436 159604 165488 159656
rect 153016 159536 153068 159588
rect 169944 159536 169996 159588
rect 170220 159604 170272 159656
rect 171232 159604 171284 159656
rect 171324 159536 171376 159588
rect 171968 159740 172020 159792
rect 172704 159808 172756 159860
rect 173348 159808 173400 159860
rect 172888 159740 172940 159792
rect 172612 159672 172664 159724
rect 173348 159672 173400 159724
rect 174452 159672 174504 159724
rect 171876 159604 171928 159656
rect 171784 159536 171836 159588
rect 174360 159604 174412 159656
rect 174728 159876 174780 159928
rect 174820 159876 174872 159928
rect 178500 159876 178552 159928
rect 183100 159808 183152 159860
rect 188988 159808 189040 159860
rect 191748 159876 191800 159928
rect 193128 159876 193180 159928
rect 199292 159876 199344 159928
rect 203432 159876 203484 159928
rect 209136 160216 209188 160268
rect 182548 159740 182600 159792
rect 191104 159740 191156 159792
rect 208400 160148 208452 160200
rect 199016 159740 199068 159792
rect 199292 159740 199344 159792
rect 199384 159740 199436 159792
rect 200212 159740 200264 159792
rect 203248 159740 203300 159792
rect 208124 160080 208176 160132
rect 280804 160080 280856 160132
rect 300860 160080 300912 160132
rect 207848 160012 207900 160064
rect 207756 159944 207808 159996
rect 206192 159876 206244 159928
rect 207020 159876 207072 159928
rect 209688 159876 209740 159928
rect 207112 159808 207164 159860
rect 207572 159808 207624 159860
rect 206284 159740 206336 159792
rect 208308 159740 208360 159792
rect 174912 159604 174964 159656
rect 180064 159604 180116 159656
rect 209320 159604 209372 159656
rect 132500 159468 132552 159520
rect 158628 159468 158680 159520
rect 161296 159468 161348 159520
rect 170772 159468 170824 159520
rect 171600 159468 171652 159520
rect 128360 159400 128412 159452
rect 159272 159400 159324 159452
rect 171416 159400 171468 159452
rect 171692 159400 171744 159452
rect 173992 159400 174044 159452
rect 191012 159536 191064 159588
rect 200212 159536 200264 159588
rect 204076 159536 204128 159588
rect 207020 159536 207072 159588
rect 207480 159536 207532 159588
rect 208216 159536 208268 159588
rect 176108 159400 176160 159452
rect 176292 159400 176344 159452
rect 183744 159468 183796 159520
rect 202696 159468 202748 159520
rect 205180 159468 205232 159520
rect 205364 159468 205416 159520
rect 206192 159468 206244 159520
rect 235632 159468 235684 159520
rect 207940 159400 207992 159452
rect 96620 159332 96672 159384
rect 152740 159332 152792 159384
rect 153016 159332 153068 159384
rect 162768 159332 162820 159384
rect 163504 159332 163556 159384
rect 171876 159332 171928 159384
rect 174728 159332 174780 159384
rect 175096 159332 175148 159384
rect 187700 159332 187752 159384
rect 228364 159332 228416 159384
rect 153936 159264 153988 159316
rect 164240 159264 164292 159316
rect 164792 159264 164844 159316
rect 165804 159264 165856 159316
rect 166080 159264 166132 159316
rect 166816 159264 166868 159316
rect 170404 159264 170456 159316
rect 170588 159264 170640 159316
rect 170956 159264 171008 159316
rect 171232 159264 171284 159316
rect 175280 159264 175332 159316
rect 176108 159264 176160 159316
rect 210148 159264 210200 159316
rect 154120 159196 154172 159248
rect 164148 159196 164200 159248
rect 166172 159196 166224 159248
rect 222384 159196 222436 159248
rect 162676 159128 162728 159180
rect 164792 159128 164844 159180
rect 165896 159128 165948 159180
rect 166080 159128 166132 159180
rect 161848 159060 161900 159112
rect 162952 159060 163004 159112
rect 163136 159060 163188 159112
rect 163688 159060 163740 159112
rect 164424 159060 164476 159112
rect 164700 159060 164752 159112
rect 223304 159128 223356 159180
rect 169760 159060 169812 159112
rect 170588 159060 170640 159112
rect 155592 158992 155644 159044
rect 162216 158992 162268 159044
rect 171324 158992 171376 159044
rect 171416 158992 171468 159044
rect 172428 158992 172480 159044
rect 174728 158992 174780 159044
rect 165344 158924 165396 158976
rect 162860 158856 162912 158908
rect 163136 158856 163188 158908
rect 163228 158856 163280 158908
rect 163412 158856 163464 158908
rect 172612 158924 172664 158976
rect 175280 158992 175332 159044
rect 175648 158992 175700 159044
rect 185124 159060 185176 159112
rect 245016 159060 245068 159112
rect 229192 158992 229244 159044
rect 180064 158924 180116 158976
rect 190920 158924 190972 158976
rect 200212 158924 200264 158976
rect 158628 158788 158680 158840
rect 170772 158856 170824 158908
rect 176660 158856 176712 158908
rect 192944 158856 192996 158908
rect 193312 158856 193364 158908
rect 253664 158924 253716 158976
rect 200856 158856 200908 158908
rect 269120 158856 269172 158908
rect 270224 158856 270276 158908
rect 164792 158788 164844 158840
rect 171232 158788 171284 158840
rect 171324 158788 171376 158840
rect 162860 158720 162912 158772
rect 164056 158720 164108 158772
rect 167368 158720 167420 158772
rect 167828 158720 167880 158772
rect 168748 158720 168800 158772
rect 174728 158720 174780 158772
rect 158352 158652 158404 158704
rect 164700 158652 164752 158704
rect 167092 158652 167144 158704
rect 171692 158652 171744 158704
rect 156696 158516 156748 158568
rect 168564 158584 168616 158636
rect 171324 158584 171376 158636
rect 171600 158584 171652 158636
rect 171968 158584 172020 158636
rect 172428 158584 172480 158636
rect 174084 158584 174136 158636
rect 174820 158584 174872 158636
rect 175004 158584 175056 158636
rect 163136 158516 163188 158568
rect 163596 158516 163648 158568
rect 161020 158448 161072 158500
rect 163688 158448 163740 158500
rect 156604 158380 156656 158432
rect 163872 158380 163924 158432
rect 151084 158312 151136 158364
rect 165160 158516 165212 158568
rect 166080 158516 166132 158568
rect 176384 158788 176436 158840
rect 193128 158788 193180 158840
rect 199384 158788 199436 158840
rect 272340 158788 272392 158840
rect 175740 158720 175792 158772
rect 176016 158720 176068 158772
rect 185860 158720 185912 158772
rect 175464 158652 175516 158704
rect 176384 158652 176436 158704
rect 182732 158652 182784 158704
rect 187424 158652 187476 158704
rect 190460 158652 190512 158704
rect 190920 158652 190972 158704
rect 191012 158652 191064 158704
rect 191564 158652 191616 158704
rect 192392 158652 192444 158704
rect 192668 158652 192720 158704
rect 194600 158652 194652 158704
rect 187148 158584 187200 158636
rect 175464 158516 175516 158568
rect 178500 158516 178552 158568
rect 182732 158516 182784 158568
rect 186872 158516 186924 158568
rect 188528 158516 188580 158568
rect 168012 158448 168064 158500
rect 168288 158448 168340 158500
rect 168564 158448 168616 158500
rect 170220 158448 170272 158500
rect 182456 158448 182508 158500
rect 189724 158448 189776 158500
rect 192024 158584 192076 158636
rect 193680 158584 193732 158636
rect 194876 158584 194928 158636
rect 195704 158584 195756 158636
rect 198924 158584 198976 158636
rect 200028 158584 200080 158636
rect 200672 158652 200724 158704
rect 201224 158652 201276 158704
rect 280804 158720 280856 158772
rect 204260 158652 204312 158704
rect 207664 158652 207716 158704
rect 204076 158584 204128 158636
rect 193772 158516 193824 158568
rect 195244 158516 195296 158568
rect 197360 158516 197412 158568
rect 200856 158516 200908 158568
rect 202144 158516 202196 158568
rect 202604 158516 202656 158568
rect 202696 158516 202748 158568
rect 203340 158516 203392 158568
rect 234528 158584 234580 158636
rect 199660 158448 199712 158500
rect 201776 158448 201828 158500
rect 207388 158516 207440 158568
rect 208308 158516 208360 158568
rect 165988 158380 166040 158432
rect 164884 158312 164936 158364
rect 165068 158312 165120 158364
rect 168748 158312 168800 158364
rect 169300 158312 169352 158364
rect 171048 158312 171100 158364
rect 208860 158380 208912 158432
rect 162124 158244 162176 158296
rect 169392 158244 169444 158296
rect 188804 158244 188856 158296
rect 192668 158244 192720 158296
rect 194048 158244 194100 158296
rect 194508 158244 194560 158296
rect 160836 158176 160888 158228
rect 177948 158176 178000 158228
rect 78680 158108 78732 158160
rect 156696 158108 156748 158160
rect 160652 158108 160704 158160
rect 171784 158108 171836 158160
rect 180524 158108 180576 158160
rect 186320 158108 186372 158160
rect 60740 158040 60792 158092
rect 157984 158040 158036 158092
rect 158628 158040 158680 158092
rect 161388 158040 161440 158092
rect 4160 157972 4212 158024
rect 161480 157972 161532 158024
rect 162584 157972 162636 158024
rect 169392 158040 169444 158092
rect 176108 158040 176160 158092
rect 176292 158040 176344 158092
rect 176016 157972 176068 158024
rect 160744 157904 160796 157956
rect 177396 158040 177448 158092
rect 180800 158040 180852 158092
rect 189172 158176 189224 158228
rect 189356 158176 189408 158228
rect 197912 158176 197964 158228
rect 202420 158176 202472 158228
rect 203708 158244 203760 158296
rect 204168 158244 204220 158296
rect 204260 158176 204312 158228
rect 207848 158244 207900 158296
rect 227444 158244 227496 158296
rect 208032 158176 208084 158228
rect 208400 158176 208452 158228
rect 246488 158176 246540 158228
rect 181352 157972 181404 158024
rect 198280 158108 198332 158160
rect 203248 158108 203300 158160
rect 207940 158108 207992 158160
rect 246304 158108 246356 158160
rect 198004 158040 198056 158092
rect 202788 158040 202840 158092
rect 204812 158040 204864 158092
rect 205364 158040 205416 158092
rect 189172 157972 189224 158024
rect 197084 157972 197136 158024
rect 206284 158040 206336 158092
rect 208032 158040 208084 158092
rect 250444 158040 250496 158092
rect 180524 157904 180576 157956
rect 180708 157904 180760 157956
rect 185216 157904 185268 157956
rect 194876 157904 194928 157956
rect 196164 157904 196216 157956
rect 198188 157904 198240 157956
rect 148324 157836 148376 157888
rect 165620 157836 165672 157888
rect 167828 157836 167880 157888
rect 168564 157836 168616 157888
rect 176016 157836 176068 157888
rect 176292 157836 176344 157888
rect 185860 157836 185912 157888
rect 186044 157836 186096 157888
rect 186320 157836 186372 157888
rect 195520 157836 195572 157888
rect 171784 157768 171836 157820
rect 177672 157768 177724 157820
rect 181996 157768 182048 157820
rect 124864 157700 124916 157752
rect 160744 157700 160796 157752
rect 163044 157700 163096 157752
rect 165804 157700 165856 157752
rect 166080 157700 166132 157752
rect 167184 157700 167236 157752
rect 184388 157700 184440 157752
rect 186044 157700 186096 157752
rect 192116 157768 192168 157820
rect 194140 157768 194192 157820
rect 195152 157768 195204 157820
rect 197728 157768 197780 157820
rect 192208 157700 192260 157752
rect 194416 157700 194468 157752
rect 196808 157700 196860 157752
rect 160928 157632 160980 157684
rect 177120 157632 177172 157684
rect 181352 157632 181404 157684
rect 183284 157632 183336 157684
rect 184480 157632 184532 157684
rect 185768 157632 185820 157684
rect 187148 157632 187200 157684
rect 190460 157632 190512 157684
rect 191104 157632 191156 157684
rect 195428 157632 195480 157684
rect 199384 157632 199436 157684
rect 165068 157564 165120 157616
rect 202604 157904 202656 157956
rect 202788 157904 202840 157956
rect 207480 157972 207532 158024
rect 208492 157972 208544 158024
rect 253572 157972 253624 158024
rect 207020 157904 207072 157956
rect 221556 157904 221608 157956
rect 199568 157836 199620 157888
rect 207112 157836 207164 157888
rect 208216 157836 208268 157888
rect 260288 157768 260340 157820
rect 202144 157700 202196 157752
rect 210792 157700 210844 157752
rect 200948 157632 201000 157684
rect 209596 157632 209648 157684
rect 152924 157292 152976 157344
rect 163412 157496 163464 157548
rect 164332 157496 164384 157548
rect 164884 157496 164936 157548
rect 165620 157496 165672 157548
rect 198280 157496 198332 157548
rect 158628 157428 158680 157480
rect 166080 157428 166132 157480
rect 170404 157428 170456 157480
rect 171048 157428 171100 157480
rect 210884 157564 210936 157616
rect 205640 157496 205692 157548
rect 205824 157496 205876 157548
rect 207204 157496 207256 157548
rect 214932 157496 214984 157548
rect 161020 157360 161072 157412
rect 164056 157360 164108 157412
rect 162768 157292 162820 157344
rect 163044 157292 163096 157344
rect 163504 157292 163556 157344
rect 170128 157292 170180 157344
rect 154304 157224 154356 157276
rect 159640 157156 159692 157208
rect 161848 157156 161900 157208
rect 162124 157224 162176 157276
rect 166540 157224 166592 157276
rect 169944 157224 169996 157276
rect 171048 157224 171100 157276
rect 163412 157156 163464 157208
rect 163964 157156 164016 157208
rect 164884 157156 164936 157208
rect 211068 157360 211120 157412
rect 187976 157292 188028 157344
rect 208400 157292 208452 157344
rect 190736 157224 190788 157276
rect 200948 157224 201000 157276
rect 202236 157224 202288 157276
rect 202788 157224 202840 157276
rect 190184 157156 190236 157208
rect 191656 157156 191708 157208
rect 192392 157156 192444 157208
rect 206192 157156 206244 157208
rect 160744 157088 160796 157140
rect 171600 157088 171652 157140
rect 183100 157088 183152 157140
rect 242164 157088 242216 157140
rect 143540 157020 143592 157072
rect 173532 157020 173584 157072
rect 213184 157020 213236 157072
rect 130384 156952 130436 157004
rect 161480 156952 161532 157004
rect 99380 156884 99432 156936
rect 163504 156952 163556 157004
rect 163596 156952 163648 157004
rect 164148 156952 164200 157004
rect 165804 156952 165856 157004
rect 166172 156952 166224 157004
rect 170496 156952 170548 157004
rect 171048 156952 171100 157004
rect 179052 156952 179104 157004
rect 213920 156952 213972 157004
rect 161848 156884 161900 156936
rect 165620 156884 165672 156936
rect 166632 156884 166684 156936
rect 196256 156884 196308 156936
rect 202236 156884 202288 156936
rect 205824 156884 205876 156936
rect 239864 156884 239916 156936
rect 85580 156816 85632 156868
rect 169024 156816 169076 156868
rect 179604 156816 179656 156868
rect 200672 156816 200724 156868
rect 200948 156816 201000 156868
rect 209228 156816 209280 156868
rect 81440 156748 81492 156800
rect 168656 156748 168708 156800
rect 178776 156748 178828 156800
rect 209688 156748 209740 156800
rect 215852 156748 215904 156800
rect 74540 156680 74592 156732
rect 168196 156680 168248 156732
rect 67640 156612 67692 156664
rect 167644 156612 167696 156664
rect 182548 156680 182600 156732
rect 191380 156680 191432 156732
rect 220360 156680 220412 156732
rect 220268 156612 220320 156664
rect 245016 156612 245068 156664
rect 267004 156612 267056 156664
rect 161480 156544 161532 156596
rect 169944 156544 169996 156596
rect 176568 156544 176620 156596
rect 176844 156544 176896 156596
rect 185768 156544 185820 156596
rect 191380 156544 191432 156596
rect 200672 156544 200724 156596
rect 211804 156544 211856 156596
rect 212356 156544 212408 156596
rect 154212 156476 154264 156528
rect 164240 156476 164292 156528
rect 165252 156476 165304 156528
rect 185400 156476 185452 156528
rect 275928 156476 275980 156528
rect 289176 156612 289228 156664
rect 159548 156408 159600 156460
rect 167000 156408 167052 156460
rect 168012 156408 168064 156460
rect 169668 156408 169720 156460
rect 170680 156408 170732 156460
rect 172980 156408 173032 156460
rect 232964 156408 233016 156460
rect 175372 156340 175424 156392
rect 176384 156340 176436 156392
rect 235172 156340 235224 156392
rect 184112 156272 184164 156324
rect 207020 156272 207072 156324
rect 176292 156068 176344 156120
rect 179420 156068 179472 156120
rect 191012 156000 191064 156052
rect 191196 156000 191248 156052
rect 164424 155932 164476 155984
rect 165528 155932 165580 155984
rect 189908 155932 189960 155984
rect 191380 155932 191432 155984
rect 149060 155864 149112 155916
rect 150348 155864 150400 155916
rect 164700 155864 164752 155916
rect 193588 155864 193640 155916
rect 195888 155864 195940 155916
rect 206376 155932 206428 155984
rect 206928 155932 206980 155984
rect 269764 155932 269816 155984
rect 518900 155932 518952 155984
rect 272156 155864 272208 155916
rect 272340 155864 272392 155916
rect 125600 155592 125652 155644
rect 159824 155592 159876 155644
rect 171968 155796 172020 155848
rect 185492 155796 185544 155848
rect 191012 155796 191064 155848
rect 196992 155796 197044 155848
rect 203064 155796 203116 155848
rect 271236 155796 271288 155848
rect 271788 155796 271840 155848
rect 164700 155728 164752 155780
rect 165344 155728 165396 155780
rect 190276 155728 190328 155780
rect 214840 155728 214892 155780
rect 200672 155660 200724 155712
rect 207204 155660 207256 155712
rect 168564 155592 168616 155644
rect 175372 155592 175424 155644
rect 180156 155592 180208 155644
rect 222108 155592 222160 155644
rect 225604 155592 225656 155644
rect 137284 155524 137336 155576
rect 172796 155524 172848 155576
rect 175188 155524 175240 155576
rect 216128 155524 216180 155576
rect 115204 155456 115256 155508
rect 150440 155456 150492 155508
rect 175372 155456 175424 155508
rect 175740 155456 175792 155508
rect 216036 155456 216088 155508
rect 135260 155388 135312 155440
rect 172980 155388 173032 155440
rect 179328 155388 179380 155440
rect 210424 155388 210476 155440
rect 106280 155320 106332 155372
rect 169760 155320 169812 155372
rect 191012 155320 191064 155372
rect 207848 155320 207900 155372
rect 272340 155320 272392 155372
rect 355324 155320 355376 155372
rect 26240 155252 26292 155304
rect 149060 155252 149112 155304
rect 150440 155252 150492 155304
rect 174176 155252 174228 155304
rect 177948 155252 178000 155304
rect 193588 155252 193640 155304
rect 270224 155252 270276 155304
rect 494060 155252 494112 155304
rect 13084 155184 13136 155236
rect 152924 155184 152976 155236
rect 178040 155184 178092 155236
rect 191012 155184 191064 155236
rect 271788 155184 271840 155236
rect 522304 155184 522356 155236
rect 193036 155116 193088 155168
rect 200672 155116 200724 155168
rect 201684 155116 201736 155168
rect 202696 155116 202748 155168
rect 267924 155116 267976 155168
rect 179880 155048 179932 155100
rect 212448 155048 212500 155100
rect 213184 155048 213236 155100
rect 174176 154980 174228 155032
rect 234436 154980 234488 155032
rect 185860 154912 185912 154964
rect 207940 154912 207992 154964
rect 184664 154844 184716 154896
rect 190276 154844 190328 154896
rect 190920 154844 190972 154896
rect 208032 154844 208084 154896
rect 191012 154708 191064 154760
rect 201960 154708 202012 154760
rect 200580 154640 200632 154692
rect 203064 154640 203116 154692
rect 174728 154572 174780 154624
rect 175188 154572 175240 154624
rect 194508 154572 194560 154624
rect 200672 154572 200724 154624
rect 201224 154504 201276 154556
rect 215116 154504 215168 154556
rect 196532 154436 196584 154488
rect 210700 154436 210752 154488
rect 188436 154368 188488 154420
rect 249248 154368 249300 154420
rect 181628 154300 181680 154352
rect 240784 154300 240836 154352
rect 157064 154232 157116 154284
rect 160192 154232 160244 154284
rect 174912 154232 174964 154284
rect 183836 154232 183888 154284
rect 243544 154232 243596 154284
rect 153200 154164 153252 154216
rect 173348 154164 173400 154216
rect 176292 154164 176344 154216
rect 182916 154164 182968 154216
rect 151820 154096 151872 154148
rect 174268 154096 174320 154148
rect 180432 154096 180484 154148
rect 227812 154096 227864 154148
rect 139400 153960 139452 154012
rect 173256 154028 173308 154080
rect 217324 154028 217376 154080
rect 180524 153960 180576 154012
rect 220728 153960 220780 154012
rect 228364 153960 228416 154012
rect 91100 153892 91152 153944
rect 169484 153892 169536 153944
rect 46940 153824 46992 153876
rect 155776 153824 155828 153876
rect 157340 153824 157392 153876
rect 174636 153892 174688 153944
rect 213000 153892 213052 153944
rect 178868 153824 178920 153876
rect 211160 153824 211212 153876
rect 212172 153824 212224 153876
rect 269120 154096 269172 154148
rect 270040 154096 270092 154148
rect 287244 154096 287296 154148
rect 288348 154096 288400 154148
rect 241336 153824 241388 153876
rect 253204 153824 253256 153876
rect 178592 153756 178644 153808
rect 208400 153756 208452 153808
rect 209412 153756 209464 153808
rect 176292 153620 176344 153672
rect 236000 153620 236052 153672
rect 191196 153552 191248 153604
rect 252192 153552 252244 153604
rect 270040 153280 270092 153332
rect 483020 153280 483072 153332
rect 195612 153212 195664 153264
rect 200580 153212 200632 153264
rect 204352 153212 204404 153264
rect 204628 153212 204680 153264
rect 205364 153212 205416 153264
rect 205548 153212 205600 153264
rect 227812 153212 227864 153264
rect 228916 153212 228968 153264
rect 229744 153212 229796 153264
rect 288348 153212 288400 153264
rect 507860 153212 507912 153264
rect 181904 153144 181956 153196
rect 182088 153144 182140 153196
rect 204444 153144 204496 153196
rect 273812 153144 273864 153196
rect 276480 153144 276532 153196
rect 579896 153144 579948 153196
rect 186504 153076 186556 153128
rect 280252 153076 280304 153128
rect 281448 153076 281500 153128
rect 202328 153008 202380 153060
rect 269028 153008 269080 153060
rect 178684 152940 178736 152992
rect 183284 152940 183336 152992
rect 189264 152940 189316 152992
rect 190184 152940 190236 152992
rect 190552 152940 190604 152992
rect 191564 152940 191616 152992
rect 196072 152940 196124 152992
rect 196532 152940 196584 152992
rect 199016 152940 199068 152992
rect 258632 152940 258684 152992
rect 182364 152872 182416 152924
rect 241428 152872 241480 152924
rect 246304 152872 246356 152924
rect 181812 152804 181864 152856
rect 239404 152804 239456 152856
rect 180984 152736 181036 152788
rect 185492 152736 185544 152788
rect 173164 152668 173216 152720
rect 173808 152668 173860 152720
rect 187148 152736 187200 152788
rect 193036 152736 193088 152788
rect 193312 152736 193364 152788
rect 193956 152736 194008 152788
rect 194876 152736 194928 152788
rect 247316 152736 247368 152788
rect 214564 152668 214616 152720
rect 217324 152668 217376 152720
rect 217784 152668 217836 152720
rect 133880 152600 133932 152652
rect 129004 152532 129056 152584
rect 34520 152464 34572 152516
rect 149152 152464 149204 152516
rect 168656 152600 168708 152652
rect 169208 152600 169260 152652
rect 177672 152600 177724 152652
rect 182916 152600 182968 152652
rect 185492 152600 185544 152652
rect 281448 152600 281500 152652
rect 307208 152600 307260 152652
rect 171140 152532 171192 152584
rect 172336 152532 172388 152584
rect 182456 152532 182508 152584
rect 183192 152532 183244 152584
rect 183284 152532 183336 152584
rect 167276 152464 167328 152516
rect 167644 152464 167696 152516
rect 171692 152464 171744 152516
rect 171876 152464 171928 152516
rect 175556 152464 175608 152516
rect 176200 152464 176252 152516
rect 176844 152464 176896 152516
rect 177580 152464 177632 152516
rect 182272 152464 182324 152516
rect 182824 152464 182876 152516
rect 185124 152464 185176 152516
rect 185952 152464 186004 152516
rect 186596 152532 186648 152584
rect 187056 152532 187108 152584
rect 187700 152532 187752 152584
rect 188712 152532 188764 152584
rect 189172 152532 189224 152584
rect 189816 152532 189868 152584
rect 190552 152532 190604 152584
rect 191472 152532 191524 152584
rect 191932 152532 191984 152584
rect 192576 152532 192628 152584
rect 193220 152532 193272 152584
rect 194232 152532 194284 152584
rect 194692 152532 194744 152584
rect 195060 152532 195112 152584
rect 195152 152532 195204 152584
rect 212908 152532 212960 152584
rect 269028 152532 269080 152584
rect 512000 152532 512052 152584
rect 209872 152464 209924 152516
rect 273812 152464 273864 152516
rect 274548 152464 274600 152516
rect 536104 152464 536156 152516
rect 167460 152396 167512 152448
rect 167920 152396 167972 152448
rect 168380 152396 168432 152448
rect 169116 152396 169168 152448
rect 172980 152396 173032 152448
rect 173624 152396 173676 152448
rect 175464 152396 175516 152448
rect 176476 152396 176528 152448
rect 172796 152328 172848 152380
rect 220084 152396 220136 152448
rect 181168 152328 181220 152380
rect 181996 152328 182048 152380
rect 182364 152328 182416 152380
rect 183468 152328 183520 152380
rect 185308 152328 185360 152380
rect 186136 152328 186188 152380
rect 186504 152328 186556 152380
rect 187332 152328 187384 152380
rect 188344 152328 188396 152380
rect 188896 152328 188948 152380
rect 192024 152328 192076 152380
rect 192852 152328 192904 152380
rect 193036 152328 193088 152380
rect 210608 152328 210660 152380
rect 172244 152260 172296 152312
rect 210516 152260 210568 152312
rect 185032 152192 185084 152244
rect 186228 152192 186280 152244
rect 186412 152192 186464 152244
rect 187608 152192 187660 152244
rect 191840 152192 191892 152244
rect 192944 152192 192996 152244
rect 194968 152192 195020 152244
rect 195888 152192 195940 152244
rect 196072 152192 196124 152244
rect 196716 152192 196768 152244
rect 197360 152192 197412 152244
rect 198096 152192 198148 152244
rect 198832 152192 198884 152244
rect 199936 152192 199988 152244
rect 200212 152192 200264 152244
rect 200764 152192 200816 152244
rect 201684 152192 201736 152244
rect 202512 152192 202564 152244
rect 203340 152192 203392 152244
rect 203800 152192 203852 152244
rect 204812 152192 204864 152244
rect 205456 152192 205508 152244
rect 188896 152124 188948 152176
rect 195152 152124 195204 152176
rect 196256 152124 196308 152176
rect 196900 152124 196952 152176
rect 197452 152124 197504 152176
rect 198556 152124 198608 152176
rect 202880 152124 202932 152176
rect 203892 152124 203944 152176
rect 165988 151852 166040 151904
rect 166264 151852 166316 151904
rect 176660 151716 176712 151768
rect 181536 151716 181588 151768
rect 189632 151716 189684 151768
rect 190092 151716 190144 151768
rect 203064 151716 203116 151768
rect 280160 151716 280212 151768
rect 182640 151648 182692 151700
rect 244924 151648 244976 151700
rect 174544 151580 174596 151632
rect 175648 151580 175700 151632
rect 235540 151580 235592 151632
rect 185676 151512 185728 151564
rect 242808 151512 242860 151564
rect 181076 151444 181128 151496
rect 236644 151444 236696 151496
rect 181260 151376 181312 151428
rect 232504 151376 232556 151428
rect 180248 151308 180300 151360
rect 229100 151308 229152 151360
rect 230020 151308 230072 151360
rect 140780 151240 140832 151292
rect 158444 151240 158496 151292
rect 184940 151240 184992 151292
rect 233976 151240 234028 151292
rect 82820 151172 82872 151224
rect 152832 151172 152884 151224
rect 189080 151172 189132 151224
rect 189540 151172 189592 151224
rect 192208 151172 192260 151224
rect 240876 151172 240928 151224
rect 64880 151104 64932 151156
rect 155500 151104 155552 151156
rect 189448 151104 189500 151156
rect 190000 151104 190052 151156
rect 198004 151104 198056 151156
rect 242992 151104 243044 151156
rect 29000 151036 29052 151088
rect 164516 151036 164568 151088
rect 189080 151036 189132 151088
rect 190368 151036 190420 151088
rect 197084 151036 197136 151088
rect 236000 151036 236052 151088
rect 242808 151036 242860 151088
rect 295984 151036 296036 151088
rect 195520 150968 195572 151020
rect 233240 150968 233292 151020
rect 199660 150900 199712 150952
rect 223212 150900 223264 150952
rect 190092 150832 190144 150884
rect 211620 150832 211672 150884
rect 233240 150492 233292 150544
rect 234252 150492 234304 150544
rect 236000 150424 236052 150476
rect 236920 150424 236972 150476
rect 244924 150424 244976 150476
rect 250444 150424 250496 150476
rect 280160 150424 280212 150476
rect 280804 150424 280856 150476
rect 3332 150356 3384 150408
rect 11704 150356 11756 150408
rect 186688 150356 186740 150408
rect 215944 150356 215996 150408
rect 204260 150288 204312 150340
rect 291292 150288 291344 150340
rect 187792 150220 187844 150272
rect 272524 150220 272576 150272
rect 187424 150152 187476 150204
rect 259460 150152 259512 150204
rect 175004 150084 175056 150136
rect 235448 150084 235500 150136
rect 197636 150016 197688 150068
rect 257436 150016 257488 150068
rect 196624 149948 196676 150000
rect 252100 149948 252152 150000
rect 181628 149880 181680 149932
rect 235264 149880 235316 149932
rect 177488 149812 177540 149864
rect 218704 149812 218756 149864
rect 56600 149744 56652 149796
rect 165712 149744 165764 149796
rect 179144 149744 179196 149796
rect 213736 149744 213788 149796
rect 215944 149744 215996 149796
rect 234068 149744 234120 149796
rect 272524 149744 272576 149796
rect 327080 149744 327132 149796
rect 15200 149676 15252 149728
rect 163136 149676 163188 149728
rect 186688 149676 186740 149728
rect 186964 149676 187016 149728
rect 201960 149676 202012 149728
rect 232872 149676 232924 149728
rect 291292 149676 291344 149728
rect 451280 149676 451332 149728
rect 188528 149608 188580 149660
rect 217508 149608 217560 149660
rect 184020 149540 184072 149592
rect 274824 149540 274876 149592
rect 172520 149472 172572 149524
rect 175832 149472 175884 149524
rect 214012 149472 214064 149524
rect 187792 149268 187844 149320
rect 188988 149268 189040 149320
rect 213736 149064 213788 149116
rect 214564 149064 214616 149116
rect 259460 149064 259512 149116
rect 260104 149064 260156 149116
rect 274824 149064 274876 149116
rect 275284 149064 275336 149116
rect 181904 148996 181956 149048
rect 217140 148996 217192 149048
rect 220084 148996 220136 149048
rect 183560 148928 183612 148980
rect 271880 148928 271932 148980
rect 186044 148860 186096 148912
rect 267832 148860 267884 148912
rect 268384 148860 268436 148912
rect 182180 148792 182232 148844
rect 243728 148792 243780 148844
rect 184296 148724 184348 148776
rect 244096 148724 244148 148776
rect 182180 148656 182232 148708
rect 182548 148656 182600 148708
rect 184480 148656 184532 148708
rect 243636 148656 243688 148708
rect 194140 148588 194192 148640
rect 252008 148588 252060 148640
rect 191656 148520 191708 148572
rect 246396 148520 246448 148572
rect 189724 148452 189776 148504
rect 244280 148452 244332 148504
rect 271880 148452 271932 148504
rect 272432 148452 272484 148504
rect 144920 148384 144972 148436
rect 173716 148384 173768 148436
rect 202236 148384 202288 148436
rect 256056 148384 256108 148436
rect 57980 148316 58032 148368
rect 165896 148316 165948 148368
rect 192668 148316 192720 148368
rect 237012 148316 237064 148368
rect 244096 148316 244148 148368
rect 278044 148316 278096 148368
rect 191564 148248 191616 148300
rect 230204 148248 230256 148300
rect 179512 148180 179564 148232
rect 215300 148180 215352 148232
rect 190184 148112 190236 148164
rect 278412 148112 278464 148164
rect 345020 148316 345072 148368
rect 244280 147636 244332 147688
rect 244924 147636 244976 147688
rect 200856 147568 200908 147620
rect 228548 147568 228600 147620
rect 201776 147500 201828 147552
rect 287244 147500 287296 147552
rect 194784 147432 194836 147484
rect 278964 147432 279016 147484
rect 279976 147432 280028 147484
rect 182456 147364 182508 147416
rect 260196 147364 260248 147416
rect 264244 147364 264296 147416
rect 168380 147296 168432 147348
rect 168564 147296 168616 147348
rect 184756 147296 184808 147348
rect 245200 147296 245252 147348
rect 185308 147228 185360 147280
rect 246580 147228 246632 147280
rect 190736 147160 190788 147212
rect 251916 147160 251968 147212
rect 188068 147092 188120 147144
rect 247684 147092 247736 147144
rect 153844 147024 153896 147076
rect 175096 147024 175148 147076
rect 196348 147024 196400 147076
rect 255412 147024 255464 147076
rect 126244 146956 126296 147008
rect 161756 146956 161808 147008
rect 191104 146956 191156 147008
rect 250536 146956 250588 147008
rect 104900 146888 104952 146940
rect 170956 146888 171008 146940
rect 189540 146888 189592 146940
rect 235816 146888 235868 146940
rect 179696 146820 179748 146872
rect 222200 146820 222252 146872
rect 223028 146820 223080 146872
rect 215300 146752 215352 146804
rect 216588 146752 216640 146804
rect 239588 146752 239640 146804
rect 187976 146684 188028 146736
rect 276204 146684 276256 146736
rect 316684 146956 316736 147008
rect 279976 146888 280028 146940
rect 415400 146888 415452 146940
rect 177396 146276 177448 146328
rect 180064 146276 180116 146328
rect 201684 146208 201736 146260
rect 294052 146208 294104 146260
rect 294880 146208 294932 146260
rect 183652 146140 183704 146192
rect 245476 146140 245528 146192
rect 282184 146140 282236 146192
rect 189448 146072 189500 146124
rect 251088 146072 251140 146124
rect 190644 146004 190696 146056
rect 250996 146004 251048 146056
rect 195336 145936 195388 145988
rect 253388 145936 253440 145988
rect 196716 145868 196768 145920
rect 254860 145868 254912 145920
rect 197728 145800 197780 145852
rect 254952 145800 255004 145852
rect 199384 145732 199436 145784
rect 255964 145732 256016 145784
rect 251088 145664 251140 145716
rect 356060 145664 356112 145716
rect 138020 145596 138072 145648
rect 172888 145596 172940 145648
rect 250996 145596 251048 145648
rect 369860 145596 369912 145648
rect 46204 145528 46256 145580
rect 152464 145528 152516 145580
rect 155960 145528 156012 145580
rect 174820 145528 174872 145580
rect 202420 145528 202472 145580
rect 257344 145528 257396 145580
rect 294880 145528 294932 145580
rect 514024 145528 514076 145580
rect 170036 145460 170088 145512
rect 170496 145460 170548 145512
rect 222844 145460 222896 145512
rect 200488 145392 200540 145444
rect 251824 145392 251876 145444
rect 199476 145324 199528 145376
rect 226984 145324 227036 145376
rect 200948 145256 201000 145308
rect 254768 145256 254820 145308
rect 200764 145188 200816 145240
rect 254676 145188 254728 145240
rect 196164 144848 196216 144900
rect 289268 144848 289320 144900
rect 289728 144848 289780 144900
rect 185124 144780 185176 144832
rect 278136 144780 278188 144832
rect 284944 144780 284996 144832
rect 189356 144712 189408 144764
rect 274640 144712 274692 144764
rect 175556 144644 175608 144696
rect 176568 144644 176620 144696
rect 202880 144644 202932 144696
rect 270316 144644 270368 144696
rect 198832 144576 198884 144628
rect 260380 144576 260432 144628
rect 175464 144508 175516 144560
rect 176476 144508 176528 144560
rect 238116 144508 238168 144560
rect 196256 144440 196308 144492
rect 257528 144440 257580 144492
rect 176844 144372 176896 144424
rect 177948 144372 178000 144424
rect 185216 144372 185268 144424
rect 245108 144372 245160 144424
rect 205824 144304 205876 144356
rect 206652 144304 206704 144356
rect 265440 144304 265492 144356
rect 274640 144304 274692 144356
rect 341524 144304 341576 144356
rect 142160 144236 142212 144288
rect 173440 144236 173492 144288
rect 177764 144236 177816 144288
rect 231124 144236 231176 144288
rect 289728 144236 289780 144288
rect 436744 144236 436796 144288
rect 75920 144168 75972 144220
rect 167000 144168 167052 144220
rect 176476 144168 176528 144220
rect 225788 144168 225840 144220
rect 270316 144168 270368 144220
rect 532700 144168 532752 144220
rect 176568 143964 176620 144016
rect 222936 144100 222988 144152
rect 177028 143556 177080 143608
rect 177764 143556 177816 143608
rect 193312 143488 193364 143540
rect 288532 143488 288584 143540
rect 186780 143420 186832 143472
rect 277584 143420 277636 143472
rect 278688 143420 278740 143472
rect 197544 143352 197596 143404
rect 282920 143352 282972 143404
rect 193956 143284 194008 143336
rect 273260 143284 273312 143336
rect 203800 143216 203852 143268
rect 271144 143216 271196 143268
rect 182364 143148 182416 143200
rect 244188 143148 244240 143200
rect 177856 143080 177908 143132
rect 220176 143080 220228 143132
rect 204444 143012 204496 143064
rect 205272 143012 205324 143064
rect 118700 142944 118752 142996
rect 172152 142944 172204 142996
rect 174636 142944 174688 142996
rect 224224 142944 224276 142996
rect 60832 142876 60884 142928
rect 167368 142876 167420 142928
rect 177304 142876 177356 142928
rect 177856 142876 177908 142928
rect 35900 142808 35952 142860
rect 164240 142808 164292 142860
rect 176752 142808 176804 142860
rect 179328 142808 179380 142860
rect 229836 142876 229888 142928
rect 278688 142944 278740 142996
rect 309876 142944 309928 142996
rect 261484 142876 261536 142928
rect 273260 142876 273312 142928
rect 380900 142876 380952 142928
rect 205272 142808 205324 142860
rect 263600 142808 263652 142860
rect 282920 142808 282972 142860
rect 283748 142808 283800 142860
rect 449900 142808 449952 142860
rect 202696 142128 202748 142180
rect 260840 142128 260892 142180
rect 193220 142060 193272 142112
rect 285864 142060 285916 142112
rect 194692 141992 194744 142044
rect 287520 141992 287572 142044
rect 198464 141924 198516 141976
rect 287796 141924 287848 141976
rect 204904 141856 204956 141908
rect 267740 141856 267792 141908
rect 269028 141856 269080 141908
rect 185032 141788 185084 141840
rect 246948 141788 247000 141840
rect 164424 141720 164476 141772
rect 223856 141720 223908 141772
rect 188988 141652 189040 141704
rect 225880 141652 225932 141704
rect 189264 141584 189316 141636
rect 190368 141584 190420 141636
rect 227076 141584 227128 141636
rect 246948 141584 247000 141636
rect 302884 141584 302936 141636
rect 287520 141516 287572 141568
rect 419540 141516 419592 141568
rect 92480 141448 92532 141500
rect 168932 141448 168984 141500
rect 187792 141448 187844 141500
rect 323584 141448 323636 141500
rect 48320 141380 48372 141432
rect 165804 141380 165856 141432
rect 187884 141380 187936 141432
rect 188988 141380 189040 141432
rect 269028 141380 269080 141432
rect 550640 141380 550692 141432
rect 285864 140768 285916 140820
rect 286324 140768 286376 140820
rect 182272 140700 182324 140752
rect 183376 140700 183428 140752
rect 186596 140700 186648 140752
rect 281540 140700 281592 140752
rect 197360 140632 197412 140684
rect 261576 140632 261628 140684
rect 198648 140564 198700 140616
rect 258816 140564 258868 140616
rect 183376 140496 183428 140548
rect 241796 140496 241848 140548
rect 191656 140428 191708 140480
rect 231216 140428 231268 140480
rect 190000 140360 190052 140412
rect 225972 140360 226024 140412
rect 281540 140088 281592 140140
rect 314016 140088 314068 140140
rect 20720 140020 20772 140072
rect 162860 140020 162912 140072
rect 280804 140020 280856 140072
rect 363604 140020 363656 140072
rect 186504 139340 186556 139392
rect 282276 139340 282328 139392
rect 192116 139272 192168 139324
rect 284392 139272 284444 139324
rect 184848 139204 184900 139256
rect 244740 139204 244792 139256
rect 249064 139204 249116 139256
rect 167276 139136 167328 139188
rect 167644 139136 167696 139188
rect 227720 139136 227772 139188
rect 166448 139068 166500 139120
rect 225696 139068 225748 139120
rect 168564 139000 168616 139052
rect 169116 139000 169168 139052
rect 228456 139000 228508 139052
rect 122840 138728 122892 138780
rect 171692 138728 171744 138780
rect 282276 138728 282328 138780
rect 320180 138728 320232 138780
rect 40040 138660 40092 138712
rect 164424 138660 164476 138712
rect 284392 138660 284444 138712
rect 383660 138660 383712 138712
rect 3056 137912 3108 137964
rect 159364 137912 159416 137964
rect 187700 137912 187752 137964
rect 282920 137912 282972 137964
rect 205180 137844 205232 137896
rect 272708 137844 272760 137896
rect 167736 137776 167788 137828
rect 168012 137776 168064 137828
rect 223764 137776 223816 137828
rect 282920 137368 282972 137420
rect 283564 137368 283616 137420
rect 338120 137368 338172 137420
rect 288532 137300 288584 137352
rect 405740 137300 405792 137352
rect 146300 137232 146352 137284
rect 173164 137232 173216 137284
rect 180616 137232 180668 137284
rect 219440 137232 219492 137284
rect 272708 137232 272760 137284
rect 554780 137232 554832 137284
rect 205732 136552 205784 136604
rect 272248 136552 272300 136604
rect 196072 136484 196124 136536
rect 255872 136484 255924 136536
rect 189172 136416 189224 136468
rect 247316 136416 247368 136468
rect 79324 135940 79376 135992
rect 168564 135940 168616 135992
rect 247316 135940 247368 135992
rect 248236 135940 248288 135992
rect 351920 135940 351972 135992
rect 55220 135872 55272 135924
rect 166448 135872 166500 135924
rect 255872 135872 255924 135924
rect 256608 135872 256660 135924
rect 440240 135872 440292 135924
rect 272248 135260 272300 135312
rect 568580 135260 568632 135312
rect 206376 135192 206428 135244
rect 270500 135192 270552 135244
rect 271788 135192 271840 135244
rect 190552 135124 190604 135176
rect 249708 135124 249760 135176
rect 249708 134648 249760 134700
rect 351184 134648 351236 134700
rect 287796 134580 287848 134632
rect 455420 134580 455472 134632
rect 18604 134512 18656 134564
rect 161664 134512 161716 134564
rect 181996 134512 182048 134564
rect 241520 134512 241572 134564
rect 271788 134512 271840 134564
rect 549904 134512 549956 134564
rect 192024 133832 192076 133884
rect 252468 133832 252520 133884
rect 102140 133220 102192 133272
rect 169852 133220 169904 133272
rect 252468 133220 252520 133272
rect 390560 133220 390612 133272
rect 8300 133152 8352 133204
rect 163688 133152 163740 133204
rect 208124 133152 208176 133204
rect 575480 133152 575532 133204
rect 191932 132404 191984 132456
rect 287152 132404 287204 132456
rect 288348 132404 288400 132456
rect 186412 132336 186464 132388
rect 248328 132336 248380 132388
rect 248328 131792 248380 131844
rect 287704 131792 287756 131844
rect 111800 131724 111852 131776
rect 172336 131724 172388 131776
rect 288348 131724 288400 131776
rect 387800 131724 387852 131776
rect 84200 130364 84252 130416
rect 169208 130364 169260 130416
rect 286324 130364 286376 130416
rect 408500 130364 408552 130416
rect 199844 129684 199896 129736
rect 270408 129684 270460 129736
rect 195612 129616 195664 129668
rect 253848 129616 253900 129668
rect 98000 129072 98052 129124
rect 170496 129072 170548 129124
rect 253848 129072 253900 129124
rect 422944 129072 422996 129124
rect 25504 129004 25556 129056
rect 163044 129004 163096 129056
rect 182088 129004 182140 129056
rect 237380 129004 237432 129056
rect 270408 129004 270460 129056
rect 480260 129004 480312 129056
rect 189080 128256 189132 128308
rect 284300 128256 284352 128308
rect 195980 128188 196032 128240
rect 291200 128188 291252 128240
rect 291660 128188 291712 128240
rect 117320 127644 117372 127696
rect 171416 127644 171468 127696
rect 284300 127644 284352 127696
rect 358820 127644 358872 127696
rect 66260 127576 66312 127628
rect 167644 127576 167696 127628
rect 291660 127576 291712 127628
rect 444380 127576 444432 127628
rect 200120 126896 200172 126948
rect 273904 126896 273956 126948
rect 274088 126896 274140 126948
rect 261576 126284 261628 126336
rect 458180 126284 458232 126336
rect 69020 126216 69072 126268
rect 167828 126216 167880 126268
rect 274088 126216 274140 126268
rect 489920 126216 489972 126268
rect 190460 125536 190512 125588
rect 285772 125536 285824 125588
rect 286232 125536 286284 125588
rect 115940 124924 115992 124976
rect 171324 124924 171376 124976
rect 15844 124856 15896 124908
rect 162952 124856 163004 124908
rect 286232 124856 286284 124908
rect 376760 124856 376812 124908
rect 201592 124108 201644 124160
rect 294512 124108 294564 124160
rect 111064 123496 111116 123548
rect 170772 123496 170824 123548
rect 191840 123496 191892 123548
rect 394700 123496 394752 123548
rect 14464 123428 14516 123480
rect 161572 123428 161624 123480
rect 294512 123428 294564 123480
rect 503720 123428 503772 123480
rect 86960 122068 87012 122120
rect 169024 122068 169076 122120
rect 203892 122068 203944 122120
rect 520924 122068 520976 122120
rect 23480 120708 23532 120760
rect 164608 120708 164660 120760
rect 205272 120708 205324 120760
rect 539692 120708 539744 120760
rect 19340 119348 19392 119400
rect 161020 119348 161072 119400
rect 22744 117920 22796 117972
rect 163412 117920 163464 117972
rect 163504 117920 163556 117972
rect 174820 117920 174872 117972
rect 187516 116628 187568 116680
rect 307852 116628 307904 116680
rect 22100 116560 22152 116612
rect 163596 116560 163648 116612
rect 198556 116560 198608 116612
rect 462320 116560 462372 116612
rect 39304 115200 39356 115252
rect 164700 115200 164752 115252
rect 166356 112412 166408 112464
rect 174084 112412 174136 112464
rect 194416 112412 194468 112464
rect 404360 112412 404412 112464
rect 3332 111732 3384 111784
rect 142804 111732 142856 111784
rect 183376 111052 183428 111104
rect 262220 111052 262272 111104
rect 9680 109692 9732 109744
rect 163320 109692 163372 109744
rect 49700 108264 49752 108316
rect 166080 108264 166132 108316
rect 178040 108264 178092 108316
rect 200764 108264 200816 108316
rect 201316 108264 201368 108316
rect 492680 108264 492732 108316
rect 63500 106904 63552 106956
rect 167552 106904 167604 106956
rect 167644 106904 167696 106956
rect 174728 106904 174780 106956
rect 70400 105544 70452 105596
rect 167460 105544 167512 105596
rect 201408 105544 201460 105596
rect 499580 105544 499632 105596
rect 88340 104116 88392 104168
rect 168748 104116 168800 104168
rect 177672 104116 177724 104168
rect 189724 104116 189776 104168
rect 190368 104116 190420 104168
rect 347780 104116 347832 104168
rect 102232 102756 102284 102808
rect 171048 102756 171100 102808
rect 202696 102756 202748 102808
rect 510620 102756 510672 102808
rect 120080 101396 120132 101448
rect 171876 101396 171928 101448
rect 337384 100648 337436 100700
rect 580172 100648 580224 100700
rect 31760 99968 31812 100020
rect 164976 99968 165028 100020
rect 176476 99288 176528 99340
rect 180800 99288 180852 99340
rect 27620 98608 27672 98660
rect 158352 98608 158404 98660
rect 53840 97316 53892 97368
rect 165620 97316 165672 97368
rect 161940 97248 161992 97300
rect 580264 97248 580316 97300
rect 11704 95888 11756 95940
rect 163228 95888 163280 95940
rect 183468 94528 183520 94580
rect 269120 94528 269172 94580
rect 42800 94460 42852 94512
rect 148324 94460 148376 94512
rect 203984 94460 204036 94512
rect 535460 94460 535512 94512
rect 180708 93168 180760 93220
rect 234712 93168 234764 93220
rect 204352 93100 204404 93152
rect 542360 93100 542412 93152
rect 205456 91740 205508 91792
rect 546500 91740 546552 91792
rect 206652 88952 206704 89004
rect 552664 88952 552716 89004
rect 205548 87592 205600 87644
rect 553400 87592 553452 87644
rect 206560 86232 206612 86284
rect 560300 86232 560352 86284
rect 208216 83444 208268 83496
rect 574100 83444 574152 83496
rect 206836 82084 206888 82136
rect 567200 82084 567252 82136
rect 208308 80656 208360 80708
rect 578240 80656 578292 80708
rect 194508 79296 194560 79348
rect 400220 79296 400272 79348
rect 162032 73788 162084 73840
rect 580264 73788 580316 73840
rect 188896 72428 188948 72480
rect 331864 72428 331916 72480
rect 3516 71680 3568 71732
rect 120724 71680 120776 71732
rect 177764 66852 177816 66904
rect 187700 66852 187752 66904
rect 95976 59984 96028 60036
rect 170588 59984 170640 60036
rect 177856 59984 177908 60036
rect 191104 59984 191156 60036
rect 3056 59304 3108 59356
rect 95884 59304 95936 59356
rect 3516 45500 3568 45552
rect 155224 45500 155276 45552
rect 75184 37884 75236 37936
rect 167736 37884 167788 37936
rect 204076 36524 204128 36576
rect 525800 36524 525852 36576
rect 179236 33736 179288 33788
rect 205640 33736 205692 33788
rect 206928 33736 206980 33788
rect 564532 33736 564584 33788
rect 2872 33056 2924 33108
rect 43444 33056 43496 33108
rect 280068 33056 280120 33108
rect 580172 33056 580224 33108
rect 203616 28228 203668 28280
rect 524420 28228 524472 28280
rect 175924 23468 175976 23520
rect 176660 23468 176712 23520
rect 187608 22720 187660 22772
rect 315396 22720 315448 22772
rect 334624 20612 334676 20664
rect 580080 20612 580132 20664
rect 202788 17212 202840 17264
rect 505100 17212 505152 17264
rect 39120 15852 39172 15904
rect 164792 15852 164844 15904
rect 177948 15852 178000 15904
rect 195152 15852 195204 15904
rect 195796 15852 195848 15904
rect 429200 15852 429252 15904
rect 11152 14424 11204 14476
rect 124864 14424 124916 14476
rect 25320 13064 25372 13116
rect 164884 13064 164936 13116
rect 197452 13064 197504 13116
rect 465172 13064 465224 13116
rect 160100 11772 160152 11824
rect 161296 11772 161348 11824
rect 46112 11704 46164 11756
rect 166264 11704 166316 11756
rect 198740 11704 198792 11756
rect 478880 11704 478932 11756
rect 35992 10276 36044 10328
rect 151084 10276 151136 10328
rect 200028 10276 200080 10328
rect 472256 10276 472308 10328
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 193128 8984 193180 9036
rect 383568 8984 383620 9036
rect 110512 8916 110564 8968
rect 170404 8916 170456 8968
rect 195888 8916 195940 8968
rect 418988 8916 419040 8968
rect 176568 8236 176620 8288
rect 177856 8236 177908 8288
rect 78588 7556 78640 7608
rect 168472 7556 168524 7608
rect 3424 6808 3476 6860
rect 146944 6808 146996 6860
rect 191748 6264 191800 6316
rect 369400 6264 369452 6316
rect 191656 6196 191708 6248
rect 372896 6196 372948 6248
rect 197268 6128 197320 6180
rect 436652 6128 436704 6180
rect 19432 4768 19484 4820
rect 156604 4768 156656 4820
rect 188988 4768 189040 4820
rect 330392 4768 330444 4820
rect 315304 4156 315356 4208
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 149520 4088 149572 4140
rect 153844 4088 153896 4140
rect 209688 4088 209740 4140
rect 210976 4088 211028 4140
rect 243728 4088 243780 4140
rect 254676 4088 254728 4140
rect 275284 4088 275336 4140
rect 278320 4088 278372 4140
rect 315396 4088 315448 4140
rect 316040 4088 316092 4140
rect 171416 4020 171468 4072
rect 171784 4020 171836 4072
rect 193864 4020 193916 4072
rect 200304 4020 200356 4072
rect 240876 4020 240928 4072
rect 251180 4020 251232 4072
rect 314016 4020 314068 4072
rect 316684 4088 316736 4140
rect 323676 4088 323728 4140
rect 571984 4088 572036 4140
rect 577412 4088 577464 4140
rect 239404 3952 239456 4004
rect 249984 3952 250036 4004
rect 250444 3952 250496 4004
rect 260656 3952 260708 4004
rect 313188 3952 313240 4004
rect 326804 4020 326856 4072
rect 507124 4020 507176 4072
rect 510068 4020 510120 4072
rect 235264 3884 235316 3936
rect 246396 3884 246448 3936
rect 246580 3884 246632 3936
rect 257068 3884 257120 3936
rect 264244 3884 264296 3936
rect 267740 3884 267792 3936
rect 302884 3884 302936 3936
rect 306748 3884 306800 3936
rect 317328 3952 317380 4004
rect 325608 3952 325660 4004
rect 431224 3952 431276 4004
rect 434444 3952 434496 4004
rect 323676 3884 323728 3936
rect 331588 3884 331640 3936
rect 363604 3884 363656 3936
rect 367008 3884 367060 3936
rect 44272 3816 44324 3868
rect 46204 3816 46256 3868
rect 244924 3816 244976 3868
rect 258264 3816 258316 3868
rect 261484 3816 261536 3868
rect 271236 3816 271288 3868
rect 305644 3816 305696 3868
rect 314016 3816 314068 3868
rect 323584 3816 323636 3868
rect 342168 3816 342220 3868
rect 179328 3748 179380 3800
rect 184940 3748 184992 3800
rect 213184 3748 213236 3800
rect 225144 3748 225196 3800
rect 236644 3748 236696 3800
rect 240508 3748 240560 3800
rect 242164 3748 242216 3800
rect 265348 3748 265400 3800
rect 268384 3748 268436 3800
rect 283104 3748 283156 3800
rect 307116 3748 307168 3800
rect 329196 3748 329248 3800
rect 118792 3680 118844 3732
rect 127624 3680 127676 3732
rect 189816 3680 189868 3732
rect 194416 3680 194468 3732
rect 211804 3680 211856 3732
rect 221556 3680 221608 3732
rect 228364 3680 228416 3732
rect 235816 3680 235868 3732
rect 243636 3680 243688 3732
rect 268844 3680 268896 3732
rect 284944 3680 284996 3732
rect 303160 3680 303212 3732
rect 308404 3680 308456 3732
rect 332600 3680 332652 3732
rect 374092 3680 374144 3732
rect 375288 3680 375340 3732
rect 376024 3680 376076 3732
rect 398840 3680 398892 3732
rect 6460 3612 6512 3664
rect 11704 3612 11756 3664
rect 1676 3544 1728 3596
rect 14464 3612 14516 3664
rect 14740 3612 14792 3664
rect 25504 3612 25556 3664
rect 96252 3612 96304 3664
rect 130384 3612 130436 3664
rect 180156 3612 180208 3664
rect 190828 3612 190880 3664
rect 13544 3544 13596 3596
rect 15844 3544 15896 3596
rect 60740 3544 60792 3596
rect 61660 3544 61712 3596
rect 69112 3544 69164 3596
rect 71044 3544 71096 3596
rect 86868 3544 86920 3596
rect 88984 3544 89036 3596
rect 95148 3544 95200 3596
rect 95976 3544 96028 3596
rect 110420 3544 110472 3596
rect 111616 3544 111668 3596
rect 114008 3544 114060 3596
rect 115204 3544 115256 3596
rect 118700 3544 118752 3596
rect 119896 3544 119948 3596
rect 124680 3544 124732 3596
rect 160744 3544 160796 3596
rect 162768 3544 162820 3596
rect 166080 3544 166132 3596
rect 180064 3544 180116 3596
rect 182916 3544 182968 3596
rect 196808 3612 196860 3664
rect 220084 3612 220136 3664
rect 4068 3476 4120 3528
rect 18604 3476 18656 3528
rect 31300 3476 31352 3528
rect 32404 3476 32456 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 38384 3476 38436 3528
rect 39304 3476 39356 3528
rect 53748 3476 53800 3528
rect 162124 3476 162176 3528
rect 162492 3476 162544 3528
rect 163504 3476 163556 3528
rect 164884 3476 164936 3528
rect 167644 3476 167696 3528
rect 170772 3476 170824 3528
rect 174636 3476 174688 3528
rect 193220 3544 193272 3596
rect 225604 3544 225656 3596
rect 228732 3544 228784 3596
rect 232504 3612 232556 3664
rect 242900 3612 242952 3664
rect 243544 3612 243596 3664
rect 276020 3612 276072 3664
rect 287704 3612 287756 3664
rect 324412 3612 324464 3664
rect 327724 3612 327776 3664
rect 339868 3612 339920 3664
rect 341524 3612 341576 3664
rect 349160 3612 349212 3664
rect 355324 3612 355376 3664
rect 402520 3612 402572 3664
rect 423772 3612 423824 3664
rect 424968 3612 425020 3664
rect 448612 3612 448664 3664
rect 449808 3612 449860 3664
rect 552664 3612 552716 3664
rect 557356 3612 557408 3664
rect 253480 3544 253532 3596
rect 253572 3544 253624 3596
rect 260012 3544 260064 3596
rect 260104 3544 260156 3596
rect 261760 3544 261812 3596
rect 265624 3544 265676 3596
rect 266544 3544 266596 3596
rect 267004 3544 267056 3596
rect 292580 3544 292632 3596
rect 295984 3544 296036 3596
rect 299664 3544 299716 3596
rect 307852 3544 307904 3596
rect 309048 3544 309100 3596
rect 191104 3476 191156 3528
rect 192024 3476 192076 3528
rect 198004 3476 198056 3528
rect 199108 3476 199160 3528
rect 217324 3476 217376 3528
rect 239312 3476 239364 3528
rect 240784 3476 240836 3528
rect 247592 3476 247644 3528
rect 249064 3476 249116 3528
rect 288992 3476 289044 3528
rect 289084 3476 289136 3528
rect 290188 3476 290240 3528
rect 305736 3476 305788 3528
rect 311440 3544 311492 3596
rect 320824 3544 320876 3596
rect 346952 3544 347004 3596
rect 349252 3544 349304 3596
rect 350448 3544 350500 3596
rect 351276 3544 351328 3596
rect 374092 3544 374144 3596
rect 378048 3544 378100 3596
rect 463976 3544 464028 3596
rect 471244 3544 471296 3596
rect 474556 3544 474608 3596
rect 547880 3544 547932 3596
rect 548708 3544 548760 3596
rect 549904 3544 549956 3596
rect 572720 3544 572772 3596
rect 311164 3476 311216 3528
rect 312636 3476 312688 3528
rect 313924 3476 313976 3528
rect 2872 3408 2924 3460
rect 126244 3408 126296 3460
rect 126980 3408 127032 3460
rect 128176 3408 128228 3460
rect 135260 3408 135312 3460
rect 136456 3408 136508 3460
rect 169576 3408 169628 3460
rect 174544 3408 174596 3460
rect 181536 3408 181588 3460
rect 183744 3408 183796 3460
rect 109316 3340 109368 3392
rect 111064 3340 111116 3392
rect 182824 3340 182876 3392
rect 207388 3408 207440 3460
rect 210424 3408 210476 3460
rect 218060 3408 218112 3460
rect 215944 3340 215996 3392
rect 258724 3340 258776 3392
rect 259460 3340 259512 3392
rect 260012 3340 260064 3392
rect 264152 3340 264204 3392
rect 271144 3340 271196 3392
rect 274824 3340 274876 3392
rect 278044 3340 278096 3392
rect 281908 3340 281960 3392
rect 309876 3340 309928 3392
rect 313832 3340 313884 3392
rect 18236 3272 18288 3324
rect 22744 3272 22796 3324
rect 77392 3272 77444 3324
rect 79324 3272 79376 3324
rect 126980 3272 127032 3324
rect 129004 3272 129056 3324
rect 135260 3272 135312 3324
rect 137284 3272 137336 3324
rect 214564 3272 214616 3324
rect 215668 3272 215720 3324
rect 309784 3272 309836 3324
rect 320824 3340 320876 3392
rect 332692 3340 332744 3392
rect 333888 3340 333940 3392
rect 357532 3408 357584 3460
rect 358728 3408 358780 3460
rect 390560 3408 390612 3460
rect 391848 3408 391900 3460
rect 363512 3340 363564 3392
rect 387064 3340 387116 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 415400 3476 415452 3528
rect 416688 3476 416740 3528
rect 422944 3476 422996 3528
rect 423772 3476 423824 3528
rect 432052 3476 432104 3528
rect 433248 3476 433300 3528
rect 436744 3476 436796 3528
rect 437940 3476 437992 3528
rect 440240 3476 440292 3528
rect 441528 3476 441580 3528
rect 447784 3476 447836 3528
rect 448612 3476 448664 3528
rect 456892 3476 456944 3528
rect 458088 3476 458140 3528
rect 465080 3476 465132 3528
rect 465908 3476 465960 3528
rect 468484 3476 468536 3528
rect 469864 3476 469916 3528
rect 472624 3476 472676 3528
rect 473452 3476 473504 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 520924 3476 520976 3528
rect 521844 3476 521896 3528
rect 522304 3476 522356 3528
rect 523040 3476 523092 3528
rect 527916 3476 527968 3528
rect 552664 3476 552716 3528
rect 421380 3340 421432 3392
rect 566832 3408 566884 3460
rect 27712 3204 27764 3256
rect 31024 3204 31076 3256
rect 163688 3204 163740 3256
rect 166356 3204 166408 3256
rect 175280 3204 175332 3256
rect 179052 3204 179104 3256
rect 314016 3204 314068 3256
rect 318524 3204 318576 3256
rect 216588 3136 216640 3188
rect 219256 3136 219308 3188
rect 282184 3136 282236 3188
rect 285404 3136 285456 3188
rect 307208 3136 307260 3188
rect 310244 3136 310296 3188
rect 331864 3136 331916 3188
rect 335084 3136 335136 3188
rect 12348 3068 12400 3120
rect 13084 3068 13136 3120
rect 229744 3068 229796 3120
rect 232228 3068 232280 3120
rect 247684 3068 247736 3120
rect 248788 3068 248840 3120
rect 543004 3068 543056 3120
rect 545488 3068 545540 3120
rect 41880 3000 41932 3052
rect 44824 3000 44876 3052
rect 167184 3000 167236 3052
rect 171416 3000 171468 3052
rect 181444 3000 181496 3052
rect 189724 3000 189776 3052
rect 196624 3000 196676 3052
rect 197912 3000 197964 3052
rect 200764 3000 200816 3052
rect 202696 3000 202748 3052
rect 289176 3000 289228 3052
rect 296076 3000 296128 3052
rect 307024 3000 307076 3052
rect 315028 3000 315080 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 536196 3000 536248 3052
rect 540796 3000 540848 3052
rect 291844 2932 291896 2984
rect 293684 2932 293736 2984
rect 548524 2932 548576 2984
rect 550272 2932 550324 2984
rect 115204 2864 115256 2916
rect 116584 2864 116636 2916
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3436 402286 3464 566879
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 4816 413914 4844 553794
rect 6932 450537 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 10324 656940 10376 656946
rect 10324 656882 10376 656888
rect 6918 450528 6974 450537
rect 6918 450463 6974 450472
rect 8944 448588 8996 448594
rect 8944 448530 8996 448536
rect 8956 416770 8984 448530
rect 8944 416764 8996 416770
rect 8944 416706 8996 416712
rect 4804 413908 4856 413914
rect 4804 413850 4856 413856
rect 10336 410582 10364 656882
rect 40052 467158 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 51724 501016 51776 501022
rect 51724 500958 51776 500964
rect 40040 467152 40092 467158
rect 40040 467094 40092 467100
rect 51736 414730 51764 500958
rect 51724 414724 51776 414730
rect 51724 414666 51776 414672
rect 10324 410576 10376 410582
rect 4066 410544 4122 410553
rect 4122 410502 4200 410530
rect 10324 410518 10376 410524
rect 4066 410479 4122 410488
rect 4172 405686 4200 410502
rect 4160 405680 4212 405686
rect 4160 405622 4212 405628
rect 71792 404297 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 406434 88380 702406
rect 104912 465730 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 104900 465724 104952 465730
rect 104900 465666 104952 465672
rect 136652 450566 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 136640 450560 136692 450566
rect 136640 450502 136692 450508
rect 88340 406428 88392 406434
rect 88340 406370 88392 406376
rect 71778 404288 71834 404297
rect 71778 404223 71834 404232
rect 3424 402280 3476 402286
rect 3424 402222 3476 402228
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 385694 3464 397423
rect 3424 385688 3476 385694
rect 3424 385630 3476 385636
rect 153212 373998 153240 702406
rect 169772 464370 169800 702406
rect 180064 605872 180116 605878
rect 180064 605814 180116 605820
rect 169760 464364 169812 464370
rect 169760 464306 169812 464312
rect 180076 411942 180104 605814
rect 201512 450634 201540 702986
rect 218992 699718 219020 703520
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 220084 699712 220136 699718
rect 220084 699654 220136 699660
rect 201500 450628 201552 450634
rect 201500 450570 201552 450576
rect 180064 411936 180116 411942
rect 180064 411878 180116 411884
rect 220096 374678 220124 699654
rect 234632 461650 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700330 283880 703520
rect 280804 700324 280856 700330
rect 280804 700266 280856 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 262864 514820 262916 514826
rect 262864 514762 262916 514768
rect 234620 461644 234672 461650
rect 234620 461586 234672 461592
rect 262876 417450 262904 514762
rect 266372 450702 266400 697546
rect 273260 465724 273312 465730
rect 273260 465666 273312 465672
rect 273272 465118 273300 465666
rect 273260 465112 273312 465118
rect 273260 465054 273312 465060
rect 274548 465112 274600 465118
rect 274548 465054 274600 465060
rect 266360 450696 266412 450702
rect 266360 450638 266412 450644
rect 262864 417444 262916 417450
rect 262864 417386 262916 417392
rect 265806 402112 265862 402121
rect 265806 402047 265862 402056
rect 263322 401840 263378 401849
rect 263322 401775 263378 401784
rect 260748 398268 260800 398274
rect 260748 398210 260800 398216
rect 256606 398168 256662 398177
rect 256606 398103 256662 398112
rect 257988 398132 258040 398138
rect 255320 385688 255372 385694
rect 255320 385630 255372 385636
rect 255332 385082 255360 385630
rect 255320 385076 255372 385082
rect 255320 385018 255372 385024
rect 253204 382424 253256 382430
rect 253204 382366 253256 382372
rect 246304 380996 246356 381002
rect 246304 380938 246356 380944
rect 243544 379636 243596 379642
rect 243544 379578 243596 379584
rect 232504 375828 232556 375834
rect 232504 375770 232556 375776
rect 220728 375420 220780 375426
rect 220728 375362 220780 375368
rect 220084 374672 220136 374678
rect 220084 374614 220136 374620
rect 153200 373992 153252 373998
rect 153200 373934 153252 373940
rect 220450 373280 220506 373289
rect 220360 373244 220412 373250
rect 220450 373215 220506 373224
rect 220360 373186 220412 373192
rect 219900 372632 219952 372638
rect 219900 372574 219952 372580
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 209688 322312 209740 322318
rect 209688 322254 209740 322260
rect 204166 322144 204222 322153
rect 204166 322079 204222 322088
rect 204076 321632 204128 321638
rect 204076 321574 204128 321580
rect 3424 319456 3476 319462
rect 3424 319398 3476 319404
rect 3436 319297 3464 319398
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 202696 312792 202748 312798
rect 202696 312734 202748 312740
rect 4066 306232 4122 306241
rect 4122 306190 4200 306218
rect 4066 306167 4122 306176
rect 4172 298858 4200 306190
rect 201408 303680 201460 303686
rect 201408 303622 201460 303628
rect 200120 302252 200172 302258
rect 200120 302194 200172 302200
rect 197360 300960 197412 300966
rect 197360 300902 197412 300908
rect 195980 299668 196032 299674
rect 195980 299610 196032 299616
rect 4160 298852 4212 298858
rect 4160 298794 4212 298800
rect 194600 298172 194652 298178
rect 194600 298114 194652 298120
rect 179420 297220 179472 297226
rect 179420 297162 179472 297168
rect 173900 297084 173952 297090
rect 173900 297026 173952 297032
rect 169760 295928 169812 295934
rect 169760 295870 169812 295876
rect 167000 294704 167052 294710
rect 167000 294646 167052 294652
rect 164516 294636 164568 294642
rect 164516 294578 164568 294584
rect 162676 293276 162728 293282
rect 162676 293218 162728 293224
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 14464 266416 14516 266422
rect 14464 266358 14516 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 14476 241466 14504 266358
rect 158626 241768 158682 241777
rect 158626 241703 158682 241712
rect 151726 241632 151782 241641
rect 151726 241567 151782 241576
rect 157248 241596 157300 241602
rect 14464 241460 14516 241466
rect 14464 241402 14516 241408
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 239426 3372 241023
rect 3332 239420 3384 239426
rect 3332 239362 3384 239368
rect 150348 236768 150400 236774
rect 150348 236710 150400 236716
rect 150254 228440 150310 228449
rect 150254 228375 150310 228384
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 11704 211812 11756 211818
rect 11704 211754 11756 211760
rect 3424 210656 3476 210662
rect 3424 210598 3476 210604
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3056 137964 3108 137970
rect 3056 137906 3108 137912
rect 3068 136785 3096 137906
rect 3054 136776 3110 136785
rect 3054 136711 3110 136720
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 19417 3464 210598
rect 3608 210588 3660 210594
rect 3608 210530 3660 210536
rect 3516 210520 3568 210526
rect 3516 210462 3568 210468
rect 3528 84697 3556 210462
rect 3620 97617 3648 210530
rect 3700 210452 3752 210458
rect 3700 210394 3752 210400
rect 3712 162897 3740 210394
rect 3698 162888 3754 162897
rect 3698 162823 3754 162832
rect 4160 158024 4212 158030
rect 4160 157966 4212 157972
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 157966
rect 6918 153776 6974 153785
rect 6918 153711 6974 153720
rect 6932 16574 6960 153711
rect 11716 150414 11744 211754
rect 95884 211540 95936 211546
rect 95884 211482 95936 211488
rect 43444 209092 43496 209098
rect 43444 209034 43496 209040
rect 26240 155304 26292 155310
rect 26240 155246 26292 155252
rect 13084 155236 13136 155242
rect 13084 155178 13136 155184
rect 11704 150408 11756 150414
rect 11704 150350 11756 150356
rect 8300 133204 8352 133210
rect 8300 133146 8352 133152
rect 8312 16574 8340 133146
rect 9680 109744 9732 109750
rect 9680 109686 9732 109692
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 480 1716 3538
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2884 480 2912 3402
rect 4080 480 4108 3470
rect 5276 480 5304 16546
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 480 6500 3606
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 109686
rect 11704 95940 11756 95946
rect 11704 95882 11756 95888
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11164 480 11192 14418
rect 11716 3670 11744 95882
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 13096 3126 13124 155178
rect 15200 149728 15252 149734
rect 15200 149670 15252 149676
rect 14464 123480 14516 123486
rect 14464 123422 14516 123428
rect 14476 3670 14504 123422
rect 15212 16574 15240 149670
rect 16578 146976 16634 146985
rect 16578 146911 16634 146920
rect 15844 124908 15896 124914
rect 15844 124850 15896 124856
rect 15212 16546 15792 16574
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 12360 480 12388 3062
rect 13556 480 13584 3538
rect 14752 480 14780 3606
rect 15764 3482 15792 16546
rect 15856 3602 15884 124850
rect 16592 16574 16620 146911
rect 20720 140072 20772 140078
rect 20720 140014 20772 140020
rect 18604 134564 18656 134570
rect 18604 134506 18656 134512
rect 16592 16546 17080 16574
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15764 3454 15976 3482
rect 15948 480 15976 3454
rect 17052 480 17080 16546
rect 18616 3534 18644 134506
rect 19340 119400 19392 119406
rect 19340 119342 19392 119348
rect 19352 16574 19380 119342
rect 20732 16574 20760 140014
rect 25504 129056 25556 129062
rect 25504 128998 25556 129004
rect 23480 120760 23532 120766
rect 23480 120702 23532 120708
rect 22744 117972 22796 117978
rect 22744 117914 22796 117920
rect 22100 116612 22152 116618
rect 22100 116554 22152 116560
rect 22112 16574 22140 116554
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18236 3324 18288 3330
rect 18236 3266 18288 3272
rect 18248 480 18276 3266
rect 19444 480 19472 4762
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 3330 22784 117914
rect 23492 16574 23520 120702
rect 23492 16546 24256 16574
rect 22744 3324 22796 3330
rect 22744 3266 22796 3272
rect 24228 480 24256 16546
rect 25320 13116 25372 13122
rect 25320 13058 25372 13064
rect 25332 480 25360 13058
rect 25516 3670 25544 128998
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 155246
rect 34520 152516 34572 152522
rect 34520 152458 34572 152464
rect 29000 151088 29052 151094
rect 29000 151030 29052 151036
rect 27620 98660 27672 98666
rect 27620 98602 27672 98608
rect 27632 16574 27660 98602
rect 29012 16574 29040 151030
rect 31022 148336 31078 148345
rect 31022 148271 31078 148280
rect 27632 16546 28488 16574
rect 29012 16546 30144 16574
rect 27712 3256 27764 3262
rect 27712 3198 27764 3204
rect 27724 480 27752 3198
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 31036 3262 31064 148271
rect 33138 144120 33194 144129
rect 33138 144055 33194 144064
rect 32402 130384 32458 130393
rect 32402 130319 32458 130328
rect 31760 100020 31812 100026
rect 31760 99962 31812 99968
rect 31772 16574 31800 99962
rect 31772 16546 31984 16574
rect 31300 3528 31352 3534
rect 31300 3470 31352 3476
rect 31024 3256 31076 3262
rect 31024 3198 31076 3204
rect 31312 480 31340 3470
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 32416 3534 32444 130319
rect 33152 16574 33180 144055
rect 33152 16546 33640 16574
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 152458
rect 35900 142860 35952 142866
rect 35900 142802 35952 142808
rect 35912 3534 35940 142802
rect 40040 138712 40092 138718
rect 40040 138654 40092 138660
rect 39304 115252 39356 115258
rect 39304 115194 39356 115200
rect 39120 15904 39172 15910
rect 39120 15846 39172 15852
rect 35992 10328 36044 10334
rect 35992 10270 36044 10276
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 10270
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 3470
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 15846
rect 39316 3534 39344 115194
rect 40052 16574 40080 138654
rect 42800 94512 42852 94518
rect 42800 94454 42852 94460
rect 40052 16546 40264 16574
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 3052 41932 3058
rect 41880 2994 41932 3000
rect 41892 480 41920 2994
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 94454
rect 43456 33114 43484 209034
rect 78680 158160 78732 158166
rect 78680 158102 78732 158108
rect 60740 158092 60792 158098
rect 60740 158034 60792 158040
rect 46940 153876 46992 153882
rect 46940 153818 46992 153824
rect 46204 145580 46256 145586
rect 46204 145522 46256 145528
rect 44822 113792 44878 113801
rect 44822 113727 44878 113736
rect 44178 112432 44234 112441
rect 44178 112367 44234 112376
rect 43444 33108 43496 33114
rect 43444 33050 43496 33056
rect 44192 16574 44220 112367
rect 44192 16546 44772 16574
rect 44272 3868 44324 3874
rect 44272 3810 44324 3816
rect 44284 480 44312 3810
rect 44744 490 44772 16546
rect 44836 3058 44864 113727
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 46124 3482 46152 11698
rect 46216 3874 46244 145522
rect 46952 16574 46980 153818
rect 51078 152416 51134 152425
rect 51078 152351 51134 152360
rect 48320 141432 48372 141438
rect 48320 141374 48372 141380
rect 48332 16574 48360 141374
rect 49700 108316 49752 108322
rect 49700 108258 49752 108264
rect 49712 16574 49740 108258
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 3868 46256 3874
rect 46204 3810 46256 3816
rect 46124 3454 46704 3482
rect 44824 3052 44876 3058
rect 44824 2994 44876 3000
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 44744 462 45140 490
rect 46676 480 46704 3454
rect 45112 354 45140 462
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 152351
rect 56600 149796 56652 149802
rect 56600 149738 56652 149744
rect 55220 135924 55272 135930
rect 55220 135866 55272 135872
rect 52458 131744 52514 131753
rect 52458 131679 52514 131688
rect 52472 16574 52500 131679
rect 53840 97368 53892 97374
rect 53840 97310 53892 97316
rect 53852 16574 53880 97310
rect 55232 16574 55260 135866
rect 56612 16574 56640 149738
rect 57980 148368 58032 148374
rect 57980 148310 58032 148316
rect 57992 16574 58020 148310
rect 59358 137320 59414 137329
rect 59358 137255 59414 137264
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52564 480 52592 16546
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 53760 480 53788 3470
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 137255
rect 60752 3602 60780 158034
rect 74540 156732 74592 156738
rect 74540 156674 74592 156680
rect 67640 156664 67692 156670
rect 67640 156606 67692 156612
rect 64880 151156 64932 151162
rect 64880 151098 64932 151104
rect 60832 142928 60884 142934
rect 60832 142870 60884 142876
rect 60740 3596 60792 3602
rect 60740 3538 60792 3544
rect 60844 480 60872 142870
rect 62118 138680 62174 138689
rect 62118 138615 62174 138624
rect 62132 16574 62160 138615
rect 63500 106956 63552 106962
rect 63500 106898 63552 106904
rect 63512 16574 63540 106898
rect 64892 16574 64920 151098
rect 66260 127628 66312 127634
rect 66260 127570 66312 127576
rect 66272 16574 66300 127570
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3596 61712 3602
rect 61660 3538 61712 3544
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3538
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 156606
rect 71778 153912 71834 153921
rect 71778 153847 71834 153856
rect 71042 149696 71098 149705
rect 71042 149631 71098 149640
rect 69020 126268 69072 126274
rect 69020 126210 69072 126216
rect 69032 16574 69060 126210
rect 70400 105596 70452 105602
rect 70400 105538 70452 105544
rect 70412 16574 70440 105538
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69124 480 69152 3538
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3602 71084 149631
rect 71792 16574 71820 153847
rect 74552 16574 74580 156674
rect 75920 144220 75972 144226
rect 75920 144162 75972 144168
rect 75184 37936 75236 37942
rect 75184 37878 75236 37884
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 37878
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 144162
rect 78692 16574 78720 158102
rect 85580 156868 85632 156874
rect 85580 156810 85632 156816
rect 81440 156800 81492 156806
rect 81440 156742 81492 156748
rect 80058 140040 80114 140049
rect 80058 139975 80114 139984
rect 79324 135992 79376 135998
rect 79324 135934 79376 135940
rect 78692 16546 79272 16574
rect 78588 7608 78640 7614
rect 78588 7550 78640 7556
rect 77392 3324 77444 3330
rect 77392 3266 77444 3272
rect 77404 480 77432 3266
rect 78600 480 78628 7550
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 79336 3330 79364 135934
rect 80072 16574 80100 139975
rect 81452 16574 81480 156742
rect 82820 151224 82872 151230
rect 82820 151166 82872 151172
rect 82832 16574 82860 151166
rect 84200 130416 84252 130422
rect 84200 130358 84252 130364
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 79324 3324 79376 3330
rect 79324 3266 79376 3272
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 130358
rect 85592 16574 85620 156810
rect 91100 153944 91152 153950
rect 91100 153886 91152 153892
rect 89718 147112 89774 147121
rect 89718 147047 89774 147056
rect 88982 145616 89038 145625
rect 88982 145551 89038 145560
rect 86960 122120 87012 122126
rect 86960 122062 87012 122068
rect 86972 16574 87000 122062
rect 88340 104168 88392 104174
rect 88340 104110 88392 104116
rect 88352 16574 88380 104110
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 88352 16546 88932 16574
rect 85684 480 85712 16546
rect 86868 3596 86920 3602
rect 86868 3538 86920 3544
rect 86880 480 86908 3538
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 88904 3482 88932 16546
rect 88996 3602 89024 145551
rect 89732 16574 89760 147047
rect 91112 16574 91140 153886
rect 93858 145752 93914 145761
rect 93858 145687 93914 145696
rect 92480 141500 92532 141506
rect 92480 141442 92532 141448
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 88984 3596 89036 3602
rect 88984 3538 89036 3544
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 141442
rect 93872 16574 93900 145687
rect 95896 59362 95924 211482
rect 142804 209228 142856 209234
rect 142804 209170 142856 209176
rect 120724 209160 120776 209166
rect 120724 209102 120776 209108
rect 96620 159384 96672 159390
rect 96620 159326 96672 159332
rect 95976 60036 96028 60042
rect 95976 59978 96028 59984
rect 95884 59356 95936 59362
rect 95884 59298 95936 59304
rect 93872 16546 93992 16574
rect 93964 480 93992 16546
rect 95988 3602 96016 59978
rect 96632 16574 96660 159326
rect 99380 156936 99432 156942
rect 99380 156878 99432 156884
rect 98000 129124 98052 129130
rect 98000 129066 98052 129072
rect 98012 16574 98040 129066
rect 99392 16574 99420 156878
rect 115204 155508 115256 155514
rect 115204 155450 115256 155456
rect 106280 155372 106332 155378
rect 106280 155314 106332 155320
rect 100758 149832 100814 149841
rect 100758 149767 100814 149776
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 95148 3596 95200 3602
rect 95148 3538 95200 3544
rect 95976 3596 96028 3602
rect 95976 3538 96028 3544
rect 95160 480 95188 3538
rect 96264 480 96292 3606
rect 97460 480 97488 16546
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 149767
rect 103518 148472 103574 148481
rect 103518 148407 103574 148416
rect 102140 133272 102192 133278
rect 102140 133214 102192 133220
rect 102152 6914 102180 133214
rect 102232 102808 102284 102814
rect 102232 102750 102284 102756
rect 102244 16574 102272 102750
rect 103532 16574 103560 148407
rect 104900 146940 104952 146946
rect 104900 146882 104952 146888
rect 104912 16574 104940 146882
rect 106292 16574 106320 155314
rect 107658 144256 107714 144265
rect 107658 144191 107714 144200
rect 107672 16574 107700 144191
rect 110418 141400 110474 141409
rect 110418 141335 110474 141344
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 110432 3602 110460 141335
rect 111800 131776 111852 131782
rect 111800 131718 111852 131724
rect 111064 123548 111116 123554
rect 111064 123490 111116 123496
rect 110512 8968 110564 8974
rect 110512 8910 110564 8916
rect 110420 3596 110472 3602
rect 110420 3538 110472 3544
rect 109316 3392 109368 3398
rect 109316 3334 109368 3340
rect 109328 480 109356 3334
rect 110524 480 110552 8910
rect 111076 3398 111104 123490
rect 111812 16574 111840 131718
rect 111812 16546 112392 16574
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 111064 3392 111116 3398
rect 111064 3334 111116 3340
rect 111628 480 111656 3538
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 115216 3602 115244 155450
rect 116582 148608 116638 148617
rect 116582 148543 116638 148552
rect 115940 124976 115992 124982
rect 115940 124918 115992 124924
rect 115952 16574 115980 124918
rect 115952 16546 116440 16574
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 114020 480 114048 3538
rect 115204 2916 115256 2922
rect 115204 2858 115256 2864
rect 115216 480 115244 2858
rect 116412 480 116440 16546
rect 116596 2922 116624 148543
rect 118700 142996 118752 143002
rect 118700 142938 118752 142944
rect 117320 127696 117372 127702
rect 117320 127638 117372 127644
rect 116584 2916 116636 2922
rect 116584 2858 116636 2864
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 127638
rect 118712 3602 118740 142938
rect 120080 101448 120132 101454
rect 120080 101390 120132 101396
rect 120092 16574 120120 101390
rect 120736 71738 120764 209102
rect 132500 159520 132552 159526
rect 132500 159462 132552 159468
rect 128360 159452 128412 159458
rect 128360 159394 128412 159400
rect 124864 157752 124916 157758
rect 124864 157694 124916 157700
rect 121458 140176 121514 140185
rect 121458 140111 121514 140120
rect 120724 71732 120776 71738
rect 120724 71674 120776 71680
rect 121472 16574 121500 140111
rect 122840 138780 122892 138786
rect 122840 138722 122892 138728
rect 122852 16574 122880 138722
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 118792 3732 118844 3738
rect 118792 3674 118844 3680
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 118804 480 118832 3674
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 119908 480 119936 3538
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124876 14482 124904 157694
rect 125600 155644 125652 155650
rect 125600 155586 125652 155592
rect 124864 14476 124916 14482
rect 124864 14418 124916 14424
rect 124680 3596 124732 3602
rect 124680 3538 124732 3544
rect 124692 480 124720 3538
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 155586
rect 127622 149968 127678 149977
rect 127622 149903 127678 149912
rect 126244 147008 126296 147014
rect 126244 146950 126296 146956
rect 126256 3466 126284 146950
rect 126978 134464 127034 134473
rect 126978 134399 127034 134408
rect 126992 3466 127020 134399
rect 127636 3738 127664 149903
rect 128372 16574 128400 159394
rect 130384 157004 130436 157010
rect 130384 156946 130436 156952
rect 129004 152584 129056 152590
rect 129004 152526 129056 152532
rect 128372 16546 128952 16574
rect 127624 3732 127676 3738
rect 127624 3674 127676 3680
rect 126244 3460 126296 3466
rect 126244 3402 126296 3408
rect 126980 3460 127032 3466
rect 126980 3402 127032 3408
rect 128176 3460 128228 3466
rect 128176 3402 128228 3408
rect 126980 3324 127032 3330
rect 126980 3266 127032 3272
rect 126992 480 127020 3266
rect 128188 480 128216 3402
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 129016 3330 129044 152526
rect 129738 111072 129794 111081
rect 129738 111007 129794 111016
rect 129752 16574 129780 111007
rect 129752 16546 130332 16574
rect 130304 3482 130332 16546
rect 130396 3670 130424 156946
rect 131118 154048 131174 154057
rect 131118 153983 131174 153992
rect 131132 16574 131160 153983
rect 132512 16574 132540 159462
rect 137284 155576 137336 155582
rect 137284 155518 137336 155524
rect 135260 155440 135312 155446
rect 135260 155382 135312 155388
rect 133880 152652 133932 152658
rect 133880 152594 133932 152600
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 130384 3664 130436 3670
rect 130384 3606 130436 3612
rect 130304 3454 130608 3482
rect 129004 3324 129056 3330
rect 129004 3266 129056 3272
rect 130580 480 130608 3454
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 152594
rect 135272 3466 135300 155382
rect 136638 126304 136694 126313
rect 136638 126239 136694 126248
rect 136652 16574 136680 126239
rect 136652 16546 137232 16574
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 136456 3460 136508 3466
rect 136456 3402 136508 3408
rect 135260 3324 135312 3330
rect 135260 3266 135312 3272
rect 135272 480 135300 3266
rect 136468 480 136496 3402
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 3330 137324 155518
rect 139400 154012 139452 154018
rect 139400 153954 139452 153960
rect 138020 145648 138072 145654
rect 138020 145590 138072 145596
rect 138032 16574 138060 145590
rect 139412 16574 139440 153954
rect 140780 151292 140832 151298
rect 140780 151234 140832 151240
rect 140792 16574 140820 151234
rect 142160 144288 142212 144294
rect 142160 144230 142212 144236
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 137284 3324 137336 3330
rect 137284 3266 137336 3272
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 144230
rect 142816 111790 142844 209170
rect 146942 209128 146998 209137
rect 146942 209063 146998 209072
rect 143540 157072 143592 157078
rect 143540 157014 143592 157020
rect 142804 111784 142856 111790
rect 142804 111726 142856 111732
rect 143552 480 143580 157014
rect 144920 148436 144972 148442
rect 144920 148378 144972 148384
rect 143630 135960 143686 135969
rect 143630 135895 143686 135904
rect 143644 16574 143672 135895
rect 144932 16574 144960 148378
rect 146300 137284 146352 137290
rect 146300 137226 146352 137232
rect 146312 16574 146340 137226
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 146892 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146864 3482 146892 16546
rect 146956 6866 146984 209063
rect 150268 159089 150296 228375
rect 149150 159080 149206 159089
rect 149150 159015 149206 159024
rect 150254 159080 150310 159089
rect 150254 159015 150310 159024
rect 148324 157888 148376 157894
rect 148324 157830 148376 157836
rect 147678 141536 147734 141545
rect 147678 141471 147734 141480
rect 147692 16574 147720 141471
rect 148336 94518 148364 157830
rect 149060 155916 149112 155922
rect 149060 155858 149112 155864
rect 149072 155310 149100 155858
rect 149060 155304 149112 155310
rect 149060 155246 149112 155252
rect 149164 152522 149192 159015
rect 150360 155922 150388 236710
rect 151636 233912 151688 233918
rect 151636 233854 151688 233860
rect 151544 217320 151596 217326
rect 151544 217262 151596 217268
rect 151556 160177 151584 217262
rect 151174 160168 151230 160177
rect 151174 160103 151230 160112
rect 151542 160168 151598 160177
rect 151542 160103 151598 160112
rect 150438 158536 150494 158545
rect 150438 158471 150494 158480
rect 150348 155916 150400 155922
rect 150348 155858 150400 155864
rect 150452 155514 150480 158471
rect 151084 158364 151136 158370
rect 151084 158306 151136 158312
rect 150440 155508 150492 155514
rect 150440 155450 150492 155456
rect 150440 155304 150492 155310
rect 150440 155246 150492 155252
rect 149152 152516 149204 152522
rect 149152 152458 149204 152464
rect 148324 94512 148376 94518
rect 148324 94454 148376 94460
rect 150452 16574 150480 155246
rect 150530 140720 150586 140729
rect 150530 140655 150586 140664
rect 150544 140049 150572 140655
rect 150530 140040 150586 140049
rect 150530 139975 150586 139984
rect 147692 16546 147904 16574
rect 150452 16546 150664 16574
rect 146944 6860 146996 6866
rect 146944 6802 146996 6808
rect 146864 3454 147168 3482
rect 147140 480 147168 3454
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149520 4140 149572 4146
rect 149520 4082 149572 4088
rect 149532 480 149560 4082
rect 150636 480 150664 16546
rect 151096 10334 151124 158306
rect 151188 148345 151216 160103
rect 151648 158545 151676 233854
rect 151634 158536 151690 158545
rect 151634 158471 151690 158480
rect 151174 148336 151230 148345
rect 151174 148271 151230 148280
rect 151740 140729 151768 241567
rect 157248 241538 157300 241544
rect 154304 241528 154356 241534
rect 154304 241470 154356 241476
rect 154210 240272 154266 240281
rect 154210 240207 154266 240216
rect 153014 239456 153070 239465
rect 153014 239391 153070 239400
rect 152924 239284 152976 239290
rect 152924 239226 152976 239232
rect 152740 228812 152792 228818
rect 152740 228754 152792 228760
rect 152464 159928 152516 159934
rect 152464 159870 152516 159876
rect 151820 154148 151872 154154
rect 151820 154090 151872 154096
rect 151726 140720 151782 140729
rect 151726 140655 151782 140664
rect 151084 10328 151136 10334
rect 151084 10270 151136 10276
rect 151832 9674 151860 154090
rect 151910 150512 151966 150521
rect 151910 150447 151966 150456
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 150447
rect 152476 145586 152504 159870
rect 152752 159390 152780 228754
rect 152832 228540 152884 228546
rect 152832 228482 152884 228488
rect 152844 159934 152872 228482
rect 152832 159928 152884 159934
rect 152832 159870 152884 159876
rect 152936 159780 152964 239226
rect 152844 159752 152964 159780
rect 152844 159497 152872 159752
rect 153028 159712 153056 239391
rect 154120 239216 154172 239222
rect 154120 239158 154172 239164
rect 153108 234116 153160 234122
rect 153108 234058 153160 234064
rect 152936 159684 153056 159712
rect 152830 159488 152886 159497
rect 152830 159423 152886 159432
rect 152740 159384 152792 159390
rect 152740 159326 152792 159332
rect 152844 151230 152872 159423
rect 152936 157350 152964 159684
rect 153016 159588 153068 159594
rect 153016 159530 153068 159536
rect 153028 159390 153056 159530
rect 153016 159384 153068 159390
rect 153016 159326 153068 159332
rect 152924 157344 152976 157350
rect 152924 157286 152976 157292
rect 152936 155242 152964 157286
rect 152924 155236 152976 155242
rect 152924 155178 152976 155184
rect 152832 151224 152884 151230
rect 152832 151166 152884 151172
rect 153120 147665 153148 234058
rect 154028 228880 154080 228886
rect 154028 228822 154080 228828
rect 153936 213308 153988 213314
rect 153936 213250 153988 213256
rect 153948 159322 153976 213250
rect 153936 159316 153988 159322
rect 153936 159258 153988 159264
rect 154040 158953 154068 228822
rect 154132 159254 154160 239158
rect 154120 159248 154172 159254
rect 154120 159190 154172 159196
rect 154026 158944 154082 158953
rect 154026 158879 154082 158888
rect 153200 154216 153252 154222
rect 153200 154158 153252 154164
rect 153106 147656 153162 147665
rect 153106 147591 153162 147600
rect 152464 145580 152516 145586
rect 152464 145522 152516 145528
rect 153212 16574 153240 154158
rect 154040 149841 154068 158879
rect 154224 156534 154252 240207
rect 154316 157282 154344 241470
rect 155866 241088 155922 241097
rect 155866 241023 155922 241032
rect 154486 240952 154542 240961
rect 154486 240887 154542 240896
rect 154394 233064 154450 233073
rect 154394 232999 154450 233008
rect 154304 157276 154356 157282
rect 154304 157218 154356 157224
rect 154212 156528 154264 156534
rect 154212 156470 154264 156476
rect 154026 149832 154082 149841
rect 154026 149767 154082 149776
rect 153844 147076 153896 147082
rect 153844 147018 153896 147024
rect 153212 16546 153792 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 153856 4146 153884 147018
rect 154408 146305 154436 232999
rect 154394 146296 154450 146305
rect 154394 146231 154450 146240
rect 154500 146169 154528 240887
rect 155776 235340 155828 235346
rect 155776 235282 155828 235288
rect 155684 232620 155736 232626
rect 155684 232562 155736 232568
rect 155592 228676 155644 228682
rect 155592 228618 155644 228624
rect 155408 227044 155460 227050
rect 155408 226986 155460 226992
rect 155224 209840 155276 209846
rect 155224 209782 155276 209788
rect 154578 153096 154634 153105
rect 154578 153031 154634 153040
rect 154486 146160 154542 146169
rect 154486 146095 154542 146104
rect 154592 16574 154620 153031
rect 155236 45558 155264 209782
rect 155420 160313 155448 226986
rect 155500 222896 155552 222902
rect 155500 222838 155552 222844
rect 155406 160304 155462 160313
rect 155406 160239 155462 160248
rect 155314 158808 155370 158817
rect 155314 158743 155370 158752
rect 155328 149977 155356 158743
rect 155420 153785 155448 160239
rect 155512 156913 155540 222838
rect 155604 159050 155632 228618
rect 155696 159633 155724 232562
rect 155682 159624 155738 159633
rect 155682 159559 155738 159568
rect 155592 159044 155644 159050
rect 155592 158986 155644 158992
rect 155696 158817 155724 159559
rect 155682 158808 155738 158817
rect 155682 158743 155738 158752
rect 155788 157457 155816 235282
rect 155880 158817 155908 241023
rect 157154 239592 157210 239601
rect 157154 239527 157210 239536
rect 156972 233980 157024 233986
rect 156972 233922 157024 233928
rect 156880 232756 156932 232762
rect 156880 232698 156932 232704
rect 156788 225616 156840 225622
rect 156788 225558 156840 225564
rect 156696 214668 156748 214674
rect 156696 214610 156748 214616
rect 156604 211880 156656 211886
rect 156604 211822 156656 211828
rect 156616 202842 156644 211822
rect 156604 202836 156656 202842
rect 156604 202778 156656 202784
rect 156512 159656 156564 159662
rect 156512 159598 156564 159604
rect 155866 158808 155922 158817
rect 155866 158743 155922 158752
rect 155774 157448 155830 157457
rect 155774 157383 155830 157392
rect 155498 156904 155554 156913
rect 155498 156839 155554 156848
rect 155406 153776 155462 153785
rect 155406 153711 155462 153720
rect 155512 151162 155540 156839
rect 155788 153882 155816 157383
rect 155880 153921 155908 158743
rect 155866 153912 155922 153921
rect 155776 153876 155828 153882
rect 155866 153847 155922 153856
rect 155776 153818 155828 153824
rect 155500 151156 155552 151162
rect 155500 151098 155552 151104
rect 155314 149968 155370 149977
rect 155314 149903 155370 149912
rect 156524 149705 156552 159598
rect 156708 158574 156736 214610
rect 156696 158568 156748 158574
rect 156696 158510 156748 158516
rect 156604 158432 156656 158438
rect 156604 158374 156656 158380
rect 156510 149696 156566 149705
rect 156510 149631 156566 149640
rect 155960 145580 156012 145586
rect 155960 145522 156012 145528
rect 155224 45552 155276 45558
rect 155224 45494 155276 45500
rect 155972 16574 156000 145522
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 153844 4140 153896 4146
rect 153844 4082 153896 4088
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 156616 4826 156644 158374
rect 156708 158166 156736 158510
rect 156696 158160 156748 158166
rect 156696 158102 156748 158108
rect 156694 157040 156750 157049
rect 156694 156975 156750 156984
rect 156708 152425 156736 156975
rect 156800 156777 156828 225558
rect 156892 166274 156920 232698
rect 156984 166394 157012 233922
rect 157064 232552 157116 232558
rect 157064 232494 157116 232500
rect 156972 166388 157024 166394
rect 156972 166330 157024 166336
rect 156892 166246 157012 166274
rect 156880 166184 156932 166190
rect 156880 166126 156932 166132
rect 156892 159361 156920 166126
rect 156984 160410 157012 166246
rect 156972 160404 157024 160410
rect 156972 160346 157024 160352
rect 156984 159662 157012 160346
rect 156972 159656 157024 159662
rect 156972 159598 157024 159604
rect 156878 159352 156934 159361
rect 156878 159287 156934 159296
rect 156786 156768 156842 156777
rect 156786 156703 156842 156712
rect 156694 152416 156750 152425
rect 156694 152351 156750 152360
rect 156892 148481 156920 159287
rect 157076 154290 157104 232494
rect 157168 157049 157196 239527
rect 157260 157321 157288 241538
rect 158536 239488 158588 239494
rect 158536 239430 158588 239436
rect 158444 235272 158496 235278
rect 158444 235214 158496 235220
rect 158350 228304 158406 228313
rect 158350 228239 158406 228248
rect 158260 221536 158312 221542
rect 158260 221478 158312 221484
rect 158168 218748 158220 218754
rect 158168 218690 158220 218696
rect 158076 218068 158128 218074
rect 158076 218010 158128 218016
rect 157984 214736 158036 214742
rect 157984 214678 158036 214684
rect 157996 158098 158024 214678
rect 158088 160002 158116 218010
rect 158076 159996 158128 160002
rect 158076 159938 158128 159944
rect 157984 158092 158036 158098
rect 157984 158034 158036 158040
rect 157338 157720 157394 157729
rect 157338 157655 157394 157664
rect 157246 157312 157302 157321
rect 157246 157247 157302 157256
rect 157154 157040 157210 157049
rect 157154 156975 157210 156984
rect 157064 154284 157116 154290
rect 157064 154226 157116 154232
rect 157352 154057 157380 157655
rect 157338 154048 157394 154057
rect 157338 153983 157394 153992
rect 157340 153876 157392 153882
rect 157340 153818 157392 153824
rect 156878 148472 156934 148481
rect 156878 148407 156934 148416
rect 157352 16574 157380 153818
rect 158088 148617 158116 159938
rect 158180 157729 158208 218690
rect 158272 157865 158300 221478
rect 158364 159662 158392 228239
rect 158352 159656 158404 159662
rect 158352 159598 158404 159604
rect 158352 158704 158404 158710
rect 158352 158646 158404 158652
rect 158258 157856 158314 157865
rect 158258 157791 158314 157800
rect 158166 157720 158222 157729
rect 158166 157655 158222 157664
rect 158272 153105 158300 157791
rect 158258 153096 158314 153105
rect 158258 153031 158314 153040
rect 158074 148608 158130 148617
rect 158074 148543 158130 148552
rect 158364 98666 158392 158646
rect 158456 158001 158484 235214
rect 158548 159610 158576 239430
rect 158640 160682 158668 241703
rect 160008 241664 160060 241670
rect 160008 241606 160060 241612
rect 159914 241496 159970 241505
rect 159914 241431 159970 241440
rect 159732 239556 159784 239562
rect 159732 239498 159784 239504
rect 159640 235476 159692 235482
rect 159640 235418 159692 235424
rect 159454 235240 159510 235249
rect 159454 235175 159510 235184
rect 159272 212560 159324 212566
rect 159272 212502 159324 212508
rect 158628 160676 158680 160682
rect 158628 160618 158680 160624
rect 159180 160336 159232 160342
rect 159180 160278 159232 160284
rect 159192 159866 159220 160278
rect 159180 159860 159232 159866
rect 159180 159802 159232 159808
rect 158548 159582 158668 159610
rect 158640 159526 158668 159582
rect 158628 159520 158680 159526
rect 158628 159462 158680 159468
rect 158640 158846 158668 159462
rect 159284 159458 159312 212502
rect 159364 209908 159416 209914
rect 159364 209850 159416 209856
rect 159272 159452 159324 159458
rect 159272 159394 159324 159400
rect 158628 158840 158680 158846
rect 158628 158782 158680 158788
rect 158718 158672 158774 158681
rect 158718 158607 158774 158616
rect 158628 158092 158680 158098
rect 158628 158034 158680 158040
rect 158442 157992 158498 158001
rect 158442 157927 158498 157936
rect 158456 151298 158484 157927
rect 158640 157486 158668 158034
rect 158628 157480 158680 157486
rect 158628 157422 158680 157428
rect 158444 151292 158496 151298
rect 158444 151234 158496 151240
rect 158352 98660 158404 98666
rect 158352 98602 158404 98608
rect 158732 16574 158760 158607
rect 159376 137970 159404 209850
rect 159468 159225 159496 235175
rect 159548 232824 159600 232830
rect 159548 232766 159600 232772
rect 159454 159216 159510 159225
rect 159454 159151 159510 159160
rect 159468 150521 159496 159151
rect 159560 156466 159588 232766
rect 159652 157214 159680 235418
rect 159744 160449 159772 239498
rect 159824 236700 159876 236706
rect 159824 236642 159876 236648
rect 159730 160440 159786 160449
rect 159730 160375 159786 160384
rect 159640 157208 159692 157214
rect 159640 157150 159692 157156
rect 159548 156460 159600 156466
rect 159548 156402 159600 156408
rect 159836 155650 159864 236642
rect 159928 158681 159956 241431
rect 160020 160546 160048 241606
rect 161296 238128 161348 238134
rect 161296 238070 161348 238076
rect 161204 238060 161256 238066
rect 161204 238002 161256 238008
rect 161020 235408 161072 235414
rect 161020 235350 161072 235356
rect 160928 229764 160980 229770
rect 160928 229706 160980 229712
rect 160836 228404 160888 228410
rect 160836 228346 160888 228352
rect 160744 224256 160796 224262
rect 160744 224198 160796 224204
rect 160652 221468 160704 221474
rect 160652 221410 160704 221416
rect 160560 209976 160612 209982
rect 160560 209918 160612 209924
rect 160572 189038 160600 209918
rect 160560 189032 160612 189038
rect 160560 188974 160612 188980
rect 160008 160540 160060 160546
rect 160008 160482 160060 160488
rect 159914 158672 159970 158681
rect 159914 158607 159970 158616
rect 160098 158672 160154 158681
rect 160098 158607 160154 158616
rect 159928 158137 159956 158607
rect 159914 158128 159970 158137
rect 159914 158063 159970 158072
rect 159824 155644 159876 155650
rect 159824 155586 159876 155592
rect 159454 150512 159510 150521
rect 159454 150447 159510 150456
rect 159364 137964 159416 137970
rect 159364 137906 159416 137912
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 156604 4820 156656 4826
rect 156604 4762 156656 4768
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11830 160140 158607
rect 160664 158166 160692 221410
rect 160652 158160 160704 158166
rect 160652 158102 160704 158108
rect 160756 157962 160784 224198
rect 160848 158234 160876 228346
rect 160836 158228 160888 158234
rect 160836 158170 160888 158176
rect 160744 157956 160796 157962
rect 160744 157898 160796 157904
rect 160744 157752 160796 157758
rect 160744 157694 160796 157700
rect 160756 157593 160784 157694
rect 160940 157690 160968 229706
rect 161032 158506 161060 235350
rect 161112 234048 161164 234054
rect 161112 233990 161164 233996
rect 161124 158681 161152 233990
rect 161216 159730 161244 238002
rect 161204 159724 161256 159730
rect 161204 159666 161256 159672
rect 161308 159526 161336 238070
rect 162308 237448 162360 237454
rect 162308 237390 162360 237396
rect 161388 236836 161440 236842
rect 161388 236778 161440 236784
rect 161296 159520 161348 159526
rect 161296 159462 161348 159468
rect 161110 158672 161166 158681
rect 161110 158607 161166 158616
rect 161020 158500 161072 158506
rect 161020 158442 161072 158448
rect 161124 158273 161152 158607
rect 161110 158264 161166 158273
rect 161110 158199 161166 158208
rect 161400 158098 161428 236778
rect 161480 232688 161532 232694
rect 161480 232630 161532 232636
rect 161388 158092 161440 158098
rect 161388 158034 161440 158040
rect 161492 158030 161520 232630
rect 162216 229832 162268 229838
rect 162216 229774 162268 229780
rect 161572 228948 161624 228954
rect 161572 228890 161624 228896
rect 161584 161566 161612 228890
rect 161664 215960 161716 215966
rect 161664 215902 161716 215908
rect 161572 161560 161624 161566
rect 161572 161502 161624 161508
rect 161480 158024 161532 158030
rect 161480 157966 161532 157972
rect 160928 157684 160980 157690
rect 160928 157626 160980 157632
rect 160742 157584 160798 157593
rect 160742 157519 160798 157528
rect 161020 157412 161072 157418
rect 161020 157354 161072 157360
rect 160744 157140 160796 157146
rect 160744 157082 160796 157088
rect 160192 154284 160244 154290
rect 160192 154226 160244 154232
rect 160100 11824 160152 11830
rect 160100 11766 160152 11772
rect 160204 6914 160232 154226
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 160756 3602 160784 157082
rect 161032 119406 161060 157354
rect 161480 157004 161532 157010
rect 161480 156946 161532 156952
rect 161492 156602 161520 156946
rect 161480 156596 161532 156602
rect 161480 156538 161532 156544
rect 161584 123486 161612 161502
rect 161676 159866 161704 215902
rect 161756 214464 161808 214470
rect 161756 214406 161808 214412
rect 161768 159934 161796 214406
rect 162032 212356 162084 212362
rect 162032 212298 162084 212304
rect 161940 211948 161992 211954
rect 161940 211890 161992 211896
rect 161848 160676 161900 160682
rect 161848 160618 161900 160624
rect 161756 159928 161808 159934
rect 161756 159870 161808 159876
rect 161664 159860 161716 159866
rect 161664 159802 161716 159808
rect 161676 134570 161704 159802
rect 161768 147014 161796 159870
rect 161860 159118 161888 160618
rect 161848 159112 161900 159118
rect 161848 159054 161900 159060
rect 161848 157208 161900 157214
rect 161848 157150 161900 157156
rect 161860 156942 161888 157150
rect 161848 156936 161900 156942
rect 161848 156878 161900 156884
rect 161756 147008 161808 147014
rect 161756 146950 161808 146956
rect 161664 134564 161716 134570
rect 161664 134506 161716 134512
rect 161572 123480 161624 123486
rect 161572 123422 161624 123428
rect 161020 119400 161072 119406
rect 161020 119342 161072 119348
rect 161952 97306 161980 211890
rect 162044 211206 162072 212298
rect 162032 211200 162084 211206
rect 162032 211142 162084 211148
rect 161940 97300 161992 97306
rect 161940 97242 161992 97248
rect 162044 73846 162072 211142
rect 162228 166994 162256 229774
rect 162136 166966 162256 166994
rect 162136 158302 162164 166966
rect 162320 163010 162348 237390
rect 162688 211954 162716 293218
rect 164330 292768 164386 292777
rect 164330 292703 164386 292712
rect 162766 292632 162822 292641
rect 162766 292567 162822 292576
rect 162780 212362 162808 292567
rect 163504 239760 163556 239766
rect 163504 239702 163556 239708
rect 163516 212566 163544 239702
rect 164148 231260 164200 231266
rect 164148 231202 164200 231208
rect 163504 212560 163556 212566
rect 163504 212502 163556 212508
rect 162768 212356 162820 212362
rect 162768 212298 162820 212304
rect 162676 211948 162728 211954
rect 162676 211890 162728 211896
rect 163516 209930 163544 212502
rect 163516 209902 163990 209930
rect 164160 209545 164188 231202
rect 164344 229094 164372 292703
rect 164528 229094 164556 294578
rect 165896 294568 165948 294574
rect 165896 294510 165948 294516
rect 165710 282160 165766 282169
rect 165710 282095 165766 282104
rect 164344 229066 164464 229094
rect 164528 229066 164832 229094
rect 164330 212120 164386 212129
rect 164330 212055 164386 212064
rect 164344 209916 164372 212055
rect 164436 209930 164464 229066
rect 164804 209930 164832 229066
rect 165620 212492 165672 212498
rect 165620 212434 165672 212440
rect 165436 211200 165488 211206
rect 165436 211142 165488 211148
rect 164436 209902 164726 209930
rect 164804 209902 165094 209930
rect 165448 209916 165476 211142
rect 165632 209930 165660 212434
rect 165724 210066 165752 282095
rect 165908 229094 165936 294510
rect 166908 291848 166960 291854
rect 166908 291790 166960 291796
rect 165908 229066 166672 229094
rect 166540 211948 166592 211954
rect 166540 211890 166592 211896
rect 165724 210038 165936 210066
rect 165908 209930 165936 210038
rect 165632 209902 165830 209930
rect 165908 209902 166198 209930
rect 166552 209916 166580 211890
rect 166644 209930 166672 229066
rect 166920 212129 166948 291790
rect 167012 214606 167040 294646
rect 168380 294228 168432 294234
rect 168380 294170 168432 294176
rect 168288 290352 168340 290358
rect 168288 290294 168340 290300
rect 167092 244928 167144 244934
rect 167092 244870 167144 244876
rect 167000 214600 167052 214606
rect 167000 214542 167052 214548
rect 166906 212120 166962 212129
rect 166906 212055 166962 212064
rect 167104 209930 167132 244870
rect 167736 214600 167788 214606
rect 167736 214542 167788 214548
rect 167644 211948 167696 211954
rect 167644 211890 167696 211896
rect 166644 209902 166934 209930
rect 167104 209902 167302 209930
rect 167656 209916 167684 211890
rect 167748 209930 167776 214542
rect 168300 211954 168328 290294
rect 168392 214606 168420 294170
rect 168472 247716 168524 247722
rect 168472 247658 168524 247664
rect 168380 214600 168432 214606
rect 168380 214542 168432 214548
rect 168484 214538 168512 247658
rect 168564 246356 168616 246362
rect 168564 246298 168616 246304
rect 168472 214532 168524 214538
rect 168472 214474 168524 214480
rect 168288 211948 168340 211954
rect 168288 211890 168340 211896
rect 168300 211342 168328 211890
rect 168288 211336 168340 211342
rect 168288 211278 168340 211284
rect 168576 209930 168604 246298
rect 168840 214600 168892 214606
rect 168840 214542 168892 214548
rect 168748 211404 168800 211410
rect 168748 211346 168800 211352
rect 167748 209902 168038 209930
rect 168406 209902 168604 209930
rect 168760 209916 168788 211346
rect 168852 209930 168880 214542
rect 169208 214532 169260 214538
rect 169208 214474 169260 214480
rect 169220 209930 169248 214474
rect 169772 209953 169800 295870
rect 172520 295520 172572 295526
rect 172520 295462 172572 295468
rect 170404 294500 170456 294506
rect 170404 294442 170456 294448
rect 169852 294432 169904 294438
rect 169852 294374 169904 294380
rect 169864 214554 169892 294374
rect 169944 290012 169996 290018
rect 169944 289954 169996 289960
rect 169956 229094 169984 289954
rect 169956 229066 170352 229094
rect 169864 214526 170260 214554
rect 170128 211472 170180 211478
rect 170128 211414 170180 211420
rect 169758 209944 169814 209953
rect 168852 209902 169142 209930
rect 169220 209902 169510 209930
rect 169758 209879 169814 209888
rect 170140 209794 170168 211414
rect 170232 209916 170260 214526
rect 170324 210066 170352 229066
rect 170416 212498 170444 294442
rect 171140 294296 171192 294302
rect 171140 294238 171192 294244
rect 171152 214538 171180 294238
rect 171232 292800 171284 292806
rect 171232 292742 171284 292748
rect 171140 214532 171192 214538
rect 171140 214474 171192 214480
rect 170404 212492 170456 212498
rect 170404 212434 170456 212440
rect 170324 210038 170720 210066
rect 170402 209944 170458 209953
rect 170692 209930 170720 210038
rect 171244 209930 171272 292742
rect 171324 249076 171376 249082
rect 171324 249018 171376 249024
rect 171336 229094 171364 249018
rect 171336 229066 171456 229094
rect 171428 209930 171456 229066
rect 172532 214538 172560 295462
rect 172612 292868 172664 292874
rect 172612 292810 172664 292816
rect 172152 214532 172204 214538
rect 172152 214474 172204 214480
rect 172520 214532 172572 214538
rect 172520 214474 172572 214480
rect 172060 212016 172112 212022
rect 172060 211958 172112 211964
rect 170458 209902 170614 209930
rect 170692 209902 170982 209930
rect 171244 209902 171350 209930
rect 171428 209902 171718 209930
rect 172072 209916 172100 211958
rect 172164 209930 172192 214474
rect 172624 209930 172652 292810
rect 172704 290760 172756 290766
rect 172704 290702 172756 290708
rect 172716 229094 172744 290702
rect 172716 229066 172928 229094
rect 172900 209930 172928 229066
rect 173256 214532 173308 214538
rect 173256 214474 173308 214480
rect 173268 209930 173296 214474
rect 172164 209902 172454 209930
rect 172624 209902 172822 209930
rect 172900 209902 173190 209930
rect 173268 209902 173558 209930
rect 173912 209916 173940 297026
rect 175280 296948 175332 296954
rect 175280 296890 175332 296896
rect 173992 242208 174044 242214
rect 173992 242150 174044 242156
rect 174004 229094 174032 242150
rect 175292 229094 175320 296890
rect 178040 295588 178092 295594
rect 178040 295530 178092 295536
rect 176660 290148 176712 290154
rect 176660 290090 176712 290096
rect 174004 229066 174768 229094
rect 175292 229066 175872 229094
rect 174636 212084 174688 212090
rect 174636 212026 174688 212032
rect 174268 210724 174320 210730
rect 174268 210666 174320 210672
rect 174280 209916 174308 210666
rect 174648 209916 174676 212026
rect 174740 209930 174768 229066
rect 175740 212152 175792 212158
rect 175740 212094 175792 212100
rect 175372 211948 175424 211954
rect 175372 211890 175424 211896
rect 174740 209902 175030 209930
rect 175384 209916 175412 211890
rect 175752 209916 175780 212094
rect 175844 209930 175872 229066
rect 176476 212220 176528 212226
rect 176476 212162 176528 212168
rect 175844 209902 176134 209930
rect 176488 209916 176516 212162
rect 176672 209930 176700 290090
rect 176750 289096 176806 289105
rect 176750 289031 176806 289040
rect 176764 229094 176792 289031
rect 176764 229066 177712 229094
rect 177212 213444 177264 213450
rect 177212 213386 177264 213392
rect 176672 209902 176870 209930
rect 177224 209916 177252 213386
rect 177580 212492 177632 212498
rect 177580 212434 177632 212440
rect 177592 209916 177620 212434
rect 177684 209930 177712 229066
rect 178052 214538 178080 295530
rect 178132 293684 178184 293690
rect 178132 293626 178184 293632
rect 178040 214532 178092 214538
rect 178040 214474 178092 214480
rect 178144 209930 178172 293626
rect 178224 293616 178276 293622
rect 178224 293558 178276 293564
rect 178236 229094 178264 293558
rect 178684 292936 178736 292942
rect 178684 292878 178736 292884
rect 178236 229066 178448 229094
rect 178420 209930 178448 229066
rect 178696 212498 178724 292878
rect 178776 214532 178828 214538
rect 178776 214474 178828 214480
rect 178684 212492 178736 212498
rect 178684 212434 178736 212440
rect 178788 209930 178816 214474
rect 177684 209902 177974 209930
rect 178144 209902 178342 209930
rect 178420 209902 178710 209930
rect 178788 209902 179078 209930
rect 179432 209916 179460 297162
rect 186320 297016 186372 297022
rect 186320 296958 186372 296964
rect 183560 296812 183612 296818
rect 183560 296754 183612 296760
rect 182180 295656 182232 295662
rect 182180 295598 182232 295604
rect 180800 294364 180852 294370
rect 180800 294306 180852 294312
rect 179512 290488 179564 290494
rect 179512 290430 179564 290436
rect 179524 229094 179552 290430
rect 180064 289264 180116 289270
rect 180064 289206 180116 289212
rect 179524 229066 179920 229094
rect 179788 212288 179840 212294
rect 179788 212230 179840 212236
rect 179800 209916 179828 212230
rect 179892 209930 179920 229066
rect 180076 212158 180104 289206
rect 180812 214538 180840 294306
rect 180890 288552 180946 288561
rect 180890 288487 180946 288496
rect 180904 229094 180932 288487
rect 180904 229066 181024 229094
rect 180892 216028 180944 216034
rect 180892 215970 180944 215976
rect 180800 214532 180852 214538
rect 180800 214474 180852 214480
rect 180064 212152 180116 212158
rect 180064 212094 180116 212100
rect 180524 212016 180576 212022
rect 180524 211958 180576 211964
rect 179892 209902 180182 209930
rect 180536 209916 180564 211958
rect 180904 209916 180932 215970
rect 180996 209930 181024 229066
rect 181352 214532 181404 214538
rect 181352 214474 181404 214480
rect 181364 209930 181392 214474
rect 181996 213376 182048 213382
rect 181996 213318 182048 213324
rect 180996 209902 181286 209930
rect 181364 209902 181654 209930
rect 182008 209916 182036 213318
rect 182192 209930 182220 295598
rect 182272 289876 182324 289882
rect 182272 289818 182324 289824
rect 182284 214538 182312 289818
rect 182364 279472 182416 279478
rect 182364 279414 182416 279420
rect 182376 229094 182404 279414
rect 182916 238196 182968 238202
rect 182916 238138 182968 238144
rect 182928 235521 182956 238138
rect 182914 235512 182970 235521
rect 182914 235447 182970 235456
rect 182376 229066 182496 229094
rect 182272 214532 182324 214538
rect 182272 214474 182324 214480
rect 182468 209930 182496 229066
rect 183100 214804 183152 214810
rect 183100 214746 183152 214752
rect 182548 211404 182600 211410
rect 182548 211346 182600 211352
rect 182560 210089 182588 211346
rect 182546 210080 182602 210089
rect 182546 210015 182602 210024
rect 182192 209902 182390 209930
rect 182468 209902 182758 209930
rect 183112 209916 183140 214746
rect 183572 214538 183600 296754
rect 184940 289196 184992 289202
rect 184940 289138 184992 289144
rect 183652 288448 183704 288454
rect 183652 288390 183704 288396
rect 183192 214532 183244 214538
rect 183192 214474 183244 214480
rect 183560 214532 183612 214538
rect 183560 214474 183612 214480
rect 183204 209930 183232 214474
rect 183664 214470 183692 288390
rect 183744 286340 183796 286346
rect 183744 286282 183796 286288
rect 183756 229094 183784 286282
rect 183756 229066 183876 229094
rect 183652 214464 183704 214470
rect 183652 214406 183704 214412
rect 183468 211268 183520 211274
rect 183468 211210 183520 211216
rect 183480 210662 183508 211210
rect 183468 210656 183520 210662
rect 183468 210598 183520 210604
rect 183204 209902 183494 209930
rect 183848 209916 183876 229066
rect 184296 214532 184348 214538
rect 184296 214474 184348 214480
rect 183928 214464 183980 214470
rect 183928 214406 183980 214412
rect 183940 209930 183968 214406
rect 184308 209930 184336 214474
rect 184952 214470 184980 289138
rect 185032 289128 185084 289134
rect 185032 289070 185084 289076
rect 185044 214538 185072 289070
rect 185124 276684 185176 276690
rect 185124 276626 185176 276632
rect 185032 214532 185084 214538
rect 185032 214474 185084 214480
rect 184940 214464 184992 214470
rect 184940 214406 184992 214412
rect 184848 213240 184900 213246
rect 184848 213182 184900 213188
rect 183940 209902 184230 209930
rect 184308 209902 184598 209930
rect 170402 209879 170458 209888
rect 169878 209766 170168 209794
rect 184860 209545 184888 213182
rect 185136 209930 185164 276626
rect 186332 214538 186360 296958
rect 187700 296880 187752 296886
rect 187700 296822 187752 296828
rect 186964 295792 187016 295798
rect 186964 295734 187016 295740
rect 186410 288688 186466 288697
rect 186410 288623 186466 288632
rect 185400 214532 185452 214538
rect 185400 214474 185452 214480
rect 186320 214532 186372 214538
rect 186320 214474 186372 214480
rect 185216 214464 185268 214470
rect 185216 214406 185268 214412
rect 184966 209902 185164 209930
rect 185228 209930 185256 214406
rect 185412 209930 185440 214474
rect 186044 214260 186096 214266
rect 186044 214202 186096 214208
rect 185228 209902 185334 209930
rect 185412 209902 185702 209930
rect 186056 209916 186084 214202
rect 186320 212424 186372 212430
rect 186320 212366 186372 212372
rect 186332 210594 186360 212366
rect 186320 210588 186372 210594
rect 186320 210530 186372 210536
rect 186424 209916 186452 288623
rect 186504 239624 186556 239630
rect 186504 239566 186556 239572
rect 186516 229094 186544 239566
rect 186516 229066 186912 229094
rect 186504 214532 186556 214538
rect 186504 214474 186556 214480
rect 186516 209930 186544 214474
rect 186884 209930 186912 229066
rect 186976 212158 187004 295734
rect 187516 217388 187568 217394
rect 187516 217330 187568 217336
rect 186964 212152 187016 212158
rect 186964 212094 187016 212100
rect 186516 209902 186806 209930
rect 186884 209902 187174 209930
rect 187528 209916 187556 217330
rect 187712 214538 187740 296822
rect 189080 295384 189132 295390
rect 189080 295326 189132 295332
rect 187790 289232 187846 289241
rect 187790 289167 187846 289176
rect 187700 214532 187752 214538
rect 187700 214474 187752 214480
rect 187804 214470 187832 289167
rect 187884 273964 187936 273970
rect 187884 273906 187936 273912
rect 187896 229094 187924 273906
rect 187896 229066 188016 229094
rect 187792 214464 187844 214470
rect 187792 214406 187844 214412
rect 187884 212492 187936 212498
rect 187884 212434 187936 212440
rect 187608 211472 187660 211478
rect 187608 211414 187660 211420
rect 187620 209774 187648 211414
rect 187896 209916 187924 212434
rect 187988 209930 188016 229066
rect 189092 214538 189120 295326
rect 193220 294840 193272 294846
rect 193220 294782 193272 294788
rect 189724 293004 189776 293010
rect 189724 292946 189776 292952
rect 189172 240780 189224 240786
rect 189172 240722 189224 240728
rect 188344 214532 188396 214538
rect 188344 214474 188396 214480
rect 189080 214532 189132 214538
rect 189080 214474 189132 214480
rect 188356 209930 188384 214474
rect 188712 214464 188764 214470
rect 188712 214406 188764 214412
rect 188724 209930 188752 214406
rect 189080 211744 189132 211750
rect 189080 211686 189132 211692
rect 189092 210526 189120 211686
rect 189080 210520 189132 210526
rect 189080 210462 189132 210468
rect 189184 209930 189212 240722
rect 189736 219434 189764 292946
rect 189908 292188 189960 292194
rect 189908 292130 189960 292136
rect 189814 289504 189870 289513
rect 189814 289439 189870 289448
rect 189644 219406 189764 219434
rect 189644 212294 189672 219406
rect 189828 214690 189856 289439
rect 189736 214662 189856 214690
rect 189736 212498 189764 214662
rect 189816 214532 189868 214538
rect 189816 214474 189868 214480
rect 189724 212492 189776 212498
rect 189724 212434 189776 212440
rect 189632 212288 189684 212294
rect 189632 212230 189684 212236
rect 189724 212152 189776 212158
rect 189724 212094 189776 212100
rect 189540 211336 189592 211342
rect 189540 211278 189592 211284
rect 187988 209902 188278 209930
rect 188356 209902 188646 209930
rect 188724 209902 189014 209930
rect 189184 209902 189382 209930
rect 187700 209774 187752 209778
rect 187620 209772 187752 209774
rect 187620 209746 187700 209772
rect 187700 209714 187752 209720
rect 189552 209545 189580 211278
rect 189736 209916 189764 212094
rect 189828 209930 189856 214474
rect 189920 214266 189948 292130
rect 190642 290728 190698 290737
rect 190642 290663 190698 290672
rect 190458 289912 190514 289921
rect 190458 289847 190514 289856
rect 190472 214538 190500 289847
rect 190550 272504 190606 272513
rect 190550 272439 190606 272448
rect 190460 214532 190512 214538
rect 190460 214474 190512 214480
rect 189908 214260 189960 214266
rect 189908 214202 189960 214208
rect 190564 209930 190592 272439
rect 189828 209902 190118 209930
rect 190486 209902 190592 209930
rect 190656 209930 190684 290663
rect 192206 290592 192262 290601
rect 192206 290527 192262 290536
rect 192022 290456 192078 290465
rect 192022 290391 192078 290400
rect 191838 290048 191894 290057
rect 191838 289983 191894 289992
rect 190734 242176 190790 242185
rect 190734 242111 190790 242120
rect 190748 229094 190776 242111
rect 191656 238332 191708 238338
rect 191656 238274 191708 238280
rect 191668 232694 191696 238274
rect 191656 232688 191708 232694
rect 191656 232630 191708 232636
rect 190748 229066 191328 229094
rect 190920 214532 190972 214538
rect 190920 214474 190972 214480
rect 190932 209930 190960 214474
rect 191300 209930 191328 229066
rect 191748 211336 191800 211342
rect 191748 211278 191800 211284
rect 191760 210458 191788 211278
rect 191748 210452 191800 210458
rect 191748 210394 191800 210400
rect 191852 209930 191880 289983
rect 191932 243568 191984 243574
rect 191932 243510 191984 243516
rect 191944 214538 191972 243510
rect 191932 214532 191984 214538
rect 191932 214474 191984 214480
rect 192036 209930 192064 290391
rect 192220 229094 192248 290527
rect 192484 238400 192536 238406
rect 192484 238342 192536 238348
rect 192496 232529 192524 238342
rect 192482 232520 192538 232529
rect 192482 232455 192538 232464
rect 192220 229066 192800 229094
rect 192392 214532 192444 214538
rect 192392 214474 192444 214480
rect 192404 209930 192432 214474
rect 192772 209930 192800 229066
rect 193232 210322 193260 294782
rect 193312 290556 193364 290562
rect 193312 290498 193364 290504
rect 193324 214538 193352 290498
rect 193404 284980 193456 284986
rect 193404 284922 193456 284928
rect 193416 229094 193444 284922
rect 194324 238264 194376 238270
rect 194324 238206 194376 238212
rect 194336 232393 194364 238206
rect 194416 232892 194468 232898
rect 194416 232834 194468 232840
rect 194322 232384 194378 232393
rect 194322 232319 194378 232328
rect 193416 229066 193536 229094
rect 193404 216096 193456 216102
rect 193404 216038 193456 216044
rect 193312 214532 193364 214538
rect 193312 214474 193364 214480
rect 193220 210316 193272 210322
rect 193220 210258 193272 210264
rect 190656 209902 190854 209930
rect 190932 209902 191222 209930
rect 191300 209902 191590 209930
rect 191852 209902 191958 209930
rect 192036 209902 192326 209930
rect 192404 209902 192694 209930
rect 192772 209902 193062 209930
rect 193416 209916 193444 216038
rect 193508 209930 193536 229066
rect 193864 214532 193916 214538
rect 193864 214474 193916 214480
rect 193876 209930 193904 214474
rect 193508 209902 193798 209930
rect 193876 209902 194166 209930
rect 194428 209545 194456 232834
rect 194612 214538 194640 298114
rect 194692 290624 194744 290630
rect 194692 290566 194744 290572
rect 194600 214532 194652 214538
rect 194600 214474 194652 214480
rect 194704 212770 194732 290566
rect 194784 286408 194836 286414
rect 194784 286350 194836 286356
rect 194796 229094 194824 286350
rect 195888 232688 195940 232694
rect 195888 232630 195940 232636
rect 194796 229066 194916 229094
rect 194692 212764 194744 212770
rect 194692 212706 194744 212712
rect 194508 210316 194560 210322
rect 194508 210258 194560 210264
rect 194520 209916 194548 210258
rect 194888 209916 194916 229066
rect 195336 214532 195388 214538
rect 195336 214474 195388 214480
rect 194968 212764 195020 212770
rect 194968 212706 195020 212712
rect 194980 209930 195008 212706
rect 195348 209930 195376 214474
rect 194980 209902 195270 209930
rect 195348 209902 195638 209930
rect 195900 209545 195928 232630
rect 195992 211070 196020 299610
rect 196072 283620 196124 283626
rect 196072 283562 196124 283568
rect 195980 211064 196032 211070
rect 195980 211006 196032 211012
rect 196084 209930 196112 283562
rect 196164 280832 196216 280838
rect 196164 280774 196216 280780
rect 196176 229094 196204 280774
rect 196176 229066 196848 229094
rect 196348 212424 196400 212430
rect 196348 212366 196400 212372
rect 196006 209902 196112 209930
rect 196360 209916 196388 212366
rect 196440 211064 196492 211070
rect 196440 211006 196492 211012
rect 196452 209930 196480 211006
rect 196820 209930 196848 229066
rect 197372 210594 197400 300902
rect 199660 293548 199712 293554
rect 199660 293490 199712 293496
rect 199672 292602 199700 293490
rect 198740 292596 198792 292602
rect 198740 292538 198792 292544
rect 199660 292596 199712 292602
rect 199660 292538 199712 292544
rect 197544 290692 197596 290698
rect 197544 290634 197596 290640
rect 197452 289944 197504 289950
rect 197452 289886 197504 289892
rect 197464 212294 197492 289886
rect 197452 212288 197504 212294
rect 197452 212230 197504 212236
rect 197556 212106 197584 290634
rect 198648 231124 198700 231130
rect 198648 231066 198700 231072
rect 198464 230512 198516 230518
rect 198464 230454 198516 230460
rect 197912 228472 197964 228478
rect 197912 228414 197964 228420
rect 197464 212078 197584 212106
rect 197360 210588 197412 210594
rect 197360 210530 197412 210536
rect 196452 209902 196742 209930
rect 196820 209902 197110 209930
rect 197464 209916 197492 212078
rect 197636 210588 197688 210594
rect 197636 210530 197688 210536
rect 197648 209930 197676 210530
rect 197924 209930 197952 228414
rect 197648 209902 197846 209930
rect 197924 209902 198214 209930
rect 198476 209545 198504 230454
rect 198556 212288 198608 212294
rect 198556 212230 198608 212236
rect 198568 209916 198596 212230
rect 198660 210089 198688 231066
rect 198646 210080 198702 210089
rect 198646 210015 198702 210024
rect 198752 209930 198780 292538
rect 199384 290080 199436 290086
rect 199384 290022 199436 290028
rect 199396 241466 199424 290022
rect 198832 241460 198884 241466
rect 198832 241402 198884 241408
rect 199384 241460 199436 241466
rect 199384 241402 199436 241408
rect 198844 212106 198872 241402
rect 198924 239692 198976 239698
rect 198924 239634 198976 239640
rect 198936 239426 198964 239634
rect 198924 239420 198976 239426
rect 198924 239362 198976 239368
rect 198936 212294 198964 239362
rect 199844 231328 199896 231334
rect 199844 231270 199896 231276
rect 199752 230580 199804 230586
rect 199752 230522 199804 230528
rect 199212 212350 199424 212378
rect 198924 212288 198976 212294
rect 198924 212230 198976 212236
rect 199212 212106 199240 212350
rect 199292 212220 199344 212226
rect 199292 212162 199344 212168
rect 198844 212078 199240 212106
rect 198752 209902 198950 209930
rect 199304 209916 199332 212162
rect 199396 209930 199424 212350
rect 199396 209902 199686 209930
rect 199200 209636 199252 209642
rect 199200 209578 199252 209584
rect 199212 209545 199240 209578
rect 164146 209536 164202 209545
rect 164146 209471 164202 209480
rect 184846 209536 184902 209545
rect 184846 209471 184902 209480
rect 189538 209536 189594 209545
rect 189538 209471 189594 209480
rect 194414 209536 194470 209545
rect 194414 209471 194470 209480
rect 195886 209536 195942 209545
rect 195886 209471 195942 209480
rect 198462 209536 198518 209545
rect 198462 209471 198518 209480
rect 199198 209536 199254 209545
rect 199764 209522 199792 230522
rect 199856 209642 199884 231270
rect 199936 231192 199988 231198
rect 199936 231134 199988 231140
rect 199948 209817 199976 231134
rect 200028 212288 200080 212294
rect 200028 212230 200080 212236
rect 200040 209916 200068 212230
rect 200132 210798 200160 302194
rect 200764 293072 200816 293078
rect 200764 293014 200816 293020
rect 200212 253904 200264 253910
rect 200212 253846 200264 253852
rect 200120 210792 200172 210798
rect 200120 210734 200172 210740
rect 200224 209930 200252 253846
rect 200672 213920 200724 213926
rect 200672 213862 200724 213868
rect 200684 212498 200712 213862
rect 200580 212492 200632 212498
rect 200580 212434 200632 212440
rect 200672 212492 200724 212498
rect 200672 212434 200724 212440
rect 200592 212294 200620 212434
rect 200580 212288 200632 212294
rect 200580 212230 200632 212236
rect 200684 209930 200712 212434
rect 200776 212362 200804 293014
rect 201224 228608 201276 228614
rect 201224 228550 201276 228556
rect 200764 212356 200816 212362
rect 200764 212298 200816 212304
rect 201236 212294 201264 228550
rect 201224 212288 201276 212294
rect 201224 212230 201276 212236
rect 201236 211818 201264 212230
rect 201420 212106 201448 303622
rect 201684 299600 201736 299606
rect 201684 299542 201736 299548
rect 201420 212078 201540 212106
rect 201512 211886 201540 212078
rect 201500 211880 201552 211886
rect 201500 211822 201552 211828
rect 201224 211812 201276 211818
rect 201224 211754 201276 211760
rect 201132 210792 201184 210798
rect 201132 210734 201184 210740
rect 200948 209976 201000 209982
rect 200224 209902 200422 209930
rect 200684 209902 200790 209930
rect 201144 209930 201172 210734
rect 201000 209924 201172 209930
rect 200948 209918 201172 209924
rect 200960 209916 201172 209918
rect 201512 209916 201540 211822
rect 200960 209902 201158 209916
rect 201696 209914 201724 299542
rect 202144 295724 202196 295730
rect 202144 295666 202196 295672
rect 202156 211342 202184 295666
rect 202604 228132 202656 228138
rect 202604 228074 202656 228080
rect 202616 215294 202644 228074
rect 202708 226302 202736 312734
rect 202788 300892 202840 300898
rect 202788 300834 202840 300840
rect 202696 226296 202748 226302
rect 202696 226238 202748 226244
rect 202708 225622 202736 226238
rect 202696 225616 202748 225622
rect 202696 225558 202748 225564
rect 202616 215266 202736 215294
rect 202708 212362 202736 215266
rect 202696 212356 202748 212362
rect 202696 212298 202748 212304
rect 202800 212294 202828 300834
rect 202880 298240 202932 298246
rect 202880 298182 202932 298188
rect 202892 214062 202920 298182
rect 202972 290216 203024 290222
rect 202972 290158 203024 290164
rect 202984 215234 203012 290158
rect 204088 218006 204116 321574
rect 204076 218000 204128 218006
rect 204076 217942 204128 217948
rect 204088 217326 204116 217942
rect 204076 217320 204128 217326
rect 204076 217262 204128 217268
rect 202984 215206 203104 215234
rect 202880 214056 202932 214062
rect 202880 213998 202932 214004
rect 202880 213920 202932 213926
rect 202880 213862 202932 213868
rect 202892 213314 202920 213862
rect 202880 213308 202932 213314
rect 202880 213250 202932 213256
rect 202604 212288 202656 212294
rect 202604 212230 202656 212236
rect 202788 212288 202840 212294
rect 202788 212230 202840 212236
rect 202144 211336 202196 211342
rect 202144 211278 202196 211284
rect 202156 209930 202184 211278
rect 202420 209976 202472 209982
rect 201684 209908 201736 209914
rect 201894 209902 202184 209930
rect 202262 209924 202420 209930
rect 202262 209918 202472 209924
rect 202262 209902 202460 209918
rect 202616 209916 202644 212230
rect 202800 211750 202828 212230
rect 202788 211744 202840 211750
rect 202788 211686 202840 211692
rect 201684 209850 201736 209856
rect 199934 209808 199990 209817
rect 199934 209743 199990 209752
rect 199844 209636 199896 209642
rect 199844 209578 199896 209584
rect 199842 209536 199898 209545
rect 199764 209494 199842 209522
rect 199198 209471 199254 209480
rect 199842 209471 199898 209480
rect 202880 209432 202932 209438
rect 203076 209386 203104 215206
rect 203156 214056 203208 214062
rect 203156 213998 203208 214004
rect 203168 209438 203196 213998
rect 204180 213926 204208 322079
rect 205546 321600 205602 321609
rect 205546 321535 205602 321544
rect 205454 316704 205510 316713
rect 205454 316639 205510 316648
rect 204902 307184 204958 307193
rect 204902 307119 204958 307128
rect 204536 303748 204588 303754
rect 204536 303690 204588 303696
rect 204352 302320 204404 302326
rect 204352 302262 204404 302268
rect 204364 219434 204392 302262
rect 204444 297152 204496 297158
rect 204444 297094 204496 297100
rect 204272 219406 204392 219434
rect 204168 213920 204220 213926
rect 204168 213862 204220 213868
rect 203708 212356 203760 212362
rect 203708 212298 203760 212304
rect 203340 212288 203392 212294
rect 203340 212230 203392 212236
rect 203352 209916 203380 212230
rect 203720 209916 203748 212298
rect 204272 209930 204300 219406
rect 204456 215294 204484 297094
rect 204180 209902 204300 209930
rect 204364 215266 204484 215294
rect 204180 209658 204208 209902
rect 204180 209630 204300 209658
rect 204272 209545 204300 209630
rect 204258 209536 204314 209545
rect 204258 209471 204314 209480
rect 204364 209438 204392 215266
rect 204548 209794 204576 303690
rect 204916 241670 204944 307119
rect 204904 241664 204956 241670
rect 204904 241606 204956 241612
rect 205468 239562 205496 316639
rect 205088 239556 205140 239562
rect 205088 239498 205140 239504
rect 205456 239556 205508 239562
rect 205456 239498 205508 239504
rect 205100 239057 205128 239498
rect 205086 239048 205142 239057
rect 205086 238983 205142 238992
rect 205560 237250 205588 321535
rect 208308 320952 208360 320958
rect 208308 320894 208360 320900
rect 208216 318912 208268 318918
rect 206926 318880 206982 318889
rect 208216 318854 208268 318860
rect 206926 318815 206982 318824
rect 206742 318200 206798 318209
rect 206742 318135 206798 318144
rect 206374 308544 206430 308553
rect 206374 308479 206430 308488
rect 206284 305040 206336 305046
rect 206284 304982 206336 304988
rect 205548 237244 205600 237250
rect 205548 237186 205600 237192
rect 205560 233209 205588 237186
rect 205546 233200 205602 233209
rect 205546 233135 205602 233144
rect 205732 215280 205784 215286
rect 205732 215222 205784 215228
rect 205640 215212 205692 215218
rect 205640 215154 205692 215160
rect 205652 214742 205680 215154
rect 205640 214736 205692 214742
rect 205640 214678 205692 214684
rect 205744 214674 205772 215222
rect 205732 214668 205784 214674
rect 205732 214610 205784 214616
rect 204812 211540 204864 211546
rect 204812 211482 204864 211488
rect 204824 209916 204852 211482
rect 206296 211274 206324 304982
rect 206388 241602 206416 308479
rect 206652 296744 206704 296750
rect 206652 296686 206704 296692
rect 206376 241596 206428 241602
rect 206376 241538 206428 241544
rect 206388 240310 206416 241538
rect 206664 240718 206692 296686
rect 206652 240712 206704 240718
rect 206652 240654 206704 240660
rect 206376 240304 206428 240310
rect 206376 240246 206428 240252
rect 206664 236745 206692 240654
rect 206650 236736 206706 236745
rect 206650 236671 206706 236680
rect 206756 219337 206784 318135
rect 206836 318096 206888 318102
rect 206836 318038 206888 318044
rect 206742 219328 206798 219337
rect 206742 219263 206798 219272
rect 206756 218929 206784 219263
rect 206742 218920 206798 218929
rect 206742 218855 206798 218864
rect 206848 215286 206876 318038
rect 206836 215280 206888 215286
rect 206836 215222 206888 215228
rect 206940 215218 206968 318815
rect 207940 308644 207992 308650
rect 207940 308586 207992 308592
rect 207848 298308 207900 298314
rect 207848 298250 207900 298256
rect 207664 241596 207716 241602
rect 207664 241538 207716 241544
rect 207020 235884 207072 235890
rect 207020 235826 207072 235832
rect 207032 235482 207060 235826
rect 207020 235476 207072 235482
rect 207020 235418 207072 235424
rect 207020 235204 207072 235210
rect 207020 235146 207072 235152
rect 207032 232762 207060 235146
rect 207020 232756 207072 232762
rect 207020 232698 207072 232704
rect 206928 215212 206980 215218
rect 206928 215154 206980 215160
rect 206284 211268 206336 211274
rect 206284 211210 206336 211216
rect 206296 209930 206324 211210
rect 205942 209902 206324 209930
rect 204628 209840 204680 209846
rect 204470 209788 204628 209794
rect 204470 209782 204680 209788
rect 204470 209766 204668 209782
rect 202932 209380 203104 209386
rect 202880 209374 203104 209380
rect 203156 209432 203208 209438
rect 203156 209374 203208 209380
rect 203892 209432 203944 209438
rect 204352 209432 204404 209438
rect 203944 209380 204102 209386
rect 203892 209374 204102 209380
rect 204352 209374 204404 209380
rect 204996 209432 205048 209438
rect 205048 209380 205206 209386
rect 204996 209374 205206 209380
rect 202892 209358 203104 209374
rect 203904 209358 204102 209374
rect 205008 209358 205206 209374
rect 205537 209208 205546 209264
rect 205602 209208 205611 209264
rect 207478 174584 207534 174593
rect 207478 174519 207534 174528
rect 207492 164234 207520 174519
rect 207492 164206 207612 164234
rect 162228 162982 162348 163010
rect 162228 159050 162256 162982
rect 162400 161560 162452 161566
rect 162452 161508 162532 161514
rect 162400 161502 162532 161508
rect 162412 161486 162532 161502
rect 162504 160684 162532 161486
rect 207480 161288 207532 161294
rect 207480 161230 207532 161236
rect 207492 160954 207520 161230
rect 207480 160948 207532 160954
rect 207480 160890 207532 160896
rect 162308 160472 162360 160478
rect 162308 160414 162360 160420
rect 162320 159780 162348 160414
rect 162596 159934 162624 160140
rect 162584 159928 162636 159934
rect 162584 159870 162636 159876
rect 162688 159866 162716 160140
rect 162676 159860 162728 159866
rect 162676 159802 162728 159808
rect 162492 159792 162544 159798
rect 162320 159752 162492 159780
rect 162780 159746 162808 160140
rect 162872 159769 162900 160140
rect 162964 159905 162992 160140
rect 162950 159896 163006 159905
rect 162950 159831 163006 159840
rect 162492 159734 162544 159740
rect 162216 159044 162268 159050
rect 162216 158986 162268 158992
rect 162124 158296 162176 158302
rect 162124 158238 162176 158244
rect 162124 157276 162176 157282
rect 162124 157218 162176 157224
rect 162032 73840 162084 73846
rect 162032 73782 162084 73788
rect 161296 11824 161348 11830
rect 161296 11766 161348 11772
rect 160744 3596 160796 3602
rect 160744 3538 160796 3544
rect 161308 480 161336 11766
rect 162136 3534 162164 157218
rect 162504 157185 162532 159734
rect 162596 159718 162808 159746
rect 162858 159760 162914 159769
rect 162596 158030 162624 159718
rect 162858 159695 162914 159704
rect 162952 159724 163004 159730
rect 162676 159656 162728 159662
rect 162676 159598 162728 159604
rect 162688 159186 162716 159598
rect 162768 159384 162820 159390
rect 162768 159326 162820 159332
rect 162676 159180 162728 159186
rect 162676 159122 162728 159128
rect 162584 158024 162636 158030
rect 162584 157966 162636 157972
rect 162490 157176 162546 157185
rect 162490 157111 162546 157120
rect 162688 151814 162716 159122
rect 162780 157350 162808 159326
rect 162872 158914 162900 159695
rect 162952 159666 163004 159672
rect 162964 159118 162992 159666
rect 163056 159508 163084 160140
rect 163148 159939 163176 160140
rect 163134 159930 163190 159939
rect 163134 159865 163190 159874
rect 163056 159480 163176 159508
rect 163148 159118 163176 159480
rect 162952 159112 163004 159118
rect 162952 159054 163004 159060
rect 163136 159112 163188 159118
rect 163136 159054 163188 159060
rect 162860 158908 162912 158914
rect 162860 158850 162912 158856
rect 162860 158772 162912 158778
rect 162860 158714 162912 158720
rect 162768 157344 162820 157350
rect 162768 157286 162820 157292
rect 162688 151786 162808 151814
rect 162780 3602 162808 151786
rect 162872 140078 162900 158714
rect 162860 140072 162912 140078
rect 162860 140014 162912 140020
rect 162964 124914 162992 159054
rect 163240 158914 163268 160140
rect 163136 158908 163188 158914
rect 163136 158850 163188 158856
rect 163228 158908 163280 158914
rect 163228 158850 163280 158856
rect 163148 158692 163176 158850
rect 163332 158760 163360 160140
rect 163424 159866 163452 160140
rect 163412 159860 163464 159866
rect 163412 159802 163464 159808
rect 163516 159390 163544 160140
rect 163608 159905 163636 160140
rect 163594 159896 163650 159905
rect 163594 159831 163650 159840
rect 163504 159384 163556 159390
rect 163504 159326 163556 159332
rect 163412 158908 163464 158914
rect 163464 158868 163544 158896
rect 163412 158850 163464 158856
rect 163332 158732 163452 158760
rect 163148 158664 163268 158692
rect 163136 158568 163188 158574
rect 163136 158510 163188 158516
rect 163044 157752 163096 157758
rect 163044 157694 163096 157700
rect 163056 157457 163084 157694
rect 163042 157448 163098 157457
rect 163042 157383 163098 157392
rect 163044 157344 163096 157350
rect 163044 157286 163096 157292
rect 163056 129062 163084 157286
rect 163148 149734 163176 158510
rect 163136 149728 163188 149734
rect 163136 149670 163188 149676
rect 163044 129056 163096 129062
rect 163044 128998 163096 129004
rect 162952 124908 163004 124914
rect 162952 124850 163004 124856
rect 163240 95946 163268 158664
rect 163318 158672 163374 158681
rect 163318 158607 163374 158616
rect 163332 109750 163360 158607
rect 163424 157554 163452 158732
rect 163516 157593 163544 158868
rect 163608 158574 163636 159831
rect 163700 159798 163728 160140
rect 163688 159792 163740 159798
rect 163688 159734 163740 159740
rect 163688 159112 163740 159118
rect 163688 159054 163740 159060
rect 163596 158568 163648 158574
rect 163596 158510 163648 158516
rect 163700 158506 163728 159054
rect 163688 158500 163740 158506
rect 163688 158442 163740 158448
rect 163502 157584 163558 157593
rect 163412 157548 163464 157554
rect 163502 157519 163558 157528
rect 163412 157490 163464 157496
rect 163504 157344 163556 157350
rect 163504 157286 163556 157292
rect 163412 157208 163464 157214
rect 163412 157150 163464 157156
rect 163424 117978 163452 157150
rect 163516 157010 163544 157286
rect 163504 157004 163556 157010
rect 163504 156946 163556 156952
rect 163596 157004 163648 157010
rect 163596 156946 163648 156952
rect 163412 117972 163464 117978
rect 163412 117914 163464 117920
rect 163504 117972 163556 117978
rect 163504 117914 163556 117920
rect 163320 109744 163372 109750
rect 163320 109686 163372 109692
rect 163228 95940 163280 95946
rect 163228 95882 163280 95888
rect 162768 3596 162820 3602
rect 162768 3538 162820 3544
rect 163516 3534 163544 117914
rect 163608 116618 163636 156946
rect 163700 133210 163728 158442
rect 163792 157334 163820 160140
rect 163884 159769 163912 160140
rect 163870 159760 163926 159769
rect 163870 159695 163926 159704
rect 163884 158438 163912 159695
rect 163872 158432 163924 158438
rect 163872 158374 163924 158380
rect 163976 158250 164004 160140
rect 164068 159905 164096 160140
rect 164054 159896 164110 159905
rect 164054 159831 164110 159840
rect 164068 158778 164096 159831
rect 164160 159254 164188 160140
rect 164252 159769 164280 160140
rect 164238 159760 164294 159769
rect 164238 159695 164294 159704
rect 164240 159316 164292 159322
rect 164240 159258 164292 159264
rect 164148 159248 164200 159254
rect 164148 159190 164200 159196
rect 164056 158772 164108 158778
rect 164056 158714 164108 158720
rect 163976 158222 164096 158250
rect 164068 157418 164096 158222
rect 164056 157412 164108 157418
rect 164056 157354 164108 157360
rect 163792 157306 164004 157334
rect 163976 157214 164004 157306
rect 163964 157208 164016 157214
rect 163964 157150 164016 157156
rect 164160 157010 164188 159190
rect 164252 158681 164280 159258
rect 164238 158672 164294 158681
rect 164238 158607 164294 158616
rect 164344 157554 164372 160140
rect 164436 159202 164464 160140
rect 164528 159905 164556 160140
rect 164514 159896 164570 159905
rect 164514 159831 164570 159840
rect 164620 159780 164648 160140
rect 164528 159752 164648 159780
rect 164528 159576 164556 159752
rect 164528 159548 164648 159576
rect 164436 159174 164556 159202
rect 164424 159112 164476 159118
rect 164424 159054 164476 159060
rect 164332 157548 164384 157554
rect 164332 157490 164384 157496
rect 164436 157332 164464 159054
rect 164528 157536 164556 159174
rect 164620 158692 164648 159548
rect 164712 159118 164740 160140
rect 164804 159934 164832 160140
rect 164792 159928 164844 159934
rect 164792 159870 164844 159876
rect 164792 159792 164844 159798
rect 164792 159734 164844 159740
rect 164804 159322 164832 159734
rect 164792 159316 164844 159322
rect 164792 159258 164844 159264
rect 164792 159180 164844 159186
rect 164792 159122 164844 159128
rect 164700 159112 164752 159118
rect 164700 159054 164752 159060
rect 164804 158846 164832 159122
rect 164792 158840 164844 158846
rect 164792 158782 164844 158788
rect 164700 158704 164752 158710
rect 164620 158664 164700 158692
rect 164700 158646 164752 158652
rect 164790 158672 164846 158681
rect 164712 158409 164740 158646
rect 164790 158607 164846 158616
rect 164698 158400 164754 158409
rect 164698 158335 164754 158344
rect 164528 157508 164740 157536
rect 164606 157448 164662 157457
rect 164606 157383 164662 157392
rect 164436 157304 164556 157332
rect 164148 157004 164200 157010
rect 164148 156946 164200 156952
rect 164240 156528 164292 156534
rect 164240 156470 164292 156476
rect 164252 142866 164280 156470
rect 164424 155984 164476 155990
rect 164424 155926 164476 155932
rect 164240 142860 164292 142866
rect 164240 142802 164292 142808
rect 164436 141778 164464 155926
rect 164528 151094 164556 157304
rect 164516 151088 164568 151094
rect 164516 151030 164568 151036
rect 164424 141772 164476 141778
rect 164424 141714 164476 141720
rect 164436 138718 164464 141714
rect 164424 138712 164476 138718
rect 164424 138654 164476 138660
rect 163688 133204 163740 133210
rect 163688 133146 163740 133152
rect 164620 120766 164648 157383
rect 164712 155922 164740 157508
rect 164700 155916 164752 155922
rect 164700 155858 164752 155864
rect 164700 155780 164752 155786
rect 164700 155722 164752 155728
rect 164608 120760 164660 120766
rect 164608 120702 164660 120708
rect 163596 116612 163648 116618
rect 163596 116554 163648 116560
rect 164712 115258 164740 155722
rect 164700 115252 164752 115258
rect 164700 115194 164752 115200
rect 164804 15910 164832 158607
rect 164896 158370 164924 160140
rect 164884 158364 164936 158370
rect 164884 158306 164936 158312
rect 164884 157548 164936 157554
rect 164884 157490 164936 157496
rect 164896 157214 164924 157490
rect 164988 157321 165016 160140
rect 165080 159089 165108 160140
rect 165066 159080 165122 159089
rect 165066 159015 165122 159024
rect 165172 158681 165200 160140
rect 165158 158672 165214 158681
rect 165158 158607 165214 158616
rect 165172 158574 165200 158607
rect 165160 158568 165212 158574
rect 165160 158510 165212 158516
rect 165068 158364 165120 158370
rect 165068 158306 165120 158312
rect 165080 157622 165108 158306
rect 165068 157616 165120 157622
rect 165068 157558 165120 157564
rect 164974 157312 165030 157321
rect 164974 157247 165030 157256
rect 164884 157208 164936 157214
rect 164884 157150 164936 157156
rect 164792 15904 164844 15910
rect 164792 15846 164844 15852
rect 164896 13122 164924 157150
rect 165080 142154 165108 157558
rect 165264 156534 165292 160140
rect 165356 158982 165384 160140
rect 165448 159905 165476 160140
rect 165434 159896 165490 159905
rect 165434 159831 165490 159840
rect 165436 159792 165488 159798
rect 165436 159734 165488 159740
rect 165448 159662 165476 159734
rect 165436 159656 165488 159662
rect 165436 159598 165488 159604
rect 165344 158976 165396 158982
rect 165344 158918 165396 158924
rect 165252 156528 165304 156534
rect 165252 156470 165304 156476
rect 165356 155786 165384 158918
rect 165540 155990 165568 160140
rect 165632 159905 165660 160140
rect 165618 159896 165674 159905
rect 165618 159831 165674 159840
rect 165620 159792 165672 159798
rect 165620 159734 165672 159740
rect 165632 159361 165660 159734
rect 165618 159352 165674 159361
rect 165618 159287 165674 159296
rect 165724 158760 165752 160140
rect 165816 159934 165844 160140
rect 165804 159928 165856 159934
rect 165804 159870 165856 159876
rect 165804 159316 165856 159322
rect 165804 159258 165856 159264
rect 165632 158732 165752 158760
rect 165632 157894 165660 158732
rect 165710 158672 165766 158681
rect 165710 158607 165766 158616
rect 165620 157888 165672 157894
rect 165620 157830 165672 157836
rect 165632 157554 165660 157830
rect 165620 157548 165672 157554
rect 165620 157490 165672 157496
rect 165620 156936 165672 156942
rect 165620 156878 165672 156884
rect 165528 155984 165580 155990
rect 165528 155926 165580 155932
rect 165344 155780 165396 155786
rect 165344 155722 165396 155728
rect 164988 142126 165108 142154
rect 164988 100026 165016 142126
rect 164976 100020 165028 100026
rect 164976 99962 165028 99968
rect 165632 97374 165660 156878
rect 165724 149802 165752 158607
rect 165816 157758 165844 159258
rect 165908 159186 165936 160140
rect 165896 159180 165948 159186
rect 165896 159122 165948 159128
rect 165894 159080 165950 159089
rect 165894 159015 165950 159024
rect 165804 157752 165856 157758
rect 165804 157694 165856 157700
rect 165804 157004 165856 157010
rect 165804 156946 165856 156952
rect 165712 149796 165764 149802
rect 165712 149738 165764 149744
rect 165816 141438 165844 156946
rect 165908 148374 165936 159015
rect 166000 158438 166028 160140
rect 166092 159322 166120 160140
rect 166080 159316 166132 159322
rect 166080 159258 166132 159264
rect 166184 159254 166212 160140
rect 166276 159769 166304 160140
rect 166262 159760 166318 159769
rect 166262 159695 166318 159704
rect 166172 159248 166224 159254
rect 166172 159190 166224 159196
rect 166080 159180 166132 159186
rect 166080 159122 166132 159128
rect 166092 158681 166120 159122
rect 166078 158672 166134 158681
rect 166078 158607 166134 158616
rect 166080 158568 166132 158574
rect 166080 158510 166132 158516
rect 165988 158432 166040 158438
rect 165988 158374 166040 158380
rect 166000 151910 166028 158374
rect 166092 158273 166120 158510
rect 166078 158264 166134 158273
rect 166078 158199 166134 158208
rect 166080 157752 166132 157758
rect 166080 157694 166132 157700
rect 166092 157486 166120 157694
rect 166080 157480 166132 157486
rect 166080 157422 166132 157428
rect 166184 157010 166212 159190
rect 166172 157004 166224 157010
rect 166172 156946 166224 156952
rect 166276 156890 166304 159695
rect 166368 157049 166396 160140
rect 166354 157040 166410 157049
rect 166354 156975 166410 156984
rect 166092 156862 166304 156890
rect 165988 151904 166040 151910
rect 165988 151846 166040 151852
rect 165896 148368 165948 148374
rect 165896 148310 165948 148316
rect 165804 141432 165856 141438
rect 165804 141374 165856 141380
rect 166092 108322 166120 156862
rect 166460 151994 166488 160140
rect 166552 159905 166580 160140
rect 166538 159896 166594 159905
rect 166538 159831 166594 159840
rect 166552 157282 166580 159831
rect 166540 157276 166592 157282
rect 166540 157218 166592 157224
rect 166644 156942 166672 160140
rect 166632 156936 166684 156942
rect 166632 156878 166684 156884
rect 166184 151966 166488 151994
rect 166184 138009 166212 151966
rect 166264 151904 166316 151910
rect 166264 151846 166316 151852
rect 166170 138000 166226 138009
rect 166170 137935 166226 137944
rect 166184 137601 166212 137935
rect 166170 137592 166226 137601
rect 166170 137527 166226 137536
rect 166080 108316 166132 108322
rect 166080 108258 166132 108264
rect 165620 97368 165672 97374
rect 165620 97310 165672 97316
rect 164884 13116 164936 13122
rect 164884 13058 164936 13064
rect 166276 11762 166304 151846
rect 166736 142154 166764 160140
rect 166828 159905 166856 160140
rect 166814 159896 166870 159905
rect 166814 159831 166870 159840
rect 166920 159769 166948 160140
rect 166906 159760 166962 159769
rect 166906 159695 166962 159704
rect 166816 159316 166868 159322
rect 166816 159258 166868 159264
rect 166828 158953 166856 159258
rect 166920 159089 166948 159695
rect 166906 159080 166962 159089
rect 166906 159015 166962 159024
rect 166814 158944 166870 158953
rect 166814 158879 166870 158888
rect 166906 158264 166962 158273
rect 166906 158199 166962 158208
rect 166920 157729 166948 158199
rect 167012 157865 167040 160140
rect 167104 158710 167132 160140
rect 167092 158704 167144 158710
rect 167092 158646 167144 158652
rect 166998 157856 167054 157865
rect 166998 157791 167054 157800
rect 166906 157720 166962 157729
rect 166906 157655 166962 157664
rect 167000 156460 167052 156466
rect 167000 156402 167052 156408
rect 167012 144226 167040 156402
rect 167104 154574 167132 158646
rect 167196 157758 167224 160140
rect 167184 157752 167236 157758
rect 167184 157694 167236 157700
rect 167288 156777 167316 160140
rect 167380 158778 167408 160140
rect 167368 158772 167420 158778
rect 167368 158714 167420 158720
rect 167274 156768 167330 156777
rect 167274 156703 167330 156712
rect 167380 155394 167408 158714
rect 167472 156913 167500 160140
rect 167458 156904 167514 156913
rect 167458 156839 167514 156848
rect 167564 155530 167592 160140
rect 167656 159905 167684 160140
rect 167748 159934 167776 160140
rect 167840 159934 167868 160140
rect 167736 159928 167788 159934
rect 167642 159896 167698 159905
rect 167736 159870 167788 159876
rect 167828 159928 167880 159934
rect 167828 159870 167880 159876
rect 167642 159831 167698 159840
rect 167656 156670 167684 159831
rect 167840 159780 167868 159870
rect 167748 159752 167868 159780
rect 167932 159769 167960 160140
rect 167918 159760 167974 159769
rect 167644 156664 167696 156670
rect 167644 156606 167696 156612
rect 167564 155502 167684 155530
rect 167380 155366 167592 155394
rect 167104 154546 167408 154574
rect 167276 152516 167328 152522
rect 167276 152458 167328 152464
rect 167000 144220 167052 144226
rect 167000 144162 167052 144168
rect 166460 142126 166764 142154
rect 166460 139126 166488 142126
rect 167288 139194 167316 152458
rect 167380 142934 167408 154546
rect 167460 152448 167512 152454
rect 167460 152390 167512 152396
rect 167368 142928 167420 142934
rect 167368 142870 167420 142876
rect 167276 139188 167328 139194
rect 167276 139130 167328 139136
rect 166448 139120 166500 139126
rect 166448 139062 166500 139068
rect 166460 135930 166488 139062
rect 166448 135924 166500 135930
rect 166448 135866 166500 135872
rect 166356 112464 166408 112470
rect 166356 112406 166408 112412
rect 166264 11756 166316 11762
rect 166264 11698 166316 11704
rect 166080 3596 166132 3602
rect 166080 3538 166132 3544
rect 162124 3528 162176 3534
rect 162124 3470 162176 3476
rect 162492 3528 162544 3534
rect 162492 3470 162544 3476
rect 163504 3528 163556 3534
rect 163504 3470 163556 3476
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 162504 480 162532 3470
rect 163688 3256 163740 3262
rect 163688 3198 163740 3204
rect 163700 480 163728 3198
rect 164896 480 164924 3470
rect 166092 480 166120 3538
rect 166368 3262 166396 112406
rect 167472 105602 167500 152390
rect 167564 106962 167592 155366
rect 167656 152522 167684 155502
rect 167644 152516 167696 152522
rect 167644 152458 167696 152464
rect 167748 151814 167776 159752
rect 167918 159695 167974 159704
rect 167826 159624 167882 159633
rect 167826 159559 167882 159568
rect 167840 159225 167868 159559
rect 167826 159216 167882 159225
rect 167826 159151 167882 159160
rect 167828 158772 167880 158778
rect 167828 158714 167880 158720
rect 167840 158681 167868 158714
rect 167826 158672 167882 158681
rect 167826 158607 167882 158616
rect 167826 157992 167882 158001
rect 167826 157927 167882 157936
rect 167840 157894 167868 157927
rect 167828 157888 167880 157894
rect 167828 157830 167880 157836
rect 167932 152454 167960 159695
rect 168024 158817 168052 160140
rect 168010 158808 168066 158817
rect 168010 158743 168066 158752
rect 168012 158500 168064 158506
rect 168012 158442 168064 158448
rect 168024 156466 168052 158442
rect 168012 156460 168064 156466
rect 168012 156402 168064 156408
rect 167920 152448 167972 152454
rect 167920 152390 167972 152396
rect 167748 151786 167868 151814
rect 167644 139188 167696 139194
rect 167644 139130 167696 139136
rect 167656 127634 167684 139130
rect 167736 137828 167788 137834
rect 167736 137770 167788 137776
rect 167644 127628 167696 127634
rect 167644 127570 167696 127576
rect 167552 106956 167604 106962
rect 167552 106898 167604 106904
rect 167644 106956 167696 106962
rect 167644 106898 167696 106904
rect 167460 105596 167512 105602
rect 167460 105538 167512 105544
rect 167656 3534 167684 106898
rect 167748 37942 167776 137770
rect 167840 126274 167868 151786
rect 168116 142154 168144 160140
rect 168208 159905 168236 160140
rect 168194 159896 168250 159905
rect 168194 159831 168250 159840
rect 168208 156738 168236 159831
rect 168300 158506 168328 160140
rect 168288 158500 168340 158506
rect 168288 158442 168340 158448
rect 168286 158400 168342 158409
rect 168286 158335 168342 158344
rect 168300 157729 168328 158335
rect 168286 157720 168342 157729
rect 168286 157655 168342 157664
rect 168196 156732 168248 156738
rect 168196 156674 168248 156680
rect 168392 152454 168420 160140
rect 168484 159905 168512 160140
rect 168470 159896 168526 159905
rect 168470 159831 168526 159840
rect 168380 152448 168432 152454
rect 168380 152390 168432 152396
rect 168484 152266 168512 159831
rect 168576 158642 168604 160140
rect 168668 158681 168696 160140
rect 168760 158778 168788 160140
rect 168852 159769 168880 160140
rect 168838 159760 168894 159769
rect 168838 159695 168894 159704
rect 168748 158772 168800 158778
rect 168748 158714 168800 158720
rect 168654 158672 168710 158681
rect 168564 158636 168616 158642
rect 168654 158607 168710 158616
rect 168564 158578 168616 158584
rect 168760 158556 168788 158714
rect 168668 158528 168788 158556
rect 168564 158500 168616 158506
rect 168564 158442 168616 158448
rect 168576 158409 168604 158442
rect 168562 158400 168618 158409
rect 168562 158335 168618 158344
rect 168564 157888 168616 157894
rect 168562 157856 168564 157865
rect 168616 157856 168618 157865
rect 168562 157791 168618 157800
rect 168668 156806 168696 158528
rect 168748 158364 168800 158370
rect 168748 158306 168800 158312
rect 168656 156800 168708 156806
rect 168656 156742 168708 156748
rect 168564 155644 168616 155650
rect 168564 155586 168616 155592
rect 168392 152238 168512 152266
rect 168392 149138 168420 152238
rect 168392 149110 168512 149138
rect 168380 147348 168432 147354
rect 168380 147290 168432 147296
rect 168024 142126 168144 142154
rect 168024 137834 168052 142126
rect 168012 137828 168064 137834
rect 168012 137770 168064 137776
rect 167828 126268 167880 126274
rect 167828 126210 167880 126216
rect 167736 37936 167788 37942
rect 167736 37878 167788 37884
rect 167644 3528 167696 3534
rect 167644 3470 167696 3476
rect 166356 3256 166408 3262
rect 166356 3198 166408 3204
rect 167184 3052 167236 3058
rect 167184 2994 167236 3000
rect 167196 480 167224 2994
rect 168392 480 168420 147290
rect 168484 7614 168512 149110
rect 168576 147354 168604 155586
rect 168656 152652 168708 152658
rect 168656 152594 168708 152600
rect 168564 147348 168616 147354
rect 168564 147290 168616 147296
rect 168668 139369 168696 152594
rect 168654 139360 168710 139369
rect 168654 139295 168710 139304
rect 168564 139052 168616 139058
rect 168564 138994 168616 139000
rect 168576 135998 168604 138994
rect 168564 135992 168616 135998
rect 168564 135934 168616 135940
rect 168760 104174 168788 158306
rect 168944 157334 168972 160140
rect 169036 159905 169064 160140
rect 169022 159896 169078 159905
rect 169022 159831 169078 159840
rect 168852 157306 168972 157334
rect 168852 139097 168880 157306
rect 169036 156874 169064 159831
rect 169128 158545 169156 160140
rect 169114 158536 169170 158545
rect 169114 158471 169170 158480
rect 169024 156868 169076 156874
rect 169024 156810 169076 156816
rect 169220 152658 169248 160140
rect 169312 159633 169340 160140
rect 169298 159624 169354 159633
rect 169298 159559 169354 159568
rect 169312 158370 169340 159559
rect 169404 158681 169432 160140
rect 169496 159769 169524 160140
rect 169588 159905 169616 160140
rect 169574 159896 169630 159905
rect 169574 159831 169630 159840
rect 169482 159760 169538 159769
rect 169482 159695 169538 159704
rect 169390 158672 169446 158681
rect 169390 158607 169446 158616
rect 169300 158364 169352 158370
rect 169300 158306 169352 158312
rect 169392 158296 169444 158302
rect 169392 158238 169444 158244
rect 169404 158098 169432 158238
rect 169392 158092 169444 158098
rect 169392 158034 169444 158040
rect 169496 153950 169524 159695
rect 169484 153944 169536 153950
rect 169484 153886 169536 153892
rect 169208 152652 169260 152658
rect 169208 152594 169260 152600
rect 169588 152538 169616 159831
rect 169680 158409 169708 160140
rect 169772 159118 169800 160140
rect 169760 159112 169812 159118
rect 169760 159054 169812 159060
rect 169758 158944 169814 158953
rect 169758 158879 169814 158888
rect 169666 158400 169722 158409
rect 169666 158335 169722 158344
rect 169668 156460 169720 156466
rect 169668 156402 169720 156408
rect 168944 152510 169616 152538
rect 168944 141506 168972 152510
rect 169116 152448 169168 152454
rect 169116 152390 169168 152396
rect 168932 141500 168984 141506
rect 168932 141442 168984 141448
rect 169022 139360 169078 139369
rect 169022 139295 169078 139304
rect 168838 139088 168894 139097
rect 168838 139023 168894 139032
rect 169036 122126 169064 139295
rect 169128 139058 169156 152390
rect 169680 144265 169708 156402
rect 169772 155378 169800 158879
rect 169864 158794 169892 160140
rect 169956 159594 169984 160140
rect 169944 159588 169996 159594
rect 169944 159530 169996 159536
rect 169864 158766 169984 158794
rect 169850 158672 169906 158681
rect 169850 158607 169906 158616
rect 169760 155372 169812 155378
rect 169760 155314 169812 155320
rect 169666 144256 169722 144265
rect 169666 144191 169722 144200
rect 169206 139088 169262 139097
rect 169116 139052 169168 139058
rect 169206 139023 169262 139032
rect 169116 138994 169168 139000
rect 169220 130422 169248 139023
rect 169864 133278 169892 158607
rect 169956 157282 169984 158766
rect 169944 157276 169996 157282
rect 169944 157218 169996 157224
rect 169956 156602 169984 157218
rect 169944 156596 169996 156602
rect 169944 156538 169996 156544
rect 170048 145518 170076 160140
rect 170140 159633 170168 160140
rect 170232 159780 170260 160140
rect 170324 159905 170352 160140
rect 170416 159934 170444 160140
rect 170404 159928 170456 159934
rect 170310 159896 170366 159905
rect 170404 159870 170456 159876
rect 170310 159831 170366 159840
rect 170232 159752 170352 159780
rect 170220 159656 170272 159662
rect 170126 159624 170182 159633
rect 170324 159644 170352 159752
rect 170416 159746 170444 159870
rect 170508 159866 170536 160140
rect 170496 159860 170548 159866
rect 170496 159802 170548 159808
rect 170416 159718 170536 159746
rect 170324 159616 170444 159644
rect 170220 159598 170272 159604
rect 170126 159559 170182 159568
rect 170140 157350 170168 159559
rect 170232 158506 170260 159598
rect 170416 159322 170444 159616
rect 170404 159316 170456 159322
rect 170404 159258 170456 159264
rect 170220 158500 170272 158506
rect 170220 158442 170272 158448
rect 170404 157480 170456 157486
rect 170404 157422 170456 157428
rect 170128 157344 170180 157350
rect 170128 157286 170180 157292
rect 170036 145512 170088 145518
rect 170036 145454 170088 145460
rect 169852 133272 169904 133278
rect 169852 133214 169904 133220
rect 169208 130416 169260 130422
rect 169208 130358 169260 130364
rect 169024 122120 169076 122126
rect 169024 122062 169076 122068
rect 168748 104168 168800 104174
rect 168748 104110 168800 104116
rect 170416 8974 170444 157422
rect 170508 157010 170536 159718
rect 170600 159322 170628 160140
rect 170692 159769 170720 160140
rect 170678 159760 170734 159769
rect 170678 159695 170734 159704
rect 170784 159610 170812 160140
rect 170876 159934 170904 160140
rect 170968 159934 170996 160140
rect 171060 159939 171088 160140
rect 170864 159928 170916 159934
rect 170864 159870 170916 159876
rect 170956 159928 171008 159934
rect 170956 159870 171008 159876
rect 171046 159930 171102 159939
rect 170692 159582 170812 159610
rect 170588 159316 170640 159322
rect 170588 159258 170640 159264
rect 170588 159112 170640 159118
rect 170588 159054 170640 159060
rect 170496 157004 170548 157010
rect 170496 156946 170548 156952
rect 170496 145512 170548 145518
rect 170496 145454 170548 145460
rect 170508 129130 170536 145454
rect 170496 129124 170548 129130
rect 170496 129066 170548 129072
rect 170600 60042 170628 159054
rect 170692 156466 170720 159582
rect 170772 159520 170824 159526
rect 170772 159462 170824 159468
rect 170784 158914 170812 159462
rect 170772 158908 170824 158914
rect 170772 158850 170824 158856
rect 170680 156460 170732 156466
rect 170680 156402 170732 156408
rect 170876 142154 170904 159870
rect 171046 159865 171102 159874
rect 171152 159769 171180 160140
rect 171138 159760 171194 159769
rect 171048 159724 171100 159730
rect 171138 159695 171194 159704
rect 171048 159666 171100 159672
rect 170954 159352 171010 159361
rect 170954 159287 170956 159296
rect 171008 159287 171010 159296
rect 170956 159258 171008 159264
rect 170968 146946 170996 159258
rect 171060 158370 171088 159666
rect 171048 158364 171100 158370
rect 171048 158306 171100 158312
rect 171060 157486 171088 158306
rect 171048 157480 171100 157486
rect 171048 157422 171100 157428
rect 171046 157312 171102 157321
rect 171046 157247 171048 157256
rect 171100 157247 171102 157256
rect 171048 157218 171100 157224
rect 171048 157004 171100 157010
rect 171048 156946 171100 156952
rect 170956 146940 171008 146946
rect 170956 146882 171008 146888
rect 170784 142126 170904 142154
rect 170784 123554 170812 142126
rect 170772 123548 170824 123554
rect 170772 123490 170824 123496
rect 171060 102814 171088 156946
rect 171152 152590 171180 159695
rect 171244 159662 171272 160140
rect 171232 159656 171284 159662
rect 171232 159598 171284 159604
rect 171336 159594 171364 160140
rect 171428 159934 171456 160140
rect 171416 159928 171468 159934
rect 171520 159905 171548 160140
rect 171416 159870 171468 159876
rect 171506 159896 171562 159905
rect 171506 159831 171562 159840
rect 171612 159610 171640 160140
rect 171704 159633 171732 160140
rect 171324 159588 171376 159594
rect 171324 159530 171376 159536
rect 171520 159582 171640 159610
rect 171690 159624 171746 159633
rect 171416 159452 171468 159458
rect 171416 159394 171468 159400
rect 171232 159316 171284 159322
rect 171232 159258 171284 159264
rect 171244 158846 171272 159258
rect 171428 159050 171456 159394
rect 171520 159225 171548 159582
rect 171796 159594 171824 160140
rect 171888 159934 171916 160140
rect 171980 159939 172008 160140
rect 171876 159928 171928 159934
rect 171876 159870 171928 159876
rect 171966 159930 172022 159939
rect 171966 159865 172022 159874
rect 171968 159792 172020 159798
rect 172072 159769 172100 160140
rect 171968 159734 172020 159740
rect 172058 159760 172114 159769
rect 171876 159656 171928 159662
rect 171876 159598 171928 159604
rect 171690 159559 171746 159568
rect 171784 159588 171836 159594
rect 171784 159530 171836 159536
rect 171600 159520 171652 159526
rect 171600 159462 171652 159468
rect 171612 159361 171640 159462
rect 171692 159452 171744 159458
rect 171692 159394 171744 159400
rect 171598 159352 171654 159361
rect 171598 159287 171654 159296
rect 171506 159216 171562 159225
rect 171506 159151 171562 159160
rect 171324 159044 171376 159050
rect 171324 158986 171376 158992
rect 171416 159044 171468 159050
rect 171416 158986 171468 158992
rect 171336 158846 171364 158986
rect 171506 158944 171562 158953
rect 171506 158879 171562 158888
rect 171232 158840 171284 158846
rect 171232 158782 171284 158788
rect 171324 158840 171376 158846
rect 171324 158782 171376 158788
rect 171324 158636 171376 158642
rect 171324 158578 171376 158584
rect 171230 155952 171286 155961
rect 171230 155887 171286 155896
rect 171140 152584 171192 152590
rect 171140 152526 171192 152532
rect 171244 147674 171272 155887
rect 171152 147646 171272 147674
rect 171048 102808 171100 102814
rect 171048 102750 171100 102756
rect 170588 60036 170640 60042
rect 170588 59978 170640 59984
rect 171152 16574 171180 147646
rect 171336 124982 171364 158578
rect 171520 142154 171548 158879
rect 171612 158642 171640 159287
rect 171704 158710 171732 159394
rect 171692 158704 171744 158710
rect 171692 158646 171744 158652
rect 171600 158636 171652 158642
rect 171600 158578 171652 158584
rect 171598 158536 171654 158545
rect 171598 158471 171654 158480
rect 171612 157146 171640 158471
rect 171796 158250 171824 159530
rect 171888 159390 171916 159598
rect 171876 159384 171928 159390
rect 171876 159326 171928 159332
rect 171874 158672 171930 158681
rect 171980 158642 172008 159734
rect 172058 159695 172114 159704
rect 172164 158794 172192 160140
rect 172072 158766 172192 158794
rect 171874 158607 171930 158616
rect 171968 158636 172020 158642
rect 171704 158222 171824 158250
rect 171600 157140 171652 157146
rect 171600 157082 171652 157088
rect 171704 154574 171732 158222
rect 171784 158160 171836 158166
rect 171784 158102 171836 158108
rect 171796 157826 171824 158102
rect 171784 157820 171836 157826
rect 171784 157762 171836 157768
rect 171704 154546 171824 154574
rect 171692 152516 171744 152522
rect 171692 152458 171744 152464
rect 171428 142126 171548 142154
rect 171428 127702 171456 142126
rect 171704 138786 171732 152458
rect 171796 147674 171824 154546
rect 171888 152522 171916 158607
rect 171968 158578 172020 158584
rect 172072 158522 172100 158766
rect 171980 158494 172100 158522
rect 172150 158536 172206 158545
rect 171980 155854 172008 158494
rect 172150 158471 172206 158480
rect 171968 155848 172020 155854
rect 171968 155790 172020 155796
rect 171876 152516 171928 152522
rect 171876 152458 171928 152464
rect 171796 147646 171916 147674
rect 171692 138780 171744 138786
rect 171692 138722 171744 138728
rect 171782 131200 171838 131209
rect 171782 131135 171838 131144
rect 171416 127696 171468 127702
rect 171416 127638 171468 127644
rect 171324 124976 171376 124982
rect 171324 124918 171376 124924
rect 171152 16546 171732 16574
rect 170404 8968 170456 8974
rect 170404 8910 170456 8916
rect 168472 7608 168524 7614
rect 168472 7550 168524 7556
rect 171416 4072 171468 4078
rect 171416 4014 171468 4020
rect 170772 3528 170824 3534
rect 170772 3470 170824 3476
rect 169576 3460 169628 3466
rect 169576 3402 169628 3408
rect 169588 480 169616 3402
rect 170784 480 170812 3470
rect 171428 3058 171456 4014
rect 171704 3482 171732 16546
rect 171796 4078 171824 131135
rect 171888 101454 171916 147646
rect 172164 143002 172192 158471
rect 172256 152318 172284 160140
rect 172348 158681 172376 160140
rect 172440 159050 172468 160140
rect 172428 159044 172480 159050
rect 172428 158986 172480 158992
rect 172334 158672 172390 158681
rect 172334 158607 172390 158616
rect 172428 158636 172480 158642
rect 172428 158578 172480 158584
rect 172336 152584 172388 152590
rect 172336 152526 172388 152532
rect 172244 152312 172296 152318
rect 172244 152254 172296 152260
rect 172152 142996 172204 143002
rect 172152 142938 172204 142944
rect 172348 131782 172376 152526
rect 172440 142089 172468 158578
rect 172532 157321 172560 160140
rect 172624 159905 172652 160140
rect 172610 159896 172666 159905
rect 172716 159866 172744 160140
rect 172610 159831 172666 159840
rect 172704 159860 172756 159866
rect 172704 159802 172756 159808
rect 172702 159760 172758 159769
rect 172612 159724 172664 159730
rect 172702 159695 172758 159704
rect 172612 159666 172664 159672
rect 172624 158982 172652 159666
rect 172612 158976 172664 158982
rect 172612 158918 172664 158924
rect 172716 157334 172744 159695
rect 172808 158964 172836 160140
rect 172900 159905 172928 160140
rect 172886 159896 172942 159905
rect 172886 159831 172942 159840
rect 172888 159792 172940 159798
rect 172888 159734 172940 159740
rect 172900 159225 172928 159734
rect 172886 159216 172942 159225
rect 172886 159151 172942 159160
rect 172808 158936 172928 158964
rect 172518 157312 172574 157321
rect 172716 157306 172836 157334
rect 172518 157247 172574 157256
rect 172808 155582 172836 157306
rect 172796 155576 172848 155582
rect 172796 155518 172848 155524
rect 172900 154170 172928 158936
rect 172992 156466 173020 160140
rect 173084 158681 173112 160140
rect 173176 159769 173204 160140
rect 173162 159760 173218 159769
rect 173162 159695 173218 159704
rect 173070 158672 173126 158681
rect 173070 158607 173126 158616
rect 173176 157334 173204 159695
rect 173084 157306 173204 157334
rect 172980 156460 173032 156466
rect 172980 156402 173032 156408
rect 172992 155446 173020 156402
rect 172980 155440 173032 155446
rect 172980 155382 173032 155388
rect 172808 154142 172928 154170
rect 172808 152386 172836 154142
rect 173084 152538 173112 157306
rect 173268 154086 173296 160140
rect 173360 159866 173388 160140
rect 173452 159905 173480 160140
rect 173438 159896 173494 159905
rect 173348 159860 173400 159866
rect 173438 159831 173494 159840
rect 173348 159802 173400 159808
rect 173348 159724 173400 159730
rect 173348 159666 173400 159672
rect 173360 154222 173388 159666
rect 173348 154216 173400 154222
rect 173348 154158 173400 154164
rect 173256 154080 173308 154086
rect 173256 154022 173308 154028
rect 173164 152720 173216 152726
rect 173164 152662 173216 152668
rect 172900 152510 173112 152538
rect 172796 152380 172848 152386
rect 172796 152322 172848 152328
rect 172520 149524 172572 149530
rect 172520 149466 172572 149472
rect 172426 142080 172482 142089
rect 172426 142015 172482 142024
rect 172440 140185 172468 142015
rect 172426 140176 172482 140185
rect 172426 140111 172482 140120
rect 172336 131776 172388 131782
rect 172336 131718 172388 131724
rect 171876 101448 171928 101454
rect 171876 101390 171928 101396
rect 172532 16574 172560 149466
rect 172900 145654 172928 152510
rect 172980 152448 173032 152454
rect 172980 152390 173032 152396
rect 172992 147257 173020 152390
rect 172978 147248 173034 147257
rect 172978 147183 173034 147192
rect 172888 145648 172940 145654
rect 172888 145590 172940 145596
rect 173176 137290 173204 152662
rect 173452 144294 173480 159831
rect 173544 157078 173572 160140
rect 173532 157072 173584 157078
rect 173532 157014 173584 157020
rect 173636 152454 173664 160140
rect 173728 159905 173756 160140
rect 173714 159896 173770 159905
rect 173714 159831 173770 159840
rect 173624 152448 173676 152454
rect 173624 152390 173676 152396
rect 173728 148442 173756 159831
rect 173820 152726 173848 160140
rect 173912 158681 173940 160140
rect 174004 159633 174032 160140
rect 173990 159624 174046 159633
rect 173990 159559 174046 159568
rect 173992 159452 174044 159458
rect 173992 159394 174044 159400
rect 174004 159225 174032 159394
rect 173990 159216 174046 159225
rect 173990 159151 174046 159160
rect 174096 158794 174124 160140
rect 174188 159089 174216 160140
rect 174280 159905 174308 160140
rect 174372 159934 174400 160140
rect 174464 159934 174492 160140
rect 174556 159939 174584 160140
rect 174360 159928 174412 159934
rect 174266 159896 174322 159905
rect 174360 159870 174412 159876
rect 174452 159928 174504 159934
rect 174452 159870 174504 159876
rect 174542 159930 174598 159939
rect 174542 159865 174598 159874
rect 174266 159831 174322 159840
rect 174174 159080 174230 159089
rect 174174 159015 174230 159024
rect 174096 158766 174216 158794
rect 173898 158672 173954 158681
rect 173898 158607 173954 158616
rect 174084 158636 174136 158642
rect 174084 158578 174136 158584
rect 173808 152720 173860 152726
rect 173808 152662 173860 152668
rect 173716 148436 173768 148442
rect 173716 148378 173768 148384
rect 173898 146296 173954 146305
rect 173898 146231 173954 146240
rect 173440 144288 173492 144294
rect 173440 144230 173492 144236
rect 173164 137284 173216 137290
rect 173164 137226 173216 137232
rect 172532 16546 172744 16574
rect 171784 4072 171836 4078
rect 171784 4014 171836 4020
rect 171704 3454 172008 3482
rect 171416 3052 171468 3058
rect 171416 2994 171468 3000
rect 171980 480 172008 3454
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 146231
rect 174096 112470 174124 158578
rect 174188 155310 174216 158766
rect 174176 155304 174228 155310
rect 174176 155246 174228 155252
rect 174188 155038 174216 155246
rect 174176 155032 174228 155038
rect 174176 154974 174228 154980
rect 174280 154154 174308 159831
rect 174452 159724 174504 159730
rect 174452 159666 174504 159672
rect 174360 159656 174412 159662
rect 174360 159598 174412 159604
rect 174372 157729 174400 159598
rect 174464 157865 174492 159666
rect 174450 157856 174506 157865
rect 174450 157791 174506 157800
rect 174358 157720 174414 157729
rect 174358 157655 174414 157664
rect 174268 154148 174320 154154
rect 174268 154090 174320 154096
rect 174648 153950 174676 160140
rect 174740 159934 174768 160140
rect 174832 159934 174860 160140
rect 174728 159928 174780 159934
rect 174728 159870 174780 159876
rect 174820 159928 174872 159934
rect 174820 159870 174872 159876
rect 174818 159760 174874 159769
rect 174924 159746 174952 160140
rect 175016 159939 175044 160140
rect 175002 159930 175058 159939
rect 175002 159865 175058 159874
rect 175108 159769 175136 160140
rect 175094 159760 175150 159769
rect 174924 159718 175044 159746
rect 174818 159695 174874 159704
rect 174726 159624 174782 159633
rect 174726 159559 174782 159568
rect 174740 159390 174768 159559
rect 174728 159384 174780 159390
rect 174728 159326 174780 159332
rect 174728 159044 174780 159050
rect 174728 158986 174780 158992
rect 174740 158778 174768 158986
rect 174728 158772 174780 158778
rect 174728 158714 174780 158720
rect 174832 158642 174860 159695
rect 174912 159656 174964 159662
rect 174912 159598 174964 159604
rect 174820 158636 174872 158642
rect 174820 158578 174872 158584
rect 174818 158536 174874 158545
rect 174818 158471 174874 158480
rect 174728 154624 174780 154630
rect 174728 154566 174780 154572
rect 174636 153944 174688 153950
rect 174636 153886 174688 153892
rect 174544 151632 174596 151638
rect 174544 151574 174596 151580
rect 174084 112464 174136 112470
rect 174084 112406 174136 112412
rect 174556 3466 174584 151574
rect 174634 143440 174690 143449
rect 174634 143375 174690 143384
rect 174648 143002 174676 143375
rect 174636 142996 174688 143002
rect 174636 142938 174688 142944
rect 174648 3534 174676 142938
rect 174740 106962 174768 154566
rect 174832 145586 174860 158471
rect 174924 154290 174952 159598
rect 175016 158642 175044 159718
rect 175094 159695 175150 159704
rect 175096 159384 175148 159390
rect 175096 159326 175148 159332
rect 175004 158636 175056 158642
rect 175004 158578 175056 158584
rect 175002 158536 175058 158545
rect 175002 158471 175058 158480
rect 174912 154284 174964 154290
rect 174912 154226 174964 154232
rect 175016 150142 175044 158471
rect 175004 150136 175056 150142
rect 175004 150078 175056 150084
rect 175016 147674 175044 150078
rect 174924 147646 175044 147674
rect 174820 145580 174872 145586
rect 174820 145522 174872 145528
rect 174924 142154 174952 147646
rect 175108 147082 175136 159326
rect 175200 155582 175228 160140
rect 175292 159322 175320 160140
rect 175280 159316 175332 159322
rect 175280 159258 175332 159264
rect 175280 159044 175332 159050
rect 175280 158986 175332 158992
rect 175292 158409 175320 158986
rect 175384 158545 175412 160140
rect 175476 158710 175504 160140
rect 175464 158704 175516 158710
rect 175464 158646 175516 158652
rect 175464 158568 175516 158574
rect 175370 158536 175426 158545
rect 175464 158510 175516 158516
rect 175370 158471 175426 158480
rect 175278 158400 175334 158409
rect 175278 158335 175334 158344
rect 175476 157334 175504 158510
rect 175292 157306 175504 157334
rect 175568 157334 175596 160140
rect 175660 159050 175688 160140
rect 175648 159044 175700 159050
rect 175648 158986 175700 158992
rect 175752 158930 175780 160140
rect 175660 158902 175780 158930
rect 175660 158681 175688 158902
rect 175740 158772 175792 158778
rect 175740 158714 175792 158720
rect 175646 158672 175702 158681
rect 175646 158607 175702 158616
rect 175568 157306 175688 157334
rect 175188 155576 175240 155582
rect 175188 155518 175240 155524
rect 175200 154630 175228 155518
rect 175188 154624 175240 154630
rect 175188 154566 175240 154572
rect 175096 147076 175148 147082
rect 175096 147018 175148 147024
rect 174832 142126 174952 142154
rect 174832 117978 174860 142126
rect 174820 117972 174872 117978
rect 174820 117914 174872 117920
rect 174728 106956 174780 106962
rect 174728 106898 174780 106904
rect 174636 3528 174688 3534
rect 174636 3470 174688 3476
rect 174544 3460 174596 3466
rect 174544 3402 174596 3408
rect 175292 3262 175320 157306
rect 175372 156392 175424 156398
rect 175372 156334 175424 156340
rect 175384 155650 175412 156334
rect 175372 155644 175424 155650
rect 175372 155586 175424 155592
rect 175372 155508 175424 155514
rect 175372 155450 175424 155456
rect 175384 16574 175412 155450
rect 175556 152516 175608 152522
rect 175556 152458 175608 152464
rect 175464 152448 175516 152454
rect 175464 152390 175516 152396
rect 175476 144566 175504 152390
rect 175568 144702 175596 152458
rect 175660 151638 175688 157306
rect 175752 155514 175780 158714
rect 175740 155508 175792 155514
rect 175740 155450 175792 155456
rect 175648 151632 175700 151638
rect 175648 151574 175700 151580
rect 175844 149530 175872 160140
rect 175936 159905 175964 160140
rect 175922 159896 175978 159905
rect 175922 159831 175978 159840
rect 175936 158273 175964 159831
rect 176028 158778 176056 160140
rect 176120 159458 176148 160140
rect 176108 159452 176160 159458
rect 176108 159394 176160 159400
rect 176108 159316 176160 159322
rect 176108 159258 176160 159264
rect 176120 159225 176148 159258
rect 176106 159216 176162 159225
rect 176106 159151 176162 159160
rect 176016 158772 176068 158778
rect 176016 158714 176068 158720
rect 176014 158672 176070 158681
rect 176014 158607 176070 158616
rect 175922 158264 175978 158273
rect 175922 158199 175978 158208
rect 176028 158030 176056 158607
rect 176108 158092 176160 158098
rect 176108 158034 176160 158040
rect 176016 158024 176068 158030
rect 176016 157966 176068 157972
rect 176028 157894 176056 157966
rect 176016 157888 176068 157894
rect 176016 157830 176068 157836
rect 175832 149524 175884 149530
rect 175832 149466 175884 149472
rect 176120 147674 176148 158034
rect 176212 152522 176240 160140
rect 176304 159610 176332 160140
rect 176396 159769 176424 160140
rect 176382 159760 176438 159769
rect 176382 159695 176438 159704
rect 176304 159582 176424 159610
rect 176292 159452 176344 159458
rect 176292 159394 176344 159400
rect 176304 158098 176332 159394
rect 176396 158846 176424 159582
rect 176384 158840 176436 158846
rect 176384 158782 176436 158788
rect 176384 158704 176436 158710
rect 176384 158646 176436 158652
rect 176292 158092 176344 158098
rect 176292 158034 176344 158040
rect 176292 157888 176344 157894
rect 176292 157830 176344 157836
rect 176304 156126 176332 157830
rect 176396 156398 176424 158646
rect 176384 156392 176436 156398
rect 176384 156334 176436 156340
rect 176292 156120 176344 156126
rect 176292 156062 176344 156068
rect 176292 154216 176344 154222
rect 176292 154158 176344 154164
rect 176304 153678 176332 154158
rect 176292 153672 176344 153678
rect 176292 153614 176344 153620
rect 176200 152516 176252 152522
rect 176200 152458 176252 152464
rect 176488 152454 176516 160140
rect 176580 156602 176608 160140
rect 176672 158914 176700 160140
rect 176660 158908 176712 158914
rect 176660 158850 176712 158856
rect 176568 156596 176620 156602
rect 176568 156538 176620 156544
rect 176476 152448 176528 152454
rect 176476 152390 176528 152396
rect 176672 151774 176700 158850
rect 176660 151768 176712 151774
rect 176660 151710 176712 151716
rect 175936 147646 176148 147674
rect 175556 144696 175608 144702
rect 175556 144638 175608 144644
rect 175464 144560 175516 144566
rect 175464 144502 175516 144508
rect 175936 23526 175964 147646
rect 176568 144696 176620 144702
rect 176568 144638 176620 144644
rect 176476 144560 176528 144566
rect 176476 144502 176528 144508
rect 176488 144226 176516 144502
rect 176476 144220 176528 144226
rect 176476 144162 176528 144168
rect 176488 99346 176516 144162
rect 176580 144022 176608 144638
rect 176568 144016 176620 144022
rect 176568 143958 176620 143964
rect 176476 99340 176528 99346
rect 176476 99282 176528 99288
rect 175924 23520 175976 23526
rect 175924 23462 175976 23468
rect 175384 16546 175504 16574
rect 175280 3256 175332 3262
rect 175280 3198 175332 3204
rect 175476 480 175504 16546
rect 176580 8294 176608 143958
rect 176764 142866 176792 160140
rect 176856 156602 176884 160140
rect 176948 157865 176976 160140
rect 176934 157856 176990 157865
rect 176934 157791 176990 157800
rect 176844 156596 176896 156602
rect 176844 156538 176896 156544
rect 176844 152516 176896 152522
rect 176844 152458 176896 152464
rect 176856 144430 176884 152458
rect 176844 144424 176896 144430
rect 176844 144366 176896 144372
rect 177040 143614 177068 160140
rect 177132 157690 177160 160140
rect 177120 157684 177172 157690
rect 177120 157626 177172 157632
rect 177224 157457 177252 160140
rect 177210 157448 177266 157457
rect 177210 157383 177266 157392
rect 177028 143608 177080 143614
rect 177028 143550 177080 143556
rect 177316 142934 177344 160140
rect 177408 158098 177436 160140
rect 177396 158092 177448 158098
rect 177396 158034 177448 158040
rect 177408 146334 177436 158034
rect 177500 149870 177528 160140
rect 177592 152522 177620 160140
rect 177684 157826 177712 160140
rect 177672 157820 177724 157826
rect 177672 157762 177724 157768
rect 177684 152658 177712 157762
rect 177776 157457 177804 160140
rect 177868 157729 177896 160140
rect 177960 158234 177988 160140
rect 177948 158228 178000 158234
rect 177948 158170 178000 158176
rect 177854 157720 177910 157729
rect 177854 157655 177910 157664
rect 177762 157448 177818 157457
rect 177762 157383 177818 157392
rect 177960 155310 177988 158170
rect 177948 155304 178000 155310
rect 177948 155246 178000 155252
rect 178052 155242 178080 160140
rect 178144 159905 178172 160140
rect 178130 159896 178186 159905
rect 178130 159831 178186 159840
rect 178040 155236 178092 155242
rect 178040 155178 178092 155184
rect 177672 152652 177724 152658
rect 177672 152594 177724 152600
rect 177580 152516 177632 152522
rect 177580 152458 177632 152464
rect 177488 149864 177540 149870
rect 177488 149806 177540 149812
rect 177500 147674 177528 149806
rect 177500 147646 177712 147674
rect 177396 146328 177448 146334
rect 177396 146270 177448 146276
rect 177304 142928 177356 142934
rect 177304 142870 177356 142876
rect 176752 142860 176804 142866
rect 176752 142802 176804 142808
rect 177684 104174 177712 147646
rect 177948 144424 178000 144430
rect 177948 144366 178000 144372
rect 177764 144288 177816 144294
rect 177764 144230 177816 144236
rect 177776 143614 177804 144230
rect 177764 143608 177816 143614
rect 177764 143550 177816 143556
rect 177672 104168 177724 104174
rect 177672 104110 177724 104116
rect 177776 66910 177804 143550
rect 177856 143132 177908 143138
rect 177856 143074 177908 143080
rect 177868 142934 177896 143074
rect 177856 142928 177908 142934
rect 177856 142870 177908 142876
rect 177764 66904 177816 66910
rect 177764 66846 177816 66852
rect 177868 60042 177896 142870
rect 177856 60036 177908 60042
rect 177856 59978 177908 59984
rect 176660 23520 176712 23526
rect 176660 23462 176712 23468
rect 176568 8288 176620 8294
rect 176568 8230 176620 8236
rect 176672 480 176700 23462
rect 177960 15910 177988 144366
rect 178144 138014 178172 159831
rect 178236 158001 178264 160140
rect 178222 157992 178278 158001
rect 178222 157927 178278 157936
rect 178328 157457 178356 160140
rect 178420 157865 178448 160140
rect 178512 159934 178540 160140
rect 178500 159928 178552 159934
rect 178500 159870 178552 159876
rect 178512 158574 178540 159870
rect 178500 158568 178552 158574
rect 178500 158510 178552 158516
rect 178406 157856 178462 157865
rect 178406 157791 178462 157800
rect 178314 157448 178370 157457
rect 178314 157383 178370 157392
rect 178604 153814 178632 160140
rect 178696 159769 178724 160140
rect 178682 159760 178738 159769
rect 178682 159695 178738 159704
rect 178592 153808 178644 153814
rect 178592 153750 178644 153756
rect 178696 152998 178724 159695
rect 178788 156806 178816 160140
rect 178776 156800 178828 156806
rect 178776 156742 178828 156748
rect 178880 153882 178908 160140
rect 178972 159769 179000 160140
rect 178958 159760 179014 159769
rect 178958 159695 179014 159704
rect 178972 157729 179000 159695
rect 178958 157720 179014 157729
rect 178958 157655 179014 157664
rect 179064 157010 179092 160140
rect 179052 157004 179104 157010
rect 179052 156946 179104 156952
rect 178868 153876 178920 153882
rect 178868 153818 178920 153824
rect 178684 152992 178736 152998
rect 178684 152934 178736 152940
rect 179156 149802 179184 160140
rect 179248 158681 179276 160140
rect 179234 158672 179290 158681
rect 179234 158607 179290 158616
rect 179234 157856 179290 157865
rect 179234 157791 179290 157800
rect 179144 149796 179196 149802
rect 179144 149738 179196 149744
rect 178052 137986 178172 138014
rect 178052 108322 178080 137986
rect 178040 108316 178092 108322
rect 178040 108258 178092 108264
rect 179248 33794 179276 157791
rect 179340 155446 179368 160140
rect 179432 157334 179460 160140
rect 179524 157729 179552 160140
rect 179510 157720 179566 157729
rect 179510 157655 179566 157664
rect 179432 157306 179552 157334
rect 179420 156120 179472 156126
rect 179420 156062 179472 156068
rect 179328 155440 179380 155446
rect 179328 155382 179380 155388
rect 179328 142860 179380 142866
rect 179328 142802 179380 142808
rect 179236 33788 179288 33794
rect 179236 33730 179288 33736
rect 177948 15904 178000 15910
rect 177948 15846 178000 15852
rect 177856 8288 177908 8294
rect 177856 8230 177908 8236
rect 177868 480 177896 8230
rect 179340 3806 179368 142802
rect 179432 16574 179460 156062
rect 179524 148238 179552 157306
rect 179616 156874 179644 160140
rect 179604 156868 179656 156874
rect 179604 156810 179656 156816
rect 179512 148232 179564 148238
rect 179512 148174 179564 148180
rect 179708 146878 179736 160140
rect 179800 158681 179828 160140
rect 179786 158672 179842 158681
rect 179786 158607 179842 158616
rect 179892 155106 179920 160140
rect 179984 157457 180012 160140
rect 180076 159905 180104 160140
rect 180062 159896 180118 159905
rect 180062 159831 180118 159840
rect 180064 159656 180116 159662
rect 180064 159598 180116 159604
rect 180076 158982 180104 159598
rect 180064 158976 180116 158982
rect 180064 158918 180116 158924
rect 179970 157448 180026 157457
rect 179970 157383 180026 157392
rect 180168 155650 180196 160140
rect 180156 155644 180208 155650
rect 180156 155586 180208 155592
rect 179880 155100 179932 155106
rect 179880 155042 179932 155048
rect 180260 151366 180288 160140
rect 180352 157457 180380 160140
rect 180338 157448 180394 157457
rect 180338 157383 180394 157392
rect 180444 154154 180472 160140
rect 180536 158166 180564 160140
rect 180628 159905 180656 160140
rect 180614 159896 180670 159905
rect 180614 159831 180670 159840
rect 180524 158160 180576 158166
rect 180524 158102 180576 158108
rect 180524 157956 180576 157962
rect 180524 157898 180576 157904
rect 180432 154148 180484 154154
rect 180432 154090 180484 154096
rect 180536 154018 180564 157898
rect 180628 157842 180656 159831
rect 180720 157962 180748 160140
rect 180812 158098 180840 160140
rect 180904 159633 180932 160140
rect 180890 159624 180946 159633
rect 180890 159559 180946 159568
rect 180800 158092 180852 158098
rect 180800 158034 180852 158040
rect 180904 158001 180932 159559
rect 180890 157992 180946 158001
rect 180708 157956 180760 157962
rect 180890 157927 180946 157936
rect 180708 157898 180760 157904
rect 180628 157814 180748 157842
rect 180614 157720 180670 157729
rect 180614 157655 180670 157664
rect 180524 154012 180576 154018
rect 180524 153954 180576 153960
rect 180248 151360 180300 151366
rect 180248 151302 180300 151308
rect 179696 146872 179748 146878
rect 179696 146814 179748 146820
rect 180064 146328 180116 146334
rect 180064 146270 180116 146276
rect 179432 16546 180012 16574
rect 179328 3800 179380 3806
rect 179328 3742 179380 3748
rect 179984 3482 180012 16546
rect 180076 3602 180104 146270
rect 180628 137290 180656 157655
rect 180616 137284 180668 137290
rect 180616 137226 180668 137232
rect 180154 136640 180210 136649
rect 180154 136575 180210 136584
rect 180168 3670 180196 136575
rect 180720 93226 180748 157814
rect 180996 152794 181024 160140
rect 180984 152788 181036 152794
rect 180984 152730 181036 152736
rect 181088 151502 181116 160140
rect 181180 159905 181208 160140
rect 181166 159896 181222 159905
rect 181166 159831 181222 159840
rect 181180 152386 181208 159831
rect 181168 152380 181220 152386
rect 181168 152322 181220 152328
rect 181076 151496 181128 151502
rect 181076 151438 181128 151444
rect 181272 151434 181300 160140
rect 181364 158030 181392 160140
rect 181352 158024 181404 158030
rect 181352 157966 181404 157972
rect 181456 157729 181484 160140
rect 181442 157720 181498 157729
rect 181352 157684 181404 157690
rect 181442 157655 181498 157664
rect 181352 157626 181404 157632
rect 181364 157334 181392 157626
rect 181364 157306 181484 157334
rect 181260 151428 181312 151434
rect 181260 151370 181312 151376
rect 180800 99340 180852 99346
rect 180800 99282 180852 99288
rect 180708 93220 180760 93226
rect 180708 93162 180760 93168
rect 180812 16574 180840 99282
rect 180812 16546 181024 16574
rect 180156 3664 180208 3670
rect 180156 3606 180208 3612
rect 180064 3596 180116 3602
rect 180064 3538 180116 3544
rect 179984 3454 180288 3482
rect 179052 3256 179104 3262
rect 179052 3198 179104 3204
rect 179064 480 179092 3198
rect 180260 480 180288 3454
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 3058 181484 157306
rect 181548 153626 181576 160140
rect 181640 154358 181668 160140
rect 181732 157457 181760 160140
rect 181718 157448 181774 157457
rect 181718 157383 181774 157392
rect 181628 154352 181680 154358
rect 181628 154294 181680 154300
rect 181548 153598 181668 153626
rect 181536 151768 181588 151774
rect 181536 151710 181588 151716
rect 181548 3466 181576 151710
rect 181640 149938 181668 153598
rect 181824 152862 181852 160140
rect 181916 158114 181944 160140
rect 182008 158681 182036 160140
rect 181994 158672 182050 158681
rect 181994 158607 182050 158616
rect 181916 158086 182036 158114
rect 181902 157992 181958 158001
rect 181902 157927 181958 157936
rect 181916 157334 181944 157927
rect 182008 157826 182036 158086
rect 181996 157820 182048 157826
rect 181996 157762 182048 157768
rect 181916 157306 182036 157334
rect 181904 153196 181956 153202
rect 181904 153138 181956 153144
rect 181812 152856 181864 152862
rect 181812 152798 181864 152804
rect 181628 149932 181680 149938
rect 181628 149874 181680 149880
rect 181916 149054 181944 153138
rect 182008 153082 182036 157306
rect 182100 153202 182128 160140
rect 182088 153196 182140 153202
rect 182088 153138 182140 153144
rect 182008 153054 182128 153082
rect 181996 152380 182048 152386
rect 181996 152322 182048 152328
rect 181904 149048 181956 149054
rect 181904 148990 181956 148996
rect 182008 134570 182036 152322
rect 181996 134564 182048 134570
rect 181996 134506 182048 134512
rect 182100 129062 182128 153054
rect 182192 148850 182220 160140
rect 182284 158681 182312 160140
rect 182270 158672 182326 158681
rect 182270 158607 182326 158616
rect 182376 152930 182404 160140
rect 182468 158506 182496 160140
rect 182560 159905 182588 160140
rect 182546 159896 182602 159905
rect 182546 159831 182602 159840
rect 182548 159792 182600 159798
rect 182546 159760 182548 159769
rect 182600 159760 182602 159769
rect 182546 159695 182602 159704
rect 182456 158500 182508 158506
rect 182456 158442 182508 158448
rect 182548 156732 182600 156738
rect 182548 156674 182600 156680
rect 182364 152924 182416 152930
rect 182364 152866 182416 152872
rect 182456 152584 182508 152590
rect 182456 152526 182508 152532
rect 182272 152516 182324 152522
rect 182272 152458 182324 152464
rect 182180 148844 182232 148850
rect 182180 148786 182232 148792
rect 182180 148708 182232 148714
rect 182180 148650 182232 148656
rect 182088 129056 182140 129062
rect 182088 128998 182140 129004
rect 181536 3460 181588 3466
rect 181536 3402 181588 3408
rect 181444 3052 181496 3058
rect 181444 2994 181496 3000
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 148650
rect 182284 140758 182312 152458
rect 182364 152380 182416 152386
rect 182364 152322 182416 152328
rect 182376 143206 182404 152322
rect 182468 147422 182496 152526
rect 182560 148714 182588 156674
rect 182652 151706 182680 160140
rect 182744 158710 182772 160140
rect 182732 158704 182784 158710
rect 182732 158646 182784 158652
rect 182732 158568 182784 158574
rect 182732 158510 182784 158516
rect 182640 151700 182692 151706
rect 182640 151642 182692 151648
rect 182548 148708 182600 148714
rect 182548 148650 182600 148656
rect 182744 147674 182772 158510
rect 182836 152522 182864 160140
rect 182928 154222 182956 160140
rect 183020 159746 183048 160140
rect 183112 159866 183140 160140
rect 183100 159860 183152 159866
rect 183100 159802 183152 159808
rect 183020 159718 183140 159746
rect 183112 157146 183140 159718
rect 183100 157140 183152 157146
rect 183100 157082 183152 157088
rect 182916 154216 182968 154222
rect 182916 154158 182968 154164
rect 182916 152652 182968 152658
rect 182916 152594 182968 152600
rect 182824 152516 182876 152522
rect 182824 152458 182876 152464
rect 182744 147646 182864 147674
rect 182456 147416 182508 147422
rect 182456 147358 182508 147364
rect 182364 143200 182416 143206
rect 182364 143142 182416 143148
rect 182272 140752 182324 140758
rect 182272 140694 182324 140700
rect 182836 3398 182864 147646
rect 182928 3602 182956 152594
rect 183204 152590 183232 160140
rect 183296 157690 183324 160140
rect 183388 159905 183416 160140
rect 183374 159896 183430 159905
rect 183374 159831 183430 159840
rect 183284 157684 183336 157690
rect 183284 157626 183336 157632
rect 183284 152992 183336 152998
rect 183284 152934 183336 152940
rect 183296 152590 183324 152934
rect 183192 152584 183244 152590
rect 183192 152526 183244 152532
rect 183284 152584 183336 152590
rect 183284 152526 183336 152532
rect 183388 147674 183416 159831
rect 183480 152386 183508 160140
rect 183468 152380 183520 152386
rect 183468 152322 183520 152328
rect 183572 148986 183600 160140
rect 183664 157457 183692 160140
rect 183756 159526 183784 160140
rect 183744 159520 183796 159526
rect 183744 159462 183796 159468
rect 183650 157448 183706 157457
rect 183650 157383 183706 157392
rect 183848 154290 183876 160140
rect 183940 159905 183968 160140
rect 183926 159896 183982 159905
rect 183926 159831 183982 159840
rect 183836 154284 183888 154290
rect 183836 154226 183888 154232
rect 184032 149598 184060 160140
rect 184124 156330 184152 160140
rect 184216 159769 184244 160140
rect 184202 159760 184258 159769
rect 184202 159695 184258 159704
rect 184112 156324 184164 156330
rect 184112 156266 184164 156272
rect 184020 149592 184072 149598
rect 184020 149534 184072 149540
rect 183560 148980 183612 148986
rect 183560 148922 183612 148928
rect 184308 148782 184336 160140
rect 184400 157758 184428 160140
rect 184492 159905 184520 160140
rect 184478 159896 184534 159905
rect 184478 159831 184534 159840
rect 184388 157752 184440 157758
rect 184388 157694 184440 157700
rect 184480 157684 184532 157690
rect 184480 157626 184532 157632
rect 184296 148776 184348 148782
rect 184296 148718 184348 148724
rect 184492 148714 184520 157626
rect 184480 148708 184532 148714
rect 184480 148650 184532 148656
rect 184584 148594 184612 160140
rect 184676 154902 184704 160140
rect 184664 154896 184716 154902
rect 184664 154838 184716 154844
rect 183664 148566 184612 148594
rect 183388 147646 183508 147674
rect 183376 140752 183428 140758
rect 183376 140694 183428 140700
rect 183388 140554 183416 140694
rect 183376 140548 183428 140554
rect 183376 140490 183428 140496
rect 183388 111110 183416 140490
rect 183376 111104 183428 111110
rect 183376 111046 183428 111052
rect 183480 94586 183508 147646
rect 183664 146198 183692 148566
rect 184768 147354 184796 160140
rect 184756 147348 184808 147354
rect 184756 147290 184808 147296
rect 183652 146192 183704 146198
rect 183652 146134 183704 146140
rect 184860 139262 184888 160140
rect 184952 151298 184980 160140
rect 185044 157457 185072 160140
rect 185136 159118 185164 160140
rect 185124 159112 185176 159118
rect 185124 159054 185176 159060
rect 185228 157962 185256 160140
rect 185320 159905 185348 160140
rect 185306 159896 185362 159905
rect 185306 159831 185362 159840
rect 185216 157956 185268 157962
rect 185216 157898 185268 157904
rect 185030 157448 185086 157457
rect 185030 157383 185086 157392
rect 185412 156534 185440 160140
rect 185400 156528 185452 156534
rect 185400 156470 185452 156476
rect 185504 155854 185532 160140
rect 185492 155848 185544 155854
rect 185492 155790 185544 155796
rect 185492 152788 185544 152794
rect 185492 152730 185544 152736
rect 185504 152658 185532 152730
rect 185492 152652 185544 152658
rect 185492 152594 185544 152600
rect 185596 152538 185624 160140
rect 185124 152516 185176 152522
rect 185124 152458 185176 152464
rect 185228 152510 185624 152538
rect 185032 152244 185084 152250
rect 185032 152186 185084 152192
rect 184940 151292 184992 151298
rect 184940 151234 184992 151240
rect 185044 141846 185072 152186
rect 185136 144838 185164 152458
rect 185124 144832 185176 144838
rect 185124 144774 185176 144780
rect 185228 144430 185256 152510
rect 185308 152380 185360 152386
rect 185308 152322 185360 152328
rect 185320 147286 185348 152322
rect 185688 151570 185716 160140
rect 185780 157690 185808 160140
rect 185872 158778 185900 160140
rect 185860 158772 185912 158778
rect 185860 158714 185912 158720
rect 185860 157888 185912 157894
rect 185860 157830 185912 157836
rect 185768 157684 185820 157690
rect 185768 157626 185820 157632
rect 185768 156596 185820 156602
rect 185768 156538 185820 156544
rect 185676 151564 185728 151570
rect 185676 151506 185728 151512
rect 185308 147280 185360 147286
rect 185308 147222 185360 147228
rect 185216 144424 185268 144430
rect 185216 144366 185268 144372
rect 185032 141840 185084 141846
rect 185032 141782 185084 141788
rect 184848 139256 184900 139262
rect 184848 139198 184900 139204
rect 183468 94580 183520 94586
rect 183468 94522 183520 94528
rect 185780 16574 185808 156538
rect 185872 154970 185900 157830
rect 185860 154964 185912 154970
rect 185860 154906 185912 154912
rect 185964 152522 185992 160140
rect 186056 157894 186084 160140
rect 186044 157888 186096 157894
rect 186044 157830 186096 157836
rect 186044 157752 186096 157758
rect 186044 157694 186096 157700
rect 185952 152516 186004 152522
rect 185952 152458 186004 152464
rect 186056 148918 186084 157694
rect 186148 152386 186176 160140
rect 186136 152380 186188 152386
rect 186136 152322 186188 152328
rect 186240 152250 186268 160140
rect 186332 158681 186360 160140
rect 186318 158672 186374 158681
rect 186318 158607 186374 158616
rect 186320 158160 186372 158166
rect 186320 158102 186372 158108
rect 186332 157894 186360 158102
rect 186320 157888 186372 157894
rect 186320 157830 186372 157836
rect 186424 157334 186452 160140
rect 186332 157306 186452 157334
rect 186228 152244 186280 152250
rect 186228 152186 186280 152192
rect 186044 148912 186096 148918
rect 186044 148854 186096 148860
rect 186332 139641 186360 157306
rect 186516 153134 186544 160140
rect 186608 157334 186636 160140
rect 186700 158545 186728 160140
rect 186686 158536 186742 158545
rect 186686 158471 186742 158480
rect 186608 157306 186728 157334
rect 186504 153128 186556 153134
rect 186504 153070 186556 153076
rect 186596 152584 186648 152590
rect 186596 152526 186648 152532
rect 186504 152380 186556 152386
rect 186504 152322 186556 152328
rect 186412 152244 186464 152250
rect 186412 152186 186464 152192
rect 186318 139632 186374 139641
rect 186318 139567 186374 139576
rect 186318 138680 186374 138689
rect 186318 138615 186374 138624
rect 186332 16574 186360 138615
rect 186424 132394 186452 152186
rect 186516 139398 186544 152322
rect 186608 140758 186636 152526
rect 186700 150414 186728 157306
rect 186792 154574 186820 160140
rect 186884 158574 186912 160140
rect 186872 158568 186924 158574
rect 186872 158510 186924 158516
rect 186792 154546 186912 154574
rect 186688 150408 186740 150414
rect 186688 150350 186740 150356
rect 186688 149728 186740 149734
rect 186688 149670 186740 149676
rect 186596 140752 186648 140758
rect 186596 140694 186648 140700
rect 186700 139505 186728 149670
rect 186884 144914 186912 154546
rect 186976 149734 187004 160140
rect 187068 152590 187096 160140
rect 187160 158642 187188 160140
rect 187252 158681 187280 160140
rect 187238 158672 187294 158681
rect 187148 158636 187200 158642
rect 187238 158607 187294 158616
rect 187148 158578 187200 158584
rect 187148 157684 187200 157690
rect 187148 157626 187200 157632
rect 187160 152794 187188 157626
rect 187148 152788 187200 152794
rect 187148 152730 187200 152736
rect 187056 152584 187108 152590
rect 187056 152526 187108 152532
rect 187344 152386 187372 160140
rect 187436 159497 187464 160140
rect 187422 159488 187478 159497
rect 187422 159423 187478 159432
rect 187424 158704 187476 158710
rect 187528 158681 187556 160140
rect 187424 158646 187476 158652
rect 187514 158672 187570 158681
rect 187332 152380 187384 152386
rect 187332 152322 187384 152328
rect 187436 150210 187464 158646
rect 187514 158607 187570 158616
rect 187620 152250 187648 160140
rect 187712 159390 187740 160140
rect 187700 159384 187752 159390
rect 187700 159326 187752 159332
rect 187804 158681 187832 160140
rect 187790 158672 187846 158681
rect 187790 158607 187846 158616
rect 187896 157334 187924 160140
rect 187988 157350 188016 160140
rect 187804 157306 187924 157334
rect 187976 157344 188028 157350
rect 187700 152584 187752 152590
rect 187700 152526 187752 152532
rect 187608 152244 187660 152250
rect 187608 152186 187660 152192
rect 187424 150204 187476 150210
rect 187424 150146 187476 150152
rect 186964 149728 187016 149734
rect 186964 149670 187016 149676
rect 186792 144886 186912 144914
rect 186792 143478 186820 144886
rect 186780 143472 186832 143478
rect 186780 143414 186832 143420
rect 187514 140312 187570 140321
rect 187514 140247 187570 140256
rect 187528 139641 187556 140247
rect 187606 140176 187662 140185
rect 187606 140111 187662 140120
rect 187514 139632 187570 139641
rect 187514 139567 187570 139576
rect 186686 139496 186742 139505
rect 186686 139431 186742 139440
rect 186504 139392 186556 139398
rect 186504 139334 186556 139340
rect 186412 132388 186464 132394
rect 186412 132330 186464 132336
rect 187528 116686 187556 139567
rect 187620 139505 187648 140111
rect 187606 139496 187662 139505
rect 187606 139431 187662 139440
rect 187516 116680 187568 116686
rect 187516 116622 187568 116628
rect 187620 22778 187648 139431
rect 187712 137970 187740 152526
rect 187804 150278 187832 157306
rect 187976 157286 188028 157292
rect 188080 152674 188108 160140
rect 187896 152646 188108 152674
rect 187792 150272 187844 150278
rect 187792 150214 187844 150220
rect 187792 149320 187844 149326
rect 187792 149262 187844 149268
rect 187804 141506 187832 149262
rect 187792 141500 187844 141506
rect 187792 141442 187844 141448
rect 187896 141438 187924 152646
rect 188172 152538 188200 160140
rect 187988 152510 188200 152538
rect 187988 146742 188016 152510
rect 188264 147674 188292 160140
rect 188356 159905 188384 160140
rect 188342 159896 188398 159905
rect 188342 159831 188398 159840
rect 188448 158760 188476 160140
rect 188356 158732 188476 158760
rect 188356 152386 188384 158732
rect 188540 158658 188568 160140
rect 188632 158681 188660 160140
rect 188448 158630 188568 158658
rect 188618 158672 188674 158681
rect 188448 154426 188476 158630
rect 188618 158607 188674 158616
rect 188528 158568 188580 158574
rect 188528 158510 188580 158516
rect 188436 154420 188488 154426
rect 188436 154362 188488 154368
rect 188344 152380 188396 152386
rect 188344 152322 188396 152328
rect 188540 149666 188568 158510
rect 188724 152590 188752 160140
rect 188816 158302 188844 160140
rect 188908 158681 188936 160140
rect 189000 159866 189028 160140
rect 188988 159860 189040 159866
rect 188988 159802 189040 159808
rect 188894 158672 188950 158681
rect 188894 158607 188950 158616
rect 188804 158296 188856 158302
rect 188804 158238 188856 158244
rect 188712 152584 188764 152590
rect 188712 152526 188764 152532
rect 188896 152380 188948 152386
rect 188896 152322 188948 152328
rect 188908 152182 188936 152322
rect 188896 152176 188948 152182
rect 188896 152118 188948 152124
rect 188528 149660 188580 149666
rect 188528 149602 188580 149608
rect 188080 147646 188292 147674
rect 188080 147150 188108 147646
rect 188068 147144 188120 147150
rect 188068 147086 188120 147092
rect 187976 146736 188028 146742
rect 187976 146678 188028 146684
rect 187884 141432 187936 141438
rect 187884 141374 187936 141380
rect 187700 137964 187752 137970
rect 187700 137906 187752 137912
rect 188908 72486 188936 152118
rect 189000 149326 189028 159802
rect 189092 151230 189120 160140
rect 189184 158681 189212 160140
rect 189170 158672 189226 158681
rect 189170 158607 189226 158616
rect 189172 158228 189224 158234
rect 189172 158170 189224 158176
rect 189184 158030 189212 158170
rect 189172 158024 189224 158030
rect 189172 157966 189224 157972
rect 189276 152998 189304 160140
rect 189368 158234 189396 160140
rect 189356 158228 189408 158234
rect 189356 158170 189408 158176
rect 189460 157334 189488 160140
rect 189368 157306 189488 157334
rect 189264 152992 189316 152998
rect 189264 152934 189316 152940
rect 189172 152584 189224 152590
rect 189368 152538 189396 157306
rect 189172 152526 189224 152532
rect 189080 151224 189132 151230
rect 189080 151166 189132 151172
rect 189080 151088 189132 151094
rect 189080 151030 189132 151036
rect 188988 149320 189040 149326
rect 188988 149262 189040 149268
rect 188988 141704 189040 141710
rect 188988 141646 189040 141652
rect 189000 141438 189028 141646
rect 188988 141432 189040 141438
rect 188988 141374 189040 141380
rect 188896 72480 188948 72486
rect 188896 72422 188948 72428
rect 187700 66904 187752 66910
rect 187700 66846 187752 66852
rect 187608 22772 187660 22778
rect 187608 22714 187660 22720
rect 187712 16574 187740 66846
rect 185780 16546 186176 16574
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 184940 3800 184992 3806
rect 184940 3742 184992 3748
rect 182916 3596 182968 3602
rect 182916 3538 182968 3544
rect 183744 3460 183796 3466
rect 183744 3402 183796 3408
rect 182824 3392 182876 3398
rect 182824 3334 182876 3340
rect 183756 480 183784 3402
rect 184952 480 184980 3742
rect 186148 480 186176 16546
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189000 4826 189028 141374
rect 189092 128314 189120 151030
rect 189184 136474 189212 152526
rect 189276 152510 189396 152538
rect 189276 141642 189304 152510
rect 189552 151722 189580 160140
rect 189644 151774 189672 160140
rect 189736 159905 189764 160140
rect 189722 159896 189778 159905
rect 189722 159831 189778 159840
rect 189724 158500 189776 158506
rect 189724 158442 189776 158448
rect 189368 151694 189580 151722
rect 189632 151768 189684 151774
rect 189632 151710 189684 151716
rect 189368 144770 189396 151694
rect 189540 151224 189592 151230
rect 189540 151166 189592 151172
rect 189448 151156 189500 151162
rect 189448 151098 189500 151104
rect 189460 146130 189488 151098
rect 189552 146946 189580 151166
rect 189736 148510 189764 158442
rect 189828 152590 189856 160140
rect 189920 155990 189948 160140
rect 190012 158681 190040 160140
rect 189998 158672 190054 158681
rect 189998 158607 190054 158616
rect 190104 157334 190132 160140
rect 190012 157306 190132 157334
rect 189908 155984 189960 155990
rect 189908 155926 189960 155932
rect 189816 152584 189868 152590
rect 189816 152526 189868 152532
rect 190012 151162 190040 157306
rect 190196 157214 190224 160140
rect 190288 158681 190316 160140
rect 190274 158672 190330 158681
rect 190274 158607 190330 158616
rect 190184 157208 190236 157214
rect 190184 157150 190236 157156
rect 190276 155780 190328 155786
rect 190276 155722 190328 155728
rect 190288 154902 190316 155722
rect 190276 154896 190328 154902
rect 190276 154838 190328 154844
rect 190184 152992 190236 152998
rect 190184 152934 190236 152940
rect 190092 151768 190144 151774
rect 190092 151710 190144 151716
rect 190000 151156 190052 151162
rect 190000 151098 190052 151104
rect 190104 150890 190132 151710
rect 190092 150884 190144 150890
rect 190092 150826 190144 150832
rect 189724 148504 189776 148510
rect 189724 148446 189776 148452
rect 190196 148170 190224 152934
rect 190380 151094 190408 160140
rect 190472 158710 190500 160140
rect 190460 158704 190512 158710
rect 190460 158646 190512 158652
rect 190460 157684 190512 157690
rect 190460 157626 190512 157632
rect 190368 151088 190420 151094
rect 190368 151030 190420 151036
rect 190184 148164 190236 148170
rect 190184 148106 190236 148112
rect 189540 146940 189592 146946
rect 189540 146882 189592 146888
rect 189448 146124 189500 146130
rect 189448 146066 189500 146072
rect 189356 144764 189408 144770
rect 189356 144706 189408 144712
rect 189264 141636 189316 141642
rect 189264 141578 189316 141584
rect 190368 141636 190420 141642
rect 190368 141578 190420 141584
rect 189998 140448 190054 140457
rect 189998 140383 190000 140392
rect 190052 140383 190054 140392
rect 190000 140354 190052 140360
rect 189172 136468 189224 136474
rect 189172 136410 189224 136416
rect 189080 128308 189132 128314
rect 189080 128250 189132 128256
rect 190380 104174 190408 141578
rect 190472 125594 190500 157626
rect 190564 152998 190592 160140
rect 190656 158681 190684 160140
rect 190642 158672 190698 158681
rect 190642 158607 190698 158616
rect 190748 157282 190776 160140
rect 190840 158409 190868 160140
rect 190932 158982 190960 160140
rect 191024 159594 191052 160140
rect 191116 159905 191144 160140
rect 191102 159896 191158 159905
rect 191102 159831 191158 159840
rect 191104 159792 191156 159798
rect 191104 159734 191156 159740
rect 191012 159588 191064 159594
rect 191012 159530 191064 159536
rect 190920 158976 190972 158982
rect 190920 158918 190972 158924
rect 190920 158704 190972 158710
rect 190920 158646 190972 158652
rect 191012 158704 191064 158710
rect 191012 158646 191064 158652
rect 190826 158400 190882 158409
rect 190826 158335 190882 158344
rect 190736 157276 190788 157282
rect 190736 157218 190788 157224
rect 190932 154902 190960 158646
rect 191024 156058 191052 158646
rect 191116 157690 191144 159734
rect 191104 157684 191156 157690
rect 191104 157626 191156 157632
rect 191208 157334 191236 160140
rect 191116 157306 191236 157334
rect 191012 156052 191064 156058
rect 191012 155994 191064 156000
rect 191012 155848 191064 155854
rect 191012 155790 191064 155796
rect 191024 155378 191052 155790
rect 191012 155372 191064 155378
rect 191012 155314 191064 155320
rect 191012 155236 191064 155242
rect 191012 155178 191064 155184
rect 190920 154896 190972 154902
rect 190920 154838 190972 154844
rect 191024 154766 191052 155178
rect 191012 154760 191064 154766
rect 191012 154702 191064 154708
rect 190552 152992 190604 152998
rect 190552 152934 190604 152940
rect 190552 152584 190604 152590
rect 191116 152538 191144 157306
rect 191196 156052 191248 156058
rect 191196 155994 191248 156000
rect 191208 153610 191236 155994
rect 191196 153604 191248 153610
rect 191196 153546 191248 153552
rect 190552 152526 190604 152532
rect 190564 135182 190592 152526
rect 190656 152510 191144 152538
rect 190656 146062 190684 152510
rect 191300 152402 191328 160140
rect 191392 158545 191420 160140
rect 191378 158536 191434 158545
rect 191378 158471 191434 158480
rect 191380 156732 191432 156738
rect 191380 156674 191432 156680
rect 191392 156602 191420 156674
rect 191380 156596 191432 156602
rect 191380 156538 191432 156544
rect 191380 155984 191432 155990
rect 191380 155926 191432 155932
rect 190748 152374 191328 152402
rect 190748 147218 190776 152374
rect 191392 147674 191420 155926
rect 191484 152590 191512 160140
rect 191576 158710 191604 160140
rect 191564 158704 191616 158710
rect 191564 158646 191616 158652
rect 191668 157321 191696 160140
rect 191760 159934 191788 160140
rect 191748 159928 191800 159934
rect 191748 159870 191800 159876
rect 191746 159760 191802 159769
rect 191746 159695 191802 159704
rect 191654 157312 191710 157321
rect 191654 157247 191710 157256
rect 191656 157208 191708 157214
rect 191656 157150 191708 157156
rect 191564 152992 191616 152998
rect 191564 152934 191616 152940
rect 191472 152584 191524 152590
rect 191472 152526 191524 152532
rect 191576 148306 191604 152934
rect 191668 148578 191696 157150
rect 191656 148572 191708 148578
rect 191656 148514 191708 148520
rect 191564 148300 191616 148306
rect 191564 148242 191616 148248
rect 191116 147646 191420 147674
rect 190736 147212 190788 147218
rect 190736 147154 190788 147160
rect 191116 147014 191144 147646
rect 191104 147008 191156 147014
rect 191104 146950 191156 146956
rect 190644 146056 190696 146062
rect 190644 145998 190696 146004
rect 191654 140856 191710 140865
rect 191654 140791 191710 140800
rect 191668 140486 191696 140791
rect 191656 140480 191708 140486
rect 191656 140422 191708 140428
rect 190552 135176 190604 135182
rect 190552 135118 190604 135124
rect 190460 125588 190512 125594
rect 190460 125530 190512 125536
rect 189724 104168 189776 104174
rect 189724 104110 189776 104116
rect 190368 104168 190420 104174
rect 190368 104110 190420 104116
rect 189736 16574 189764 104110
rect 191104 60036 191156 60042
rect 191104 59978 191156 59984
rect 189736 16546 189856 16574
rect 188988 4820 189040 4826
rect 188988 4762 189040 4768
rect 189828 3738 189856 16546
rect 189816 3732 189868 3738
rect 189816 3674 189868 3680
rect 190828 3664 190880 3670
rect 190828 3606 190880 3612
rect 189724 3052 189776 3058
rect 189724 2994 189776 3000
rect 189736 480 189764 2994
rect 190840 480 190868 3606
rect 191116 3534 191144 59978
rect 191668 6254 191696 140422
rect 191760 6322 191788 159695
rect 191852 157334 191880 160140
rect 191944 158273 191972 160140
rect 192036 158642 192064 160140
rect 192024 158636 192076 158642
rect 192024 158578 192076 158584
rect 192022 158536 192078 158545
rect 192022 158471 192078 158480
rect 191930 158264 191986 158273
rect 191930 158199 191986 158208
rect 192036 158001 192064 158471
rect 192022 157992 192078 158001
rect 192022 157927 192078 157936
rect 192128 157826 192156 160140
rect 192220 159905 192248 160140
rect 192206 159896 192262 159905
rect 192206 159831 192262 159840
rect 192220 158137 192248 159831
rect 192206 158128 192262 158137
rect 192206 158063 192262 158072
rect 192116 157820 192168 157826
rect 192116 157762 192168 157768
rect 192208 157752 192260 157758
rect 192208 157694 192260 157700
rect 191852 157306 192156 157334
rect 191932 152584 191984 152590
rect 191932 152526 191984 152532
rect 191840 152244 191892 152250
rect 191840 152186 191892 152192
rect 191852 123554 191880 152186
rect 191944 132462 191972 152526
rect 192024 152380 192076 152386
rect 192024 152322 192076 152328
rect 192036 133890 192064 152322
rect 192128 151201 192156 157306
rect 192220 151230 192248 157694
rect 192208 151224 192260 151230
rect 192114 151192 192170 151201
rect 192208 151166 192260 151172
rect 192114 151127 192170 151136
rect 192312 147674 192340 160140
rect 192404 158817 192432 160140
rect 192390 158808 192446 158817
rect 192390 158743 192446 158752
rect 192392 158704 192444 158710
rect 192392 158646 192444 158652
rect 192404 157214 192432 158646
rect 192496 158545 192524 160140
rect 192482 158536 192538 158545
rect 192482 158471 192538 158480
rect 192392 157208 192444 157214
rect 192392 157150 192444 157156
rect 192588 152590 192616 160140
rect 192680 158710 192708 160140
rect 192668 158704 192720 158710
rect 192772 158681 192800 160140
rect 192668 158646 192720 158652
rect 192758 158672 192814 158681
rect 192758 158607 192814 158616
rect 192668 158296 192720 158302
rect 192668 158238 192720 158244
rect 192576 152584 192628 152590
rect 192576 152526 192628 152532
rect 192680 148374 192708 158238
rect 192864 152386 192892 160140
rect 192956 158914 192984 160140
rect 193048 159089 193076 160140
rect 193140 159934 193168 160140
rect 193128 159928 193180 159934
rect 193128 159870 193180 159876
rect 193034 159080 193090 159089
rect 193034 159015 193090 159024
rect 193140 158930 193168 159870
rect 192944 158908 192996 158914
rect 192944 158850 192996 158856
rect 193048 158902 193168 158930
rect 193048 158714 193076 158902
rect 193128 158840 193180 158846
rect 193128 158782 193180 158788
rect 192956 158686 193076 158714
rect 192852 152380 192904 152386
rect 192852 152322 192904 152328
rect 192956 152250 192984 158686
rect 193140 158658 193168 158782
rect 193048 158630 193168 158658
rect 193048 155174 193076 158630
rect 193232 158273 193260 160140
rect 193324 158914 193352 160140
rect 193312 158908 193364 158914
rect 193312 158850 193364 158856
rect 193218 158264 193274 158273
rect 193218 158199 193274 158208
rect 193126 158128 193182 158137
rect 193126 158063 193182 158072
rect 193036 155168 193088 155174
rect 193036 155110 193088 155116
rect 193036 152788 193088 152794
rect 193036 152730 193088 152736
rect 193048 152386 193076 152730
rect 193036 152380 193088 152386
rect 193036 152322 193088 152328
rect 192944 152244 192996 152250
rect 192944 152186 192996 152192
rect 192668 148368 192720 148374
rect 192668 148310 192720 148316
rect 192128 147646 192340 147674
rect 192128 139330 192156 147646
rect 192116 139324 192168 139330
rect 192116 139266 192168 139272
rect 192024 133884 192076 133890
rect 192024 133826 192076 133832
rect 191932 132456 191984 132462
rect 191932 132398 191984 132404
rect 191840 123548 191892 123554
rect 191840 123490 191892 123496
rect 193140 9042 193168 158063
rect 193312 152788 193364 152794
rect 193312 152730 193364 152736
rect 193220 152584 193272 152590
rect 193220 152526 193272 152532
rect 193232 142118 193260 152526
rect 193324 143546 193352 152730
rect 193416 151745 193444 160140
rect 193508 156641 193536 160140
rect 193600 159905 193628 160140
rect 193586 159896 193642 159905
rect 193586 159831 193642 159840
rect 193692 158760 193720 160140
rect 193600 158732 193720 158760
rect 193494 156632 193550 156641
rect 193494 156567 193550 156576
rect 193600 155922 193628 158732
rect 193680 158636 193732 158642
rect 193680 158578 193732 158584
rect 193588 155916 193640 155922
rect 193588 155858 193640 155864
rect 193588 155304 193640 155310
rect 193588 155246 193640 155252
rect 193402 151736 193458 151745
rect 193402 151671 193458 151680
rect 193600 147674 193628 155246
rect 193692 152538 193720 158578
rect 193784 158574 193812 160140
rect 193876 159905 193904 160140
rect 193862 159896 193918 159905
rect 193862 159831 193918 159840
rect 193772 158568 193824 158574
rect 193772 158510 193824 158516
rect 193876 152674 193904 159831
rect 193968 152794 193996 160140
rect 194060 158302 194088 160140
rect 194152 158681 194180 160140
rect 194138 158672 194194 158681
rect 194138 158607 194194 158616
rect 194048 158296 194100 158302
rect 194048 158238 194100 158244
rect 194140 157820 194192 157826
rect 194140 157762 194192 157768
rect 193956 152788 194008 152794
rect 193956 152730 194008 152736
rect 193876 152646 194088 152674
rect 193692 152510 193996 152538
rect 193600 147646 193904 147674
rect 193312 143540 193364 143546
rect 193312 143482 193364 143488
rect 193220 142112 193272 142118
rect 193220 142054 193272 142060
rect 193128 9036 193180 9042
rect 193128 8978 193180 8984
rect 191748 6316 191800 6322
rect 191748 6258 191800 6264
rect 191656 6248 191708 6254
rect 191656 6190 191708 6196
rect 193876 4078 193904 147646
rect 193968 143342 193996 152510
rect 194060 147674 194088 152646
rect 194152 148646 194180 157762
rect 194244 152590 194272 160140
rect 194336 158522 194364 160140
rect 194428 158681 194456 160140
rect 194414 158672 194470 158681
rect 194414 158607 194470 158616
rect 194520 158545 194548 160140
rect 194612 158710 194640 160140
rect 194600 158704 194652 158710
rect 194600 158646 194652 158652
rect 194506 158536 194562 158545
rect 194336 158494 194456 158522
rect 194322 158400 194378 158409
rect 194322 158335 194378 158344
rect 194232 152584 194284 152590
rect 194232 152526 194284 152532
rect 194336 152538 194364 158335
rect 194428 157758 194456 158494
rect 194506 158471 194562 158480
rect 194704 158409 194732 160140
rect 194690 158400 194746 158409
rect 194690 158335 194746 158344
rect 194508 158296 194560 158302
rect 194508 158238 194560 158244
rect 194416 157752 194468 157758
rect 194416 157694 194468 157700
rect 194520 157334 194548 158238
rect 194520 157306 194640 157334
rect 194612 157026 194640 157306
rect 194520 156998 194640 157026
rect 194520 154630 194548 156998
rect 194508 154624 194560 154630
rect 194508 154566 194560 154572
rect 194692 152584 194744 152590
rect 194336 152510 194548 152538
rect 194692 152526 194744 152532
rect 194140 148640 194192 148646
rect 194140 148582 194192 148588
rect 194060 147646 194456 147674
rect 193956 143336 194008 143342
rect 193956 143278 194008 143284
rect 194428 112470 194456 147646
rect 194416 112464 194468 112470
rect 194416 112406 194468 112412
rect 194520 79354 194548 152510
rect 194704 142050 194732 152526
rect 194796 147490 194824 160140
rect 194888 158642 194916 160140
rect 194980 159769 195008 160140
rect 194966 159760 195022 159769
rect 194966 159695 195022 159704
rect 194876 158636 194928 158642
rect 194876 158578 194928 158584
rect 194876 157956 194928 157962
rect 194876 157898 194928 157904
rect 194888 152794 194916 157898
rect 194876 152788 194928 152794
rect 194876 152730 194928 152736
rect 194980 152250 195008 159695
rect 195072 152590 195100 160140
rect 195164 157826 195192 160140
rect 195256 159905 195284 160140
rect 195242 159896 195298 159905
rect 195242 159831 195298 159840
rect 195244 158568 195296 158574
rect 195244 158510 195296 158516
rect 195152 157820 195204 157826
rect 195152 157762 195204 157768
rect 195060 152584 195112 152590
rect 195060 152526 195112 152532
rect 195152 152584 195204 152590
rect 195152 152526 195204 152532
rect 194968 152244 195020 152250
rect 194968 152186 195020 152192
rect 195164 152182 195192 152526
rect 195152 152176 195204 152182
rect 195152 152118 195204 152124
rect 195256 147674 195284 158510
rect 195348 155700 195376 160140
rect 195440 157690 195468 160140
rect 195532 159905 195560 160140
rect 195518 159896 195574 159905
rect 195518 159831 195574 159840
rect 195624 158930 195652 160140
rect 195532 158902 195652 158930
rect 195532 158681 195560 158902
rect 195716 158760 195744 160140
rect 195808 159905 195836 160140
rect 195794 159896 195850 159905
rect 195794 159831 195850 159840
rect 195624 158732 195744 158760
rect 195518 158672 195574 158681
rect 195518 158607 195574 158616
rect 195520 157888 195572 157894
rect 195520 157830 195572 157836
rect 195428 157684 195480 157690
rect 195428 157626 195480 157632
rect 195348 155672 195468 155700
rect 195440 147674 195468 155672
rect 195532 151026 195560 157830
rect 195624 153270 195652 158732
rect 195704 158636 195756 158642
rect 195704 158578 195756 158584
rect 195716 155145 195744 158578
rect 195702 155136 195758 155145
rect 195702 155071 195758 155080
rect 195612 153264 195664 153270
rect 195612 153206 195664 153212
rect 195520 151020 195572 151026
rect 195520 150962 195572 150968
rect 195256 147646 195376 147674
rect 195440 147646 195652 147674
rect 194784 147484 194836 147490
rect 194784 147426 194836 147432
rect 195348 145994 195376 147646
rect 195336 145988 195388 145994
rect 195336 145930 195388 145936
rect 194692 142044 194744 142050
rect 194692 141986 194744 141992
rect 195426 140312 195482 140321
rect 195426 140247 195482 140256
rect 195440 139777 195468 140247
rect 195426 139768 195482 139777
rect 195426 139703 195482 139712
rect 195624 129674 195652 147646
rect 195612 129668 195664 129674
rect 195612 129610 195664 129616
rect 194508 79348 194560 79354
rect 194508 79290 194560 79296
rect 195808 15910 195836 159831
rect 195900 158545 195928 160140
rect 195886 158536 195942 158545
rect 195886 158471 195942 158480
rect 195992 157334 196020 160140
rect 196084 158681 196112 160140
rect 196070 158672 196126 158681
rect 196070 158607 196126 158616
rect 196176 157962 196204 160140
rect 196164 157956 196216 157962
rect 196164 157898 196216 157904
rect 195992 157306 196112 157334
rect 195888 155916 195940 155922
rect 195888 155858 195940 155864
rect 195900 155666 195928 155858
rect 195900 155638 196020 155666
rect 195888 152244 195940 152250
rect 195888 152186 195940 152192
rect 195152 15904 195204 15910
rect 195152 15846 195204 15852
rect 195796 15904 195848 15910
rect 195796 15846 195848 15852
rect 193864 4072 193916 4078
rect 193864 4014 193916 4020
rect 194416 3732 194468 3738
rect 194416 3674 194468 3680
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 191104 3528 191156 3534
rect 191104 3470 191156 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 192036 480 192064 3470
rect 193232 480 193260 3538
rect 194428 480 194456 3674
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 15846
rect 195900 8974 195928 152186
rect 195992 128246 196020 155638
rect 196084 152998 196112 157306
rect 196268 156942 196296 160140
rect 196360 159769 196388 160140
rect 196346 159760 196402 159769
rect 196346 159695 196402 159704
rect 196256 156936 196308 156942
rect 196256 156878 196308 156884
rect 196072 152992 196124 152998
rect 196072 152934 196124 152940
rect 196452 152266 196480 160140
rect 196544 154494 196572 160140
rect 196636 159905 196664 160140
rect 196622 159896 196678 159905
rect 196622 159831 196678 159840
rect 196622 157992 196678 158001
rect 196622 157927 196678 157936
rect 196532 154488 196584 154494
rect 196532 154430 196584 154436
rect 196532 152992 196584 152998
rect 196532 152934 196584 152940
rect 196072 152244 196124 152250
rect 196072 152186 196124 152192
rect 196176 152238 196480 152266
rect 196084 136542 196112 152186
rect 196176 144906 196204 152238
rect 196256 152176 196308 152182
rect 196256 152118 196308 152124
rect 196164 144900 196216 144906
rect 196164 144842 196216 144848
rect 196268 144498 196296 152118
rect 196544 147674 196572 152934
rect 196636 150006 196664 157927
rect 196728 152250 196756 160140
rect 196820 158137 196848 160140
rect 196806 158128 196862 158137
rect 196806 158063 196862 158072
rect 196808 157752 196860 157758
rect 196808 157694 196860 157700
rect 196716 152244 196768 152250
rect 196716 152186 196768 152192
rect 196624 150000 196676 150006
rect 196624 149942 196676 149948
rect 196820 147674 196848 157694
rect 196912 152182 196940 160140
rect 197004 155854 197032 160140
rect 197096 159225 197124 160140
rect 197082 159216 197138 159225
rect 197082 159151 197138 159160
rect 197084 158024 197136 158030
rect 197084 157966 197136 157972
rect 196992 155848 197044 155854
rect 196992 155790 197044 155796
rect 196900 152176 196952 152182
rect 196900 152118 196952 152124
rect 197096 151094 197124 157966
rect 197188 151473 197216 160140
rect 197280 158681 197308 160140
rect 197266 158672 197322 158681
rect 197266 158607 197322 158616
rect 197372 158574 197400 160140
rect 197360 158568 197412 158574
rect 197360 158510 197412 158516
rect 197266 153232 197322 153241
rect 197266 153167 197322 153176
rect 197174 151464 197230 151473
rect 197174 151399 197230 151408
rect 197084 151088 197136 151094
rect 197084 151030 197136 151036
rect 196360 147646 196572 147674
rect 196728 147646 196848 147674
rect 196360 147082 196388 147646
rect 196348 147076 196400 147082
rect 196348 147018 196400 147024
rect 196728 145926 196756 147646
rect 196716 145920 196768 145926
rect 196716 145862 196768 145868
rect 196256 144492 196308 144498
rect 196256 144434 196308 144440
rect 196072 136536 196124 136542
rect 196072 136478 196124 136484
rect 195980 128240 196032 128246
rect 195980 128182 196032 128188
rect 196622 120864 196678 120873
rect 196622 120799 196678 120808
rect 195888 8968 195940 8974
rect 195888 8910 195940 8916
rect 196636 3058 196664 120799
rect 197280 6186 197308 153167
rect 197464 152538 197492 160140
rect 197556 154601 197584 160140
rect 197542 154592 197598 154601
rect 197542 154527 197598 154536
rect 197464 152510 197584 152538
rect 197360 152244 197412 152250
rect 197360 152186 197412 152192
rect 197372 140690 197400 152186
rect 197452 152176 197504 152182
rect 197452 152118 197504 152124
rect 197360 140684 197412 140690
rect 197360 140626 197412 140632
rect 197464 13122 197492 152118
rect 197556 143410 197584 152510
rect 197648 150074 197676 160140
rect 197740 159769 197768 160140
rect 197726 159760 197782 159769
rect 197726 159695 197782 159704
rect 197728 157820 197780 157826
rect 197728 157762 197780 157768
rect 197636 150068 197688 150074
rect 197636 150010 197688 150016
rect 197740 145858 197768 157762
rect 197832 147674 197860 160140
rect 197924 158234 197952 160140
rect 198016 159905 198044 160140
rect 198002 159896 198058 159905
rect 198002 159831 198058 159840
rect 197912 158228 197964 158234
rect 197912 158170 197964 158176
rect 198004 158092 198056 158098
rect 198004 158034 198056 158040
rect 198016 151162 198044 158034
rect 198108 152250 198136 160140
rect 198200 159633 198228 160140
rect 198186 159624 198242 159633
rect 198186 159559 198242 159568
rect 198292 158681 198320 160140
rect 198278 158672 198334 158681
rect 198278 158607 198334 158616
rect 198280 158160 198332 158166
rect 198280 158102 198332 158108
rect 198188 157956 198240 157962
rect 198188 157898 198240 157904
rect 198200 157321 198228 157898
rect 198292 157554 198320 158102
rect 198280 157548 198332 157554
rect 198280 157490 198332 157496
rect 198186 157312 198242 157321
rect 198186 157247 198242 157256
rect 198384 153921 198412 160140
rect 198476 159633 198504 160140
rect 198568 159905 198596 160140
rect 198554 159896 198610 159905
rect 198554 159831 198610 159840
rect 198462 159624 198518 159633
rect 198462 159559 198518 159568
rect 198370 153912 198426 153921
rect 198370 153847 198426 153856
rect 198096 152244 198148 152250
rect 198096 152186 198148 152192
rect 198384 151994 198412 153847
rect 198568 152182 198596 159831
rect 198660 158681 198688 160140
rect 198752 158930 198780 160140
rect 198844 159905 198872 160140
rect 198830 159896 198886 159905
rect 198830 159831 198886 159840
rect 198936 158953 198964 160140
rect 199028 159798 199056 160140
rect 199120 159905 199148 160140
rect 199106 159896 199162 159905
rect 199106 159831 199162 159840
rect 199016 159792 199068 159798
rect 199016 159734 199068 159740
rect 198922 158944 198978 158953
rect 198752 158902 198872 158930
rect 198844 158794 198872 158902
rect 198922 158879 198978 158888
rect 198844 158766 199056 158794
rect 198646 158672 198702 158681
rect 198646 158607 198702 158616
rect 198924 158636 198976 158642
rect 198924 158578 198976 158584
rect 198738 158400 198794 158409
rect 198738 158335 198794 158344
rect 198556 152176 198608 152182
rect 198556 152118 198608 152124
rect 198384 151966 198596 151994
rect 198004 151156 198056 151162
rect 198004 151098 198056 151104
rect 197832 147646 198504 147674
rect 197728 145852 197780 145858
rect 197728 145794 197780 145800
rect 197544 143404 197596 143410
rect 197544 143346 197596 143352
rect 198476 141982 198504 147646
rect 198464 141976 198516 141982
rect 198464 141918 198516 141924
rect 198568 116618 198596 151966
rect 198648 140616 198700 140622
rect 198648 140558 198700 140564
rect 198660 139777 198688 140558
rect 198646 139768 198702 139777
rect 198646 139703 198702 139712
rect 198556 116612 198608 116618
rect 198556 116554 198608 116560
rect 198002 24168 198058 24177
rect 198002 24103 198058 24112
rect 197452 13116 197504 13122
rect 197452 13058 197504 13064
rect 197268 6180 197320 6186
rect 197268 6122 197320 6128
rect 196808 3664 196860 3670
rect 196808 3606 196860 3612
rect 196624 3052 196676 3058
rect 196624 2994 196676 3000
rect 196820 480 196848 3606
rect 198016 3534 198044 24103
rect 198752 11762 198780 158335
rect 198832 152244 198884 152250
rect 198832 152186 198884 152192
rect 198844 144634 198872 152186
rect 198936 148753 198964 158578
rect 199028 152998 199056 158766
rect 199120 158273 199148 159831
rect 199212 158545 199240 160140
rect 199304 159934 199332 160140
rect 199292 159928 199344 159934
rect 199396 159905 199424 160140
rect 199292 159870 199344 159876
rect 199382 159896 199438 159905
rect 199382 159831 199438 159840
rect 199292 159792 199344 159798
rect 199292 159734 199344 159740
rect 199384 159792 199436 159798
rect 199384 159734 199436 159740
rect 199198 158536 199254 158545
rect 199198 158471 199254 158480
rect 199106 158264 199162 158273
rect 199106 158199 199162 158208
rect 199304 158001 199332 159734
rect 199396 158846 199424 159734
rect 199384 158840 199436 158846
rect 199384 158782 199436 158788
rect 199488 158681 199516 160140
rect 199474 158672 199530 158681
rect 199474 158607 199530 158616
rect 199474 158128 199530 158137
rect 199474 158063 199530 158072
rect 199290 157992 199346 158001
rect 199290 157927 199346 157936
rect 199384 157684 199436 157690
rect 199384 157626 199436 157632
rect 199016 152992 199068 152998
rect 199016 152934 199068 152940
rect 198922 148744 198978 148753
rect 198922 148679 198978 148688
rect 199396 145790 199424 157626
rect 199384 145784 199436 145790
rect 199384 145726 199436 145732
rect 199488 145382 199516 158063
rect 199580 157894 199608 160140
rect 199672 159769 199700 160140
rect 199658 159760 199714 159769
rect 199658 159695 199714 159704
rect 199660 158500 199712 158506
rect 199660 158442 199712 158448
rect 199568 157888 199620 157894
rect 199568 157830 199620 157836
rect 199672 150958 199700 158442
rect 199660 150952 199712 150958
rect 199660 150894 199712 150900
rect 199764 147674 199792 160140
rect 199856 157049 199884 160140
rect 199842 157040 199898 157049
rect 199842 156975 199898 156984
rect 199948 152250 199976 160140
rect 200040 158642 200068 160140
rect 200028 158636 200080 158642
rect 200028 158578 200080 158584
rect 200026 158264 200082 158273
rect 200026 158199 200082 158208
rect 199936 152244 199988 152250
rect 199936 152186 199988 152192
rect 199764 147646 199884 147674
rect 199476 145376 199528 145382
rect 199476 145318 199528 145324
rect 198832 144628 198884 144634
rect 198832 144570 198884 144576
rect 199856 129742 199884 147646
rect 199844 129736 199896 129742
rect 199844 129678 199896 129684
rect 198740 11756 198792 11762
rect 198740 11698 198792 11704
rect 200040 10334 200068 158199
rect 200132 156777 200160 160140
rect 200224 159905 200252 160140
rect 200210 159896 200266 159905
rect 200210 159831 200266 159840
rect 200212 159792 200264 159798
rect 200212 159734 200264 159740
rect 200224 159594 200252 159734
rect 200212 159588 200264 159594
rect 200212 159530 200264 159536
rect 200212 158976 200264 158982
rect 200212 158918 200264 158924
rect 200224 157457 200252 158918
rect 200316 158545 200344 160140
rect 200302 158536 200358 158545
rect 200302 158471 200358 158480
rect 200210 157448 200266 157457
rect 200210 157383 200266 157392
rect 200118 156768 200174 156777
rect 200118 156703 200174 156712
rect 200408 155961 200436 160140
rect 200500 158409 200528 160140
rect 200486 158400 200542 158409
rect 200486 158335 200542 158344
rect 200592 157334 200620 160140
rect 200684 158710 200712 160140
rect 200672 158704 200724 158710
rect 200672 158646 200724 158652
rect 200670 157448 200726 157457
rect 200670 157383 200726 157392
rect 200500 157306 200620 157334
rect 200394 155952 200450 155961
rect 200394 155887 200450 155896
rect 200500 152538 200528 157306
rect 200684 157026 200712 157383
rect 200592 156998 200712 157026
rect 200592 154698 200620 156998
rect 200672 156868 200724 156874
rect 200672 156810 200724 156816
rect 200684 156602 200712 156810
rect 200672 156596 200724 156602
rect 200672 156538 200724 156544
rect 200672 155712 200724 155718
rect 200672 155654 200724 155660
rect 200684 155174 200712 155654
rect 200672 155168 200724 155174
rect 200672 155110 200724 155116
rect 200580 154692 200632 154698
rect 200580 154634 200632 154640
rect 200672 154624 200724 154630
rect 200672 154566 200724 154572
rect 200580 153264 200632 153270
rect 200580 153206 200632 153212
rect 200132 152510 200528 152538
rect 200132 126954 200160 152510
rect 200212 152244 200264 152250
rect 200212 152186 200264 152192
rect 200224 143449 200252 152186
rect 200592 147674 200620 153206
rect 200500 147646 200620 147674
rect 200684 147674 200712 154566
rect 200776 152250 200804 160140
rect 200868 158914 200896 160140
rect 200960 159361 200988 160140
rect 200946 159352 201002 159361
rect 200946 159287 201002 159296
rect 200946 158944 201002 158953
rect 200856 158908 200908 158914
rect 200946 158879 201002 158888
rect 200856 158850 200908 158856
rect 200856 158568 200908 158574
rect 200856 158510 200908 158516
rect 200764 152244 200816 152250
rect 200764 152186 200816 152192
rect 200684 147646 200804 147674
rect 200500 145450 200528 147646
rect 200488 145444 200540 145450
rect 200488 145386 200540 145392
rect 200776 145246 200804 147646
rect 200868 147626 200896 158510
rect 200960 157690 200988 158879
rect 201052 158681 201080 160140
rect 201038 158672 201094 158681
rect 201038 158607 201094 158616
rect 200948 157684 201000 157690
rect 200948 157626 201000 157632
rect 200948 157276 201000 157282
rect 200948 157218 201000 157224
rect 200960 156874 200988 157218
rect 200948 156868 201000 156874
rect 200948 156810 201000 156816
rect 200946 155136 201002 155145
rect 200946 155071 201002 155080
rect 200856 147620 200908 147626
rect 200856 147562 200908 147568
rect 200960 145314 200988 155071
rect 201144 151609 201172 160140
rect 201236 159769 201264 160140
rect 201222 159760 201278 159769
rect 201222 159695 201278 159704
rect 201224 158704 201276 158710
rect 201224 158646 201276 158652
rect 201236 154562 201264 158646
rect 201328 158137 201356 160140
rect 201314 158128 201370 158137
rect 201314 158063 201370 158072
rect 201224 154556 201276 154562
rect 201224 154498 201276 154504
rect 201130 151600 201186 151609
rect 201130 151535 201186 151544
rect 201328 147674 201356 158063
rect 201420 148889 201448 160140
rect 201512 155417 201540 160140
rect 201498 155408 201554 155417
rect 201498 155343 201554 155352
rect 201406 148880 201462 148889
rect 201406 148815 201462 148824
rect 201328 147646 201448 147674
rect 200948 145308 201000 145314
rect 200948 145250 201000 145256
rect 200764 145240 200816 145246
rect 200764 145182 200816 145188
rect 200210 143440 200266 143449
rect 200210 143375 200266 143384
rect 201314 143440 201370 143449
rect 201314 143375 201370 143384
rect 201328 143041 201356 143375
rect 201314 143032 201370 143041
rect 201314 142967 201370 142976
rect 200120 126948 200172 126954
rect 200120 126890 200172 126896
rect 201328 108322 201356 142967
rect 200764 108316 200816 108322
rect 200764 108258 200816 108264
rect 201316 108316 201368 108322
rect 201316 108258 201368 108264
rect 200028 10328 200080 10334
rect 200028 10270 200080 10276
rect 200304 4072 200356 4078
rect 200304 4014 200356 4020
rect 198004 3528 198056 3534
rect 198004 3470 198056 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 197912 3052 197964 3058
rect 197912 2994 197964 3000
rect 197924 480 197952 2994
rect 199120 480 199148 3470
rect 200316 480 200344 4014
rect 200776 3058 200804 108258
rect 201420 105602 201448 147646
rect 201604 124166 201632 160140
rect 201696 155174 201724 160140
rect 201788 158506 201816 160140
rect 201880 158545 201908 160140
rect 201866 158536 201922 158545
rect 201776 158500 201828 158506
rect 201866 158471 201922 158480
rect 201776 158442 201828 158448
rect 201972 157334 202000 160140
rect 201788 157306 202000 157334
rect 201684 155168 201736 155174
rect 201684 155110 201736 155116
rect 201684 152244 201736 152250
rect 201684 152186 201736 152192
rect 201696 146266 201724 152186
rect 201788 147558 201816 157306
rect 202064 157185 202092 160140
rect 202156 158681 202184 160140
rect 202248 158760 202276 160140
rect 202340 159089 202368 160140
rect 202432 159769 202460 160140
rect 202418 159760 202474 159769
rect 202418 159695 202474 159704
rect 202326 159080 202382 159089
rect 202326 159015 202382 159024
rect 202248 158732 202368 158760
rect 202142 158672 202198 158681
rect 202142 158607 202198 158616
rect 202144 158568 202196 158574
rect 202144 158510 202196 158516
rect 202156 157865 202184 158510
rect 202234 158264 202290 158273
rect 202234 158199 202290 158208
rect 202142 157856 202198 157865
rect 202142 157791 202198 157800
rect 202144 157752 202196 157758
rect 202144 157694 202196 157700
rect 202156 157593 202184 157694
rect 202142 157584 202198 157593
rect 202142 157519 202198 157528
rect 202248 157282 202276 158199
rect 202236 157276 202288 157282
rect 202236 157218 202288 157224
rect 202050 157176 202106 157185
rect 202050 157111 202106 157120
rect 202236 156936 202288 156942
rect 202236 156878 202288 156884
rect 201960 154760 202012 154766
rect 201960 154702 202012 154708
rect 201972 149734 202000 154702
rect 201960 149728 202012 149734
rect 201960 149670 202012 149676
rect 201776 147552 201828 147558
rect 201776 147494 201828 147500
rect 201684 146260 201736 146266
rect 201684 146202 201736 146208
rect 201592 124160 201644 124166
rect 201592 124102 201644 124108
rect 201408 105596 201460 105602
rect 201408 105538 201460 105544
rect 201972 6914 202000 149670
rect 202248 148442 202276 156878
rect 202340 153066 202368 158732
rect 202420 158228 202472 158234
rect 202420 158170 202472 158176
rect 202328 153060 202380 153066
rect 202328 153002 202380 153008
rect 202236 148436 202288 148442
rect 202236 148378 202288 148384
rect 202432 145586 202460 158170
rect 202524 152250 202552 160140
rect 202616 158574 202644 160140
rect 202708 159769 202736 160140
rect 202694 159760 202750 159769
rect 202694 159695 202750 159704
rect 202696 159520 202748 159526
rect 202696 159462 202748 159468
rect 202708 158574 202736 159462
rect 202604 158568 202656 158574
rect 202604 158510 202656 158516
rect 202696 158568 202748 158574
rect 202696 158510 202748 158516
rect 202800 158273 202828 160140
rect 202892 159905 202920 160140
rect 202878 159896 202934 159905
rect 202878 159831 202934 159840
rect 202786 158264 202842 158273
rect 202786 158199 202842 158208
rect 202786 158128 202842 158137
rect 202786 158063 202788 158072
rect 202840 158063 202842 158072
rect 202788 158034 202840 158040
rect 202604 157956 202656 157962
rect 202788 157956 202840 157962
rect 202656 157916 202788 157944
rect 202604 157898 202656 157904
rect 202788 157898 202840 157904
rect 202788 157276 202840 157282
rect 202788 157218 202840 157224
rect 202696 155168 202748 155174
rect 202696 155110 202748 155116
rect 202512 152244 202564 152250
rect 202512 152186 202564 152192
rect 202708 147674 202736 155110
rect 202800 148617 202828 157218
rect 202880 152176 202932 152182
rect 202880 152118 202932 152124
rect 202786 148608 202842 148617
rect 202786 148543 202842 148552
rect 202708 147646 202828 147674
rect 202420 145580 202472 145586
rect 202420 145522 202472 145528
rect 202694 143440 202750 143449
rect 202694 143375 202750 143384
rect 202708 142186 202736 143375
rect 202696 142180 202748 142186
rect 202696 142122 202748 142128
rect 202708 102814 202736 142122
rect 202696 102808 202748 102814
rect 202696 102750 202748 102756
rect 202800 17270 202828 147646
rect 202892 144702 202920 152118
rect 202984 144809 203012 160140
rect 203076 155854 203104 160140
rect 203064 155848 203116 155854
rect 203064 155790 203116 155796
rect 203064 154692 203116 154698
rect 203064 154634 203116 154640
rect 203076 151774 203104 154634
rect 203168 154193 203196 160140
rect 203260 159939 203288 160140
rect 203246 159930 203302 159939
rect 203246 159865 203302 159874
rect 203248 159792 203300 159798
rect 203248 159734 203300 159740
rect 203260 158166 203288 159734
rect 203352 158760 203380 160140
rect 203444 159934 203472 160140
rect 203432 159928 203484 159934
rect 203432 159870 203484 159876
rect 203352 158732 203472 158760
rect 203340 158568 203392 158574
rect 203340 158510 203392 158516
rect 203248 158160 203300 158166
rect 203248 158102 203300 158108
rect 203154 154184 203210 154193
rect 203154 154119 203210 154128
rect 203352 152250 203380 158510
rect 203444 155145 203472 158732
rect 203536 158409 203564 160140
rect 203522 158400 203578 158409
rect 203522 158335 203578 158344
rect 203430 155136 203486 155145
rect 203430 155071 203486 155080
rect 203340 152244 203392 152250
rect 203340 152186 203392 152192
rect 203064 151768 203116 151774
rect 203064 151710 203116 151716
rect 203628 150385 203656 160140
rect 203720 158302 203748 160140
rect 203812 158681 203840 160140
rect 203798 158672 203854 158681
rect 203798 158607 203854 158616
rect 203708 158296 203760 158302
rect 203708 158238 203760 158244
rect 203706 158128 203762 158137
rect 203706 158063 203762 158072
rect 203614 150376 203670 150385
rect 203614 150311 203670 150320
rect 202970 144800 203026 144809
rect 202970 144735 203026 144744
rect 202880 144696 202932 144702
rect 202880 144638 202932 144644
rect 203720 142154 203748 158063
rect 203800 152244 203852 152250
rect 203800 152186 203852 152192
rect 203812 143274 203840 152186
rect 203904 152182 203932 160140
rect 203996 158953 204024 160140
rect 204088 159905 204116 160140
rect 204074 159896 204130 159905
rect 204074 159831 204130 159840
rect 204076 159588 204128 159594
rect 204076 159530 204128 159536
rect 203982 158944 204038 158953
rect 203982 158879 204038 158888
rect 203982 158808 204038 158817
rect 203982 158743 204038 158752
rect 203892 152176 203944 152182
rect 203892 152118 203944 152124
rect 203890 144800 203946 144809
rect 203890 144735 203946 144744
rect 203800 143268 203852 143274
rect 203800 143210 203852 143216
rect 203628 142126 203748 142154
rect 203628 28286 203656 142126
rect 203904 122126 203932 144735
rect 203892 122120 203944 122126
rect 203892 122062 203944 122068
rect 203996 94518 204024 158743
rect 204088 158642 204116 159530
rect 204076 158636 204128 158642
rect 204076 158578 204128 158584
rect 204180 158545 204208 160140
rect 204272 159905 204300 160140
rect 204258 159896 204314 159905
rect 204258 159831 204314 159840
rect 204260 158704 204312 158710
rect 204260 158646 204312 158652
rect 204166 158536 204222 158545
rect 204166 158471 204222 158480
rect 204168 158296 204220 158302
rect 204168 158238 204220 158244
rect 204074 155136 204130 155145
rect 204074 155071 204130 155080
rect 203984 94512 204036 94518
rect 203984 94454 204036 94460
rect 204088 36582 204116 155071
rect 204180 152833 204208 158238
rect 204272 158234 204300 158646
rect 204260 158228 204312 158234
rect 204260 158170 204312 158176
rect 204258 154592 204314 154601
rect 204258 154527 204314 154536
rect 204166 152824 204222 152833
rect 204166 152759 204222 152768
rect 204272 150346 204300 154527
rect 204364 153270 204392 160140
rect 204352 153264 204404 153270
rect 204352 153206 204404 153212
rect 204456 153202 204484 160140
rect 204548 158273 204576 160140
rect 204640 159769 204668 160140
rect 204626 159760 204682 159769
rect 204626 159695 204682 159704
rect 204534 158264 204590 158273
rect 204534 158199 204590 158208
rect 204640 157334 204668 159695
rect 204548 157306 204668 157334
rect 204444 153196 204496 153202
rect 204444 153138 204496 153144
rect 204548 152538 204576 157306
rect 204628 153264 204680 153270
rect 204628 153206 204680 153212
rect 204364 152510 204576 152538
rect 204260 150340 204312 150346
rect 204260 150282 204312 150288
rect 204364 93158 204392 152510
rect 204640 152266 204668 153206
rect 204456 152238 204668 152266
rect 204456 143070 204484 152238
rect 204732 149025 204760 160140
rect 204824 158098 204852 160140
rect 204916 159905 204944 160140
rect 204902 159896 204958 159905
rect 204902 159831 204958 159840
rect 204812 158092 204864 158098
rect 204812 158034 204864 158040
rect 204916 157334 204944 159831
rect 205008 158681 205036 160140
rect 204994 158672 205050 158681
rect 204994 158607 205050 158616
rect 205100 158409 205128 160140
rect 205192 159905 205220 160140
rect 205178 159896 205234 159905
rect 205178 159831 205234 159840
rect 205180 159520 205232 159526
rect 205180 159462 205232 159468
rect 205086 158400 205142 158409
rect 205086 158335 205142 158344
rect 204824 157306 204944 157334
rect 204824 152250 204852 157306
rect 205192 154465 205220 159462
rect 205178 154456 205234 154465
rect 205178 154391 205234 154400
rect 205284 152538 205312 160140
rect 205376 159526 205404 160140
rect 205468 159905 205496 160140
rect 205454 159896 205510 159905
rect 205454 159831 205510 159840
rect 205364 159520 205416 159526
rect 205364 159462 205416 159468
rect 205364 158092 205416 158098
rect 205364 158034 205416 158040
rect 205376 155553 205404 158034
rect 205362 155544 205418 155553
rect 205362 155479 205418 155488
rect 205364 153264 205416 153270
rect 205364 153206 205416 153212
rect 204916 152510 205312 152538
rect 204812 152244 204864 152250
rect 204812 152186 204864 152192
rect 204718 149016 204774 149025
rect 204718 148951 204774 148960
rect 204444 143064 204496 143070
rect 204444 143006 204496 143012
rect 204916 141914 204944 152510
rect 205376 147674 205404 153206
rect 205468 152538 205496 159831
rect 205560 153270 205588 160140
rect 205652 157554 205680 160140
rect 205640 157548 205692 157554
rect 205640 157490 205692 157496
rect 205638 157448 205694 157457
rect 205638 157383 205694 157392
rect 205548 153264 205600 153270
rect 205548 153206 205600 153212
rect 205468 152510 205588 152538
rect 205456 152244 205508 152250
rect 205456 152186 205508 152192
rect 205192 147646 205404 147674
rect 204904 141908 204956 141914
rect 204904 141850 204956 141856
rect 205192 137902 205220 147646
rect 205272 143064 205324 143070
rect 205272 143006 205324 143012
rect 205284 142866 205312 143006
rect 205272 142860 205324 142866
rect 205272 142802 205324 142808
rect 205180 137896 205232 137902
rect 205180 137838 205232 137844
rect 205284 120766 205312 142802
rect 205272 120760 205324 120766
rect 205272 120702 205324 120708
rect 204352 93152 204404 93158
rect 204352 93094 204404 93100
rect 205468 91798 205496 152186
rect 205456 91792 205508 91798
rect 204258 91760 204314 91769
rect 205456 91734 205508 91740
rect 204258 91695 204314 91704
rect 204076 36576 204128 36582
rect 204076 36518 204128 36524
rect 203616 28280 203668 28286
rect 203616 28222 203668 28228
rect 202788 17264 202840 17270
rect 202788 17206 202840 17212
rect 204272 16574 204300 91695
rect 205560 87650 205588 152510
rect 205652 151814 205680 157383
rect 205744 155972 205772 160140
rect 205836 157944 205864 160140
rect 205928 158817 205956 160140
rect 206020 159225 206048 160140
rect 206006 159216 206062 159225
rect 206006 159151 206062 159160
rect 205914 158808 205970 158817
rect 205914 158743 205970 158752
rect 206020 158137 206048 159151
rect 206006 158128 206062 158137
rect 206006 158063 206062 158072
rect 205836 157916 205956 157944
rect 205824 157548 205876 157554
rect 205824 157490 205876 157496
rect 205836 156942 205864 157490
rect 205824 156936 205876 156942
rect 205824 156878 205876 156884
rect 205744 155944 205864 155972
rect 205652 151786 205772 151814
rect 205744 136610 205772 151786
rect 205836 144362 205864 155944
rect 205928 154329 205956 157916
rect 205914 154320 205970 154329
rect 205914 154255 205970 154264
rect 206112 147665 206140 160140
rect 206204 159934 206232 160140
rect 206192 159928 206244 159934
rect 206296 159905 206324 160140
rect 206192 159870 206244 159876
rect 206282 159896 206338 159905
rect 206282 159831 206338 159840
rect 206284 159792 206336 159798
rect 206284 159734 206336 159740
rect 206192 159520 206244 159526
rect 206192 159462 206244 159468
rect 206204 157214 206232 159462
rect 206296 158098 206324 159734
rect 206284 158092 206336 158098
rect 206284 158034 206336 158040
rect 206192 157208 206244 157214
rect 206192 157150 206244 157156
rect 206388 156074 206416 160140
rect 206480 158545 206508 160140
rect 206572 158681 206600 160140
rect 206558 158672 206614 158681
rect 206558 158607 206614 158616
rect 206466 158536 206522 158545
rect 206466 158471 206522 158480
rect 206558 158128 206614 158137
rect 206558 158063 206614 158072
rect 206388 156046 206508 156074
rect 206376 155984 206428 155990
rect 206376 155926 206428 155932
rect 206098 147656 206154 147665
rect 206098 147591 206154 147600
rect 205824 144356 205876 144362
rect 205824 144298 205876 144304
rect 205732 136604 205784 136610
rect 205732 136546 205784 136552
rect 206388 135250 206416 155926
rect 206480 155281 206508 156046
rect 206466 155272 206522 155281
rect 206466 155207 206522 155216
rect 206376 135244 206428 135250
rect 206376 135186 206428 135192
rect 205548 87644 205600 87650
rect 205548 87586 205600 87592
rect 206572 86290 206600 158063
rect 206664 157457 206692 160140
rect 206756 159225 206784 160140
rect 206848 159769 206876 160140
rect 206834 159760 206890 159769
rect 206834 159695 206890 159704
rect 206742 159216 206798 159225
rect 206742 159151 206798 159160
rect 206742 157584 206798 157593
rect 206742 157519 206798 157528
rect 206650 157448 206706 157457
rect 206650 157383 206706 157392
rect 206756 157334 206784 157519
rect 206664 157306 206784 157334
rect 206664 151814 206692 157306
rect 206940 155990 206968 160140
rect 207032 159934 207060 160140
rect 207020 159928 207072 159934
rect 207020 159870 207072 159876
rect 207124 159866 207152 160140
rect 207112 159860 207164 159866
rect 207112 159802 207164 159808
rect 207018 159760 207074 159769
rect 207018 159695 207074 159704
rect 207032 159594 207060 159695
rect 207020 159588 207072 159594
rect 207020 159530 207072 159536
rect 207020 157956 207072 157962
rect 207020 157898 207072 157904
rect 207032 156330 207060 157898
rect 207124 157894 207152 159802
rect 207216 158137 207244 160140
rect 207308 159905 207336 160140
rect 207294 159896 207350 159905
rect 207294 159831 207350 159840
rect 207400 159769 207428 160140
rect 207584 159866 207612 164206
rect 207676 161514 207704 241538
rect 207756 238604 207808 238610
rect 207756 238546 207808 238552
rect 207768 161650 207796 238546
rect 207860 235210 207888 298250
rect 207952 241369 207980 308586
rect 208124 304496 208176 304502
rect 208124 304438 208176 304444
rect 208032 304360 208084 304366
rect 208032 304302 208084 304308
rect 207938 241360 207994 241369
rect 207938 241295 207994 241304
rect 208044 235890 208072 304302
rect 208032 235884 208084 235890
rect 208032 235826 208084 235832
rect 207848 235204 207900 235210
rect 207848 235146 207900 235152
rect 208136 233073 208164 304438
rect 208228 238105 208256 318854
rect 208214 238096 208270 238105
rect 208214 238031 208270 238040
rect 208122 233064 208178 233073
rect 208122 232999 208178 233008
rect 208320 229090 208348 320894
rect 209504 320884 209556 320890
rect 209504 320826 209556 320832
rect 209412 311160 209464 311166
rect 209412 311102 209464 311108
rect 209228 306400 209280 306406
rect 209228 306342 209280 306348
rect 209044 299736 209096 299742
rect 209044 299678 209096 299684
rect 208308 229084 208360 229090
rect 208308 229026 208360 229032
rect 208320 228886 208348 229026
rect 208308 228880 208360 228886
rect 208308 228822 208360 228828
rect 209056 216102 209084 299678
rect 209136 297424 209188 297430
rect 209136 297366 209188 297372
rect 209044 216096 209096 216102
rect 209044 216038 209096 216044
rect 209148 213450 209176 297366
rect 209240 241534 209268 306342
rect 209228 241528 209280 241534
rect 209228 241470 209280 241476
rect 209240 238746 209268 241470
rect 209424 238921 209452 311102
rect 209410 238912 209466 238921
rect 209410 238847 209466 238856
rect 209228 238740 209280 238746
rect 209228 238682 209280 238688
rect 209320 238468 209372 238474
rect 209320 238410 209372 238416
rect 209228 235612 209280 235618
rect 209228 235554 209280 235560
rect 209136 213444 209188 213450
rect 209136 213386 209188 213392
rect 209136 207800 209188 207806
rect 209136 207742 209188 207748
rect 209044 207664 209096 207670
rect 209044 207606 209096 207612
rect 207846 188320 207902 188329
rect 207846 188255 207902 188264
rect 207860 166994 207888 188255
rect 207938 184240 207994 184249
rect 207938 184175 207994 184184
rect 207952 169130 207980 184175
rect 208030 176080 208086 176089
rect 208030 176015 208086 176024
rect 208044 171134 208072 176015
rect 208952 173188 209004 173194
rect 208952 173130 209004 173136
rect 208044 171106 208256 171134
rect 207952 169102 208164 169130
rect 208030 169008 208086 169017
rect 208030 168943 208086 168952
rect 207860 166966 207980 166994
rect 207952 161786 207980 166966
rect 208044 161922 208072 168943
rect 208136 162058 208164 169102
rect 208228 166994 208256 171106
rect 208228 166966 208348 166994
rect 208136 162030 208256 162058
rect 208044 161894 208164 161922
rect 207952 161758 208072 161786
rect 207768 161622 207980 161650
rect 207676 161486 207888 161514
rect 207754 161256 207810 161265
rect 207754 161191 207810 161200
rect 207664 161152 207716 161158
rect 207664 161094 207716 161100
rect 207572 159860 207624 159866
rect 207572 159802 207624 159808
rect 207386 159760 207442 159769
rect 207386 159695 207442 159704
rect 207400 158574 207428 159695
rect 207480 159588 207532 159594
rect 207480 159530 207532 159536
rect 207388 158568 207440 158574
rect 207388 158510 207440 158516
rect 207202 158128 207258 158137
rect 207202 158063 207258 158072
rect 207492 158030 207520 159530
rect 207676 158710 207704 161094
rect 207768 160002 207796 161191
rect 207860 160070 207888 161486
rect 207848 160064 207900 160070
rect 207848 160006 207900 160012
rect 207756 159996 207808 160002
rect 207756 159938 207808 159944
rect 207952 159458 207980 161622
rect 207940 159452 207992 159458
rect 207940 159394 207992 159400
rect 207664 158704 207716 158710
rect 207664 158646 207716 158652
rect 207848 158296 207900 158302
rect 207848 158238 207900 158244
rect 207480 158024 207532 158030
rect 207480 157966 207532 157972
rect 207112 157888 207164 157894
rect 207112 157830 207164 157836
rect 207204 157548 207256 157554
rect 207204 157490 207256 157496
rect 207020 156324 207072 156330
rect 207020 156266 207072 156272
rect 206928 155984 206980 155990
rect 206928 155926 206980 155932
rect 207216 155718 207244 157490
rect 207204 155712 207256 155718
rect 207204 155654 207256 155660
rect 207860 155378 207888 158238
rect 208044 158234 208072 161758
rect 208136 160138 208164 161894
rect 208124 160132 208176 160138
rect 208124 160074 208176 160080
rect 208228 159594 208256 162030
rect 208320 159798 208348 166966
rect 208858 164792 208914 164801
rect 208858 164727 208914 164736
rect 208400 161016 208452 161022
rect 208400 160958 208452 160964
rect 208412 160206 208440 160958
rect 208400 160200 208452 160206
rect 208400 160142 208452 160148
rect 208308 159792 208360 159798
rect 208308 159734 208360 159740
rect 208216 159588 208268 159594
rect 208216 159530 208268 159536
rect 208308 158568 208360 158574
rect 208308 158510 208360 158516
rect 208032 158228 208084 158234
rect 208032 158170 208084 158176
rect 207940 158160 207992 158166
rect 207940 158102 207992 158108
rect 208122 158128 208178 158137
rect 207848 155372 207900 155378
rect 207848 155314 207900 155320
rect 206926 155272 206982 155281
rect 206926 155207 206982 155216
rect 206664 151786 206876 151814
rect 206652 144356 206704 144362
rect 206652 144298 206704 144304
rect 206664 89010 206692 144298
rect 206652 89004 206704 89010
rect 206652 88946 206704 88952
rect 206560 86284 206612 86290
rect 206560 86226 206612 86232
rect 206848 82142 206876 151786
rect 206836 82136 206888 82142
rect 206836 82078 206888 82084
rect 206940 33794 206968 155207
rect 207952 154970 207980 158102
rect 208032 158092 208084 158098
rect 208122 158063 208178 158072
rect 208032 158034 208084 158040
rect 207940 154964 207992 154970
rect 207940 154906 207992 154912
rect 208044 154902 208072 158034
rect 208032 154896 208084 154902
rect 208032 154838 208084 154844
rect 208136 133210 208164 158063
rect 208216 157888 208268 157894
rect 208216 157830 208268 157836
rect 208124 133204 208176 133210
rect 208124 133146 208176 133152
rect 208228 83502 208256 157830
rect 208216 83496 208268 83502
rect 208216 83438 208268 83444
rect 208320 80714 208348 158510
rect 208872 158438 208900 164727
rect 208964 160449 208992 173130
rect 208950 160440 209006 160449
rect 208950 160375 209006 160384
rect 208860 158432 208912 158438
rect 209056 158409 209084 207606
rect 209148 160274 209176 207742
rect 209136 160268 209188 160274
rect 209136 160210 209188 160216
rect 208860 158374 208912 158380
rect 209042 158400 209098 158409
rect 209042 158335 209098 158344
rect 208400 158228 208452 158234
rect 208400 158170 208452 158176
rect 208412 157350 208440 158170
rect 208492 158024 208544 158030
rect 208492 157966 208544 157972
rect 208674 157992 208730 158001
rect 208400 157344 208452 157350
rect 208400 157286 208452 157292
rect 208504 156641 208532 157966
rect 208674 157927 208730 157936
rect 208490 156632 208546 156641
rect 208490 156567 208546 156576
rect 208400 153808 208452 153814
rect 208400 153750 208452 153756
rect 208308 80708 208360 80714
rect 208308 80650 208360 80656
rect 205640 33788 205692 33794
rect 205640 33730 205692 33736
rect 206928 33788 206980 33794
rect 206928 33730 206980 33736
rect 205652 16574 205680 33730
rect 208412 16574 208440 153750
rect 208688 153649 208716 157927
rect 209240 156874 209268 235554
rect 209332 159662 209360 238410
rect 209424 232830 209452 238847
rect 209412 232824 209464 232830
rect 209412 232766 209464 232772
rect 209516 231810 209544 320826
rect 209594 315344 209650 315353
rect 209594 315279 209650 315288
rect 209504 231804 209556 231810
rect 209504 231746 209556 231752
rect 209516 228818 209544 231746
rect 209504 228812 209556 228818
rect 209504 228754 209556 228760
rect 209412 224324 209464 224330
rect 209412 224266 209464 224272
rect 209320 159656 209372 159662
rect 209320 159598 209372 159604
rect 209228 156868 209280 156874
rect 209228 156810 209280 156816
rect 209424 153814 209452 224266
rect 209608 222873 209636 315279
rect 209700 224913 209728 322254
rect 212448 322244 212500 322250
rect 212448 322186 212500 322192
rect 211066 319560 211122 319569
rect 211066 319495 211122 319504
rect 210790 318064 210846 318073
rect 210790 317999 210846 318008
rect 210608 312588 210660 312594
rect 210608 312530 210660 312536
rect 210238 307864 210294 307873
rect 210238 307799 210294 307808
rect 210252 233753 210280 307799
rect 210516 243500 210568 243506
rect 210516 243442 210568 243448
rect 210424 239896 210476 239902
rect 210424 239838 210476 239844
rect 210332 238536 210384 238542
rect 210332 238478 210384 238484
rect 210238 233744 210294 233753
rect 210238 233679 210294 233688
rect 209686 224904 209742 224913
rect 209686 224839 209742 224848
rect 209594 222864 209650 222873
rect 209594 222799 209650 222808
rect 209504 207732 209556 207738
rect 209504 207674 209556 207680
rect 209516 158273 209544 207674
rect 209596 202156 209648 202162
rect 209596 202098 209648 202104
rect 209502 158264 209558 158273
rect 209502 158199 209558 158208
rect 209608 157690 209636 202098
rect 209688 177336 209740 177342
rect 209688 177278 209740 177284
rect 209700 159934 209728 177278
rect 210344 166994 210372 238478
rect 210160 166966 210372 166994
rect 209780 164892 209832 164898
rect 209780 164834 209832 164840
rect 209792 164801 209820 164834
rect 209778 164792 209834 164801
rect 209778 164727 209834 164736
rect 209688 159928 209740 159934
rect 209688 159870 209740 159876
rect 210160 159322 210188 166966
rect 210238 161256 210294 161265
rect 210238 161191 210294 161200
rect 210252 160313 210280 161191
rect 210238 160304 210294 160313
rect 210238 160239 210294 160248
rect 210148 159316 210200 159322
rect 210148 159258 210200 159264
rect 209596 157684 209648 157690
rect 209596 157626 209648 157632
rect 209688 156800 209740 156806
rect 209688 156742 209740 156748
rect 209412 153808 209464 153814
rect 209412 153750 209464 153756
rect 208674 153640 208730 153649
rect 208674 153575 208730 153584
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 208412 16546 208624 16574
rect 201512 6886 202000 6914
rect 200764 3052 200816 3058
rect 200764 2994 200816 3000
rect 201512 480 201540 6886
rect 203890 3632 203946 3641
rect 203890 3567 203946 3576
rect 202696 3052 202748 3058
rect 202696 2994 202748 3000
rect 202708 480 202736 2994
rect 203904 480 203932 3567
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207388 3460 207440 3466
rect 207388 3402 207440 3408
rect 207400 480 207428 3402
rect 208596 480 208624 16546
rect 209700 4146 209728 156742
rect 210436 155446 210464 239838
rect 210424 155440 210476 155446
rect 210424 155382 210476 155388
rect 209872 152516 209924 152522
rect 209872 152458 209924 152464
rect 209884 6914 209912 152458
rect 209792 6886 209912 6914
rect 209688 4140 209740 4146
rect 209688 4082 209740 4088
rect 209792 480 209820 6886
rect 210436 3466 210464 155382
rect 210528 152318 210556 243442
rect 210620 240961 210648 312530
rect 210700 305720 210752 305726
rect 210700 305662 210752 305668
rect 210606 240952 210662 240961
rect 210606 240887 210662 240896
rect 210712 239601 210740 305662
rect 210698 239592 210754 239601
rect 210698 239527 210754 239536
rect 210712 239329 210740 239527
rect 210698 239320 210754 239329
rect 210698 239255 210754 239264
rect 210698 238640 210754 238649
rect 210698 238575 210754 238584
rect 210608 235748 210660 235754
rect 210608 235690 210660 235696
rect 210620 152386 210648 235690
rect 210712 235634 210740 238575
rect 210804 238241 210832 317999
rect 210882 315752 210938 315761
rect 210882 315687 210938 315696
rect 210790 238232 210846 238241
rect 210790 238167 210846 238176
rect 210712 235606 210832 235634
rect 210700 235476 210752 235482
rect 210700 235418 210752 235424
rect 210712 154494 210740 235418
rect 210804 234190 210832 235606
rect 210896 235521 210924 315687
rect 210976 314016 211028 314022
rect 210976 313958 211028 313964
rect 210988 238649 211016 313958
rect 211080 239873 211108 319495
rect 212172 316804 212224 316810
rect 212172 316746 212224 316752
rect 211896 313948 211948 313954
rect 211896 313890 211948 313896
rect 211804 297288 211856 297294
rect 211804 297230 211856 297236
rect 211066 239864 211122 239873
rect 211066 239799 211122 239808
rect 210974 238640 211030 238649
rect 210974 238575 211030 238584
rect 211080 238320 211108 239799
rect 210988 238292 211108 238320
rect 210882 235512 210938 235521
rect 210882 235447 210938 235456
rect 210792 234184 210844 234190
rect 210792 234126 210844 234132
rect 210988 227050 211016 238292
rect 211066 238232 211122 238241
rect 211066 238167 211122 238176
rect 211080 237425 211108 238167
rect 211066 237416 211122 237425
rect 211066 237351 211122 237360
rect 211620 235680 211672 235686
rect 211620 235622 211672 235628
rect 211066 234560 211122 234569
rect 211066 234495 211122 234504
rect 211080 233753 211108 234495
rect 211066 233744 211122 233753
rect 211066 233679 211122 233688
rect 210976 227044 211028 227050
rect 210976 226986 211028 226992
rect 210792 206304 210844 206310
rect 210792 206246 210844 206252
rect 210804 157758 210832 206246
rect 210884 196648 210936 196654
rect 210884 196590 210936 196596
rect 210792 157752 210844 157758
rect 210792 157694 210844 157700
rect 210896 157622 210924 196590
rect 210976 192500 211028 192506
rect 210976 192442 211028 192448
rect 210988 157729 211016 192442
rect 211068 186992 211120 186998
rect 211068 186934 211120 186940
rect 210974 157720 211030 157729
rect 210974 157655 211030 157664
rect 210884 157616 210936 157622
rect 210884 157558 210936 157564
rect 211080 157418 211108 186934
rect 211068 157412 211120 157418
rect 211068 157354 211120 157360
rect 210700 154488 210752 154494
rect 210700 154430 210752 154436
rect 211160 153876 211212 153882
rect 211160 153818 211212 153824
rect 210608 152380 210660 152386
rect 210608 152322 210660 152328
rect 210516 152312 210568 152318
rect 210516 152254 210568 152260
rect 211172 16574 211200 153818
rect 211632 150890 211660 235622
rect 211712 227044 211764 227050
rect 211712 226986 211764 226992
rect 211724 155961 211752 226986
rect 211816 212362 211844 297230
rect 211908 234530 211936 313890
rect 211986 298752 212042 298761
rect 211986 298687 212042 298696
rect 212000 237289 212028 298687
rect 212080 294160 212132 294166
rect 212080 294102 212132 294108
rect 211986 237280 212042 237289
rect 211986 237215 212042 237224
rect 211896 234524 211948 234530
rect 211896 234466 211948 234472
rect 211804 212356 211856 212362
rect 211804 212298 211856 212304
rect 211804 156596 211856 156602
rect 211804 156538 211856 156544
rect 211710 155952 211766 155961
rect 211710 155887 211766 155896
rect 211620 150884 211672 150890
rect 211620 150826 211672 150832
rect 211172 16546 211752 16574
rect 210976 4140 211028 4146
rect 210976 4082 211028 4088
rect 210424 3460 210476 3466
rect 210424 3402 210476 3408
rect 210988 480 211016 4082
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 211816 3738 211844 156538
rect 211908 146985 211936 234466
rect 212000 234122 212028 237215
rect 211988 234116 212040 234122
rect 211988 234058 212040 234064
rect 212092 210730 212120 294102
rect 212184 239358 212212 316746
rect 212356 316736 212408 316742
rect 212356 316678 212408 316684
rect 212264 293208 212316 293214
rect 212264 293150 212316 293156
rect 212172 239352 212224 239358
rect 212172 239294 212224 239300
rect 212172 236904 212224 236910
rect 212172 236846 212224 236852
rect 212080 210724 212132 210730
rect 212080 210666 212132 210672
rect 212184 153882 212212 236846
rect 212276 212090 212304 293150
rect 212368 236026 212396 316678
rect 212356 236020 212408 236026
rect 212356 235962 212408 235968
rect 212460 233238 212488 322186
rect 219346 321736 219402 321745
rect 216588 321700 216640 321706
rect 219346 321671 219402 321680
rect 216588 321642 216640 321648
rect 216404 320204 216456 320210
rect 216404 320146 216456 320152
rect 213092 319796 213144 319802
rect 213092 319738 213144 319744
rect 212906 239592 212962 239601
rect 212906 239527 212962 239536
rect 212540 234592 212592 234598
rect 212540 234534 212592 234540
rect 212552 234190 212580 234534
rect 212540 234184 212592 234190
rect 212540 234126 212592 234132
rect 212448 233232 212500 233238
rect 212448 233174 212500 233180
rect 212448 230172 212500 230178
rect 212448 230114 212500 230120
rect 212356 229560 212408 229566
rect 212356 229502 212408 229508
rect 212264 212084 212316 212090
rect 212264 212026 212316 212032
rect 212368 156602 212396 229502
rect 212356 156596 212408 156602
rect 212356 156538 212408 156544
rect 212460 155106 212488 230114
rect 212448 155100 212500 155106
rect 212448 155042 212500 155048
rect 212172 153876 212224 153882
rect 212172 153818 212224 153824
rect 211894 146976 211950 146985
rect 211894 146911 211950 146920
rect 212552 146305 212580 234126
rect 212920 152590 212948 239527
rect 213000 239080 213052 239086
rect 213000 239022 213052 239028
rect 213012 153950 213040 239022
rect 213104 236881 213132 319738
rect 215206 319696 215262 319705
rect 215206 319631 215262 319640
rect 213736 319524 213788 319530
rect 213736 319466 213788 319472
rect 213552 316872 213604 316878
rect 213552 316814 213604 316820
rect 213460 315376 213512 315382
rect 213460 315318 213512 315324
rect 213368 307216 213420 307222
rect 213368 307158 213420 307164
rect 213276 304292 213328 304298
rect 213276 304234 213328 304240
rect 213288 240417 213316 304234
rect 213274 240408 213330 240417
rect 213274 240343 213330 240352
rect 213184 240236 213236 240242
rect 213184 240178 213236 240184
rect 213090 236872 213146 236881
rect 213090 236807 213146 236816
rect 213196 157078 213224 240178
rect 213288 236842 213316 240343
rect 213276 236836 213328 236842
rect 213276 236778 213328 236784
rect 213380 236638 213408 307158
rect 213472 240145 213500 315318
rect 213458 240136 213514 240145
rect 213458 240071 213514 240080
rect 213472 239465 213500 240071
rect 213458 239456 213514 239465
rect 213458 239391 213514 239400
rect 213460 237312 213512 237318
rect 213460 237254 213512 237260
rect 213368 236632 213420 236638
rect 213368 236574 213420 236580
rect 213184 157072 213236 157078
rect 213184 157014 213236 157020
rect 213184 155100 213236 155106
rect 213184 155042 213236 155048
rect 213000 153944 213052 153950
rect 213000 153886 213052 153892
rect 212908 152584 212960 152590
rect 212908 152526 212960 152532
rect 212538 146296 212594 146305
rect 212538 146231 212594 146240
rect 212538 144120 212594 144129
rect 212538 144055 212594 144064
rect 212552 16574 212580 144055
rect 212552 16546 213132 16574
rect 211804 3732 211856 3738
rect 211804 3674 211856 3680
rect 213104 3482 213132 16546
rect 213196 3806 213224 155042
rect 213472 152289 213500 237254
rect 213564 236065 213592 316814
rect 213644 315512 213696 315518
rect 213644 315454 213696 315460
rect 213550 236056 213606 236065
rect 213550 235991 213606 236000
rect 213656 235929 213684 315454
rect 213748 243386 213776 319466
rect 215114 316840 215170 316849
rect 215114 316775 215170 316784
rect 214930 315888 214986 315897
rect 214930 315823 214986 315832
rect 214840 305652 214892 305658
rect 214840 305594 214892 305600
rect 213828 303000 213880 303006
rect 213828 302942 213880 302948
rect 213840 243522 213868 302942
rect 214748 295860 214800 295866
rect 214748 295802 214800 295808
rect 214656 295452 214708 295458
rect 214656 295394 214708 295400
rect 214564 291916 214616 291922
rect 214564 291858 214616 291864
rect 213840 243506 213960 243522
rect 213828 243500 213960 243506
rect 213880 243494 213960 243500
rect 213828 243442 213880 243448
rect 213748 243358 213868 243386
rect 213736 240508 213788 240514
rect 213736 240450 213788 240456
rect 213642 235920 213698 235929
rect 213642 235855 213698 235864
rect 213656 235385 213684 235855
rect 213642 235376 213698 235385
rect 213642 235311 213698 235320
rect 213748 229094 213776 240450
rect 213840 237017 213868 243358
rect 213932 241058 213960 243494
rect 214576 242214 214604 291858
rect 214564 242208 214616 242214
rect 214564 242150 214616 242156
rect 213920 241052 213972 241058
rect 213920 240994 213972 241000
rect 214472 240372 214524 240378
rect 214472 240314 214524 240320
rect 213826 237008 213882 237017
rect 213826 236943 213882 236952
rect 213840 236042 213868 236943
rect 213840 236014 214144 236042
rect 214012 235952 214064 235958
rect 214012 235894 214064 235900
rect 213748 229066 213868 229094
rect 213736 228812 213788 228818
rect 213736 228754 213788 228760
rect 213458 152280 213514 152289
rect 213458 152215 213514 152224
rect 213748 149802 213776 228754
rect 213840 157026 213868 229066
rect 213840 157010 213960 157026
rect 213840 157004 213972 157010
rect 213840 156998 213920 157004
rect 213920 156946 213972 156952
rect 213736 149796 213788 149802
rect 213736 149738 213788 149744
rect 213748 149122 213776 149738
rect 213736 149116 213788 149122
rect 213736 149058 213788 149064
rect 213932 16574 213960 156946
rect 214024 149530 214052 235894
rect 214116 149841 214144 236014
rect 214484 229094 214512 240314
rect 214484 229066 214604 229094
rect 214194 222864 214250 222873
rect 214194 222799 214250 222808
rect 214102 149832 214158 149841
rect 214102 149767 214158 149776
rect 214012 149524 214064 149530
rect 214012 149466 214064 149472
rect 214208 145897 214236 222799
rect 214576 152726 214604 229066
rect 214668 213382 214696 295394
rect 214760 214810 214788 295802
rect 214852 241194 214880 305594
rect 214944 251666 214972 315823
rect 215024 294092 215076 294098
rect 215024 294034 215076 294040
rect 214932 251660 214984 251666
rect 214932 251602 214984 251608
rect 214840 241188 214892 241194
rect 214840 241130 214892 241136
rect 214852 240242 214880 241130
rect 214840 240236 214892 240242
rect 214840 240178 214892 240184
rect 214840 236972 214892 236978
rect 214840 236914 214892 236920
rect 214852 236026 214880 236914
rect 214932 236836 214984 236842
rect 214932 236778 214984 236784
rect 214840 236020 214892 236026
rect 214840 235962 214892 235968
rect 214840 235544 214892 235550
rect 214840 235486 214892 235492
rect 214748 214804 214800 214810
rect 214748 214746 214800 214752
rect 214656 213376 214708 213382
rect 214656 213318 214708 213324
rect 214852 155786 214880 235486
rect 214944 157554 214972 236778
rect 215036 217394 215064 294034
rect 215128 239562 215156 316775
rect 215220 239970 215248 319631
rect 216312 319592 216364 319598
rect 216312 319534 216364 319540
rect 216128 307896 216180 307902
rect 216128 307838 216180 307844
rect 216036 305108 216088 305114
rect 216036 305050 216088 305056
rect 215944 302932 215996 302938
rect 215944 302874 215996 302880
rect 215852 291780 215904 291786
rect 215852 291722 215904 291728
rect 215668 251660 215720 251666
rect 215668 251602 215720 251608
rect 215680 241534 215708 251602
rect 215864 249082 215892 291722
rect 215852 249076 215904 249082
rect 215852 249018 215904 249024
rect 215668 241528 215720 241534
rect 215668 241470 215720 241476
rect 215208 239964 215260 239970
rect 215208 239906 215260 239912
rect 215116 239556 215168 239562
rect 215116 239498 215168 239504
rect 215128 236774 215156 239498
rect 215116 236768 215168 236774
rect 215116 236710 215168 236716
rect 215220 228954 215248 239906
rect 215390 236056 215446 236065
rect 215390 235991 215446 236000
rect 215208 228948 215260 228954
rect 215208 228890 215260 228896
rect 215116 227588 215168 227594
rect 215116 227530 215168 227536
rect 215024 217388 215076 217394
rect 215024 217330 215076 217336
rect 214932 157548 214984 157554
rect 214932 157490 214984 157496
rect 214840 155780 214892 155786
rect 214840 155722 214892 155728
rect 215128 154562 215156 227530
rect 215404 219434 215432 235991
rect 215680 235249 215708 241470
rect 215852 240576 215904 240582
rect 215852 240518 215904 240524
rect 215864 239018 215892 240518
rect 215852 239012 215904 239018
rect 215852 238954 215904 238960
rect 215666 235240 215722 235249
rect 215666 235175 215722 235184
rect 215312 219406 215432 219434
rect 215116 154556 215168 154562
rect 215116 154498 215168 154504
rect 214564 152720 214616 152726
rect 214564 152662 214616 152668
rect 215312 149977 215340 219406
rect 215864 156806 215892 238954
rect 215956 238134 215984 302874
rect 216048 253910 216076 305050
rect 216036 253904 216088 253910
rect 216036 253846 216088 253852
rect 216140 241330 216168 307838
rect 216220 307828 216272 307834
rect 216220 307770 216272 307776
rect 216128 241324 216180 241330
rect 216128 241266 216180 241272
rect 216140 240378 216168 241266
rect 216128 240372 216180 240378
rect 216128 240314 216180 240320
rect 216036 240236 216088 240242
rect 216036 240178 216088 240184
rect 215944 238128 215996 238134
rect 215944 238070 215996 238076
rect 215944 234660 215996 234666
rect 215944 234602 215996 234608
rect 215852 156800 215904 156806
rect 215852 156742 215904 156748
rect 215956 150414 215984 234602
rect 216048 155514 216076 240178
rect 216232 239086 216260 307770
rect 216220 239080 216272 239086
rect 216220 239022 216272 239028
rect 216324 237794 216352 319534
rect 216416 240582 216444 320146
rect 216496 319864 216548 319870
rect 216496 319806 216548 319812
rect 216404 240576 216456 240582
rect 216404 240518 216456 240524
rect 216312 237788 216364 237794
rect 216312 237730 216364 237736
rect 216128 233640 216180 233646
rect 216128 233582 216180 233588
rect 216140 155582 216168 233582
rect 216324 156913 216352 237730
rect 216508 235346 216536 319806
rect 216600 244274 216628 321642
rect 217874 320240 217930 320249
rect 217874 320175 217930 320184
rect 217784 309800 217836 309806
rect 217784 309742 217836 309748
rect 217416 308440 217468 308446
rect 217416 308382 217468 308388
rect 217232 293140 217284 293146
rect 217232 293082 217284 293088
rect 217138 291816 217194 291825
rect 217138 291751 217194 291760
rect 217152 247722 217180 291751
rect 217140 247716 217192 247722
rect 217140 247658 217192 247664
rect 216600 244246 216720 244274
rect 216692 239834 216720 244246
rect 217138 240408 217194 240417
rect 217138 240343 217194 240352
rect 216680 239828 216732 239834
rect 216680 239770 216732 239776
rect 216588 238128 216640 238134
rect 216588 238070 216640 238076
rect 216600 237862 216628 238070
rect 216588 237856 216640 237862
rect 216588 237798 216640 237804
rect 216586 236736 216642 236745
rect 216586 236671 216642 236680
rect 216600 236065 216628 236671
rect 216586 236056 216642 236065
rect 216586 235991 216642 236000
rect 216692 235414 216720 239770
rect 216680 235408 216732 235414
rect 216680 235350 216732 235356
rect 216496 235340 216548 235346
rect 216496 235282 216548 235288
rect 216310 156904 216366 156913
rect 216310 156839 216366 156848
rect 216128 155576 216180 155582
rect 216128 155518 216180 155524
rect 216036 155508 216088 155514
rect 216036 155450 216088 155456
rect 215944 150408 215996 150414
rect 215944 150350 215996 150356
rect 215298 149968 215354 149977
rect 215298 149903 215354 149912
rect 215944 149796 215996 149802
rect 215944 149738 215996 149744
rect 214564 149116 214616 149122
rect 214564 149058 214616 149064
rect 214194 145888 214250 145897
rect 214194 145823 214250 145832
rect 213932 16546 214512 16574
rect 213184 3800 213236 3806
rect 213184 3742 213236 3748
rect 213104 3454 213408 3482
rect 213380 480 213408 3454
rect 214484 480 214512 16546
rect 214576 3330 214604 149058
rect 215300 148232 215352 148238
rect 215300 148174 215352 148180
rect 215312 146810 215340 148174
rect 215300 146804 215352 146810
rect 215300 146746 215352 146752
rect 215956 144265 215984 149738
rect 217152 149054 217180 240343
rect 217244 216034 217272 293082
rect 217324 291304 217376 291310
rect 217324 291246 217376 291252
rect 217336 246362 217364 291246
rect 217324 246356 217376 246362
rect 217324 246298 217376 246304
rect 217428 241505 217456 308382
rect 217508 307148 217560 307154
rect 217508 307090 217560 307096
rect 217414 241496 217470 241505
rect 217414 241431 217470 241440
rect 217520 241380 217548 307090
rect 217600 307080 217652 307086
rect 217600 307022 217652 307028
rect 217336 241352 217548 241380
rect 217336 239193 217364 241352
rect 217322 239184 217378 239193
rect 217322 239119 217378 239128
rect 217232 216028 217284 216034
rect 217232 215970 217284 215976
rect 217336 154086 217364 239119
rect 217612 238882 217640 307022
rect 217692 292596 217744 292602
rect 217692 292538 217744 292544
rect 217600 238876 217652 238882
rect 217600 238818 217652 238824
rect 217600 236564 217652 236570
rect 217600 236506 217652 236512
rect 217508 236020 217560 236026
rect 217508 235962 217560 235968
rect 217416 233300 217468 233306
rect 217416 233242 217468 233248
rect 217324 154080 217376 154086
rect 217324 154022 217376 154028
rect 217324 152720 217376 152726
rect 217324 152662 217376 152668
rect 217140 149048 217192 149054
rect 217140 148990 217192 148996
rect 216588 146804 216640 146810
rect 216588 146746 216640 146752
rect 215942 144256 215998 144265
rect 215942 144191 215998 144200
rect 215956 3398 215984 144191
rect 215944 3392 215996 3398
rect 215944 3334 215996 3340
rect 214564 3324 214616 3330
rect 214564 3266 214616 3272
rect 215668 3324 215720 3330
rect 215668 3266 215720 3272
rect 215680 480 215708 3266
rect 216600 3194 216628 146746
rect 216678 139904 216734 139913
rect 216678 139839 216734 139848
rect 216692 16574 216720 139839
rect 216692 16546 216904 16574
rect 216588 3188 216640 3194
rect 216588 3130 216640 3136
rect 216876 480 216904 16546
rect 217336 3534 217364 152662
rect 217428 144401 217456 233242
rect 217520 149666 217548 235962
rect 217612 152425 217640 236506
rect 217704 211954 217732 292538
rect 217796 239358 217824 309742
rect 217888 240106 217916 320175
rect 217968 319660 218020 319666
rect 217968 319602 218020 319608
rect 217876 240100 217928 240106
rect 217876 240042 217928 240048
rect 217980 240038 218008 319602
rect 219164 311228 219216 311234
rect 219164 311170 219216 311176
rect 219072 309868 219124 309874
rect 219072 309810 219124 309816
rect 218978 308408 219034 308417
rect 218978 308343 219034 308352
rect 218888 304428 218940 304434
rect 218888 304370 218940 304376
rect 218796 297356 218848 297362
rect 218796 297298 218848 297304
rect 218520 292732 218572 292738
rect 218520 292674 218572 292680
rect 217968 240032 218020 240038
rect 217968 239974 218020 239980
rect 217784 239352 217836 239358
rect 217784 239294 217836 239300
rect 217796 233646 217824 239294
rect 217784 233640 217836 233646
rect 217784 233582 217836 233588
rect 217784 230308 217836 230314
rect 217784 230250 217836 230256
rect 217692 211948 217744 211954
rect 217692 211890 217744 211896
rect 217796 152726 217824 230250
rect 218532 209681 218560 292674
rect 218702 292224 218758 292233
rect 218702 292159 218758 292168
rect 218612 291984 218664 291990
rect 218612 291926 218664 291932
rect 218624 244934 218652 291926
rect 218612 244928 218664 244934
rect 218612 244870 218664 244876
rect 218716 243574 218744 292159
rect 218704 243568 218756 243574
rect 218704 243510 218756 243516
rect 218808 239698 218836 297298
rect 218900 240854 218928 304370
rect 218888 240848 218940 240854
rect 218992 240825 219020 308343
rect 219084 241126 219112 309810
rect 219072 241120 219124 241126
rect 219072 241062 219124 241068
rect 218888 240790 218940 240796
rect 218978 240816 219034 240825
rect 218796 239692 218848 239698
rect 218796 239634 218848 239640
rect 218900 239578 218928 240790
rect 218978 240751 219034 240760
rect 218992 240417 219020 240751
rect 218978 240408 219034 240417
rect 218978 240343 219034 240352
rect 219084 240242 219112 241062
rect 219072 240236 219124 240242
rect 219072 240178 219124 240184
rect 218980 239692 219032 239698
rect 218980 239634 219032 239640
rect 218716 239550 218928 239578
rect 218518 209672 218574 209681
rect 218518 209607 218574 209616
rect 218532 209137 218560 209607
rect 218518 209128 218574 209137
rect 218518 209063 218574 209072
rect 217784 152720 217836 152726
rect 217784 152662 217836 152668
rect 217598 152416 217654 152425
rect 217598 152351 217654 152360
rect 218716 149870 218744 239550
rect 218992 238202 219020 239634
rect 218980 238196 219032 238202
rect 218980 238138 219032 238144
rect 218794 236872 218850 236881
rect 218794 236807 218850 236816
rect 218704 149864 218756 149870
rect 218704 149806 218756 149812
rect 217508 149660 217560 149666
rect 217508 149602 217560 149608
rect 218058 146024 218114 146033
rect 218058 145959 218114 145968
rect 218072 145625 218100 145959
rect 218808 145625 218836 236807
rect 219176 233102 219204 311170
rect 219256 292664 219308 292670
rect 219256 292606 219308 292612
rect 219164 233096 219216 233102
rect 219164 233038 219216 233044
rect 219268 209778 219296 292606
rect 219360 285190 219388 321671
rect 219716 315308 219768 315314
rect 219716 315250 219768 315256
rect 219348 285184 219400 285190
rect 219348 285126 219400 285132
rect 219346 241360 219402 241369
rect 219346 241295 219402 241304
rect 219360 240242 219388 241295
rect 219532 240644 219584 240650
rect 219532 240586 219584 240592
rect 219348 240236 219400 240242
rect 219348 240178 219400 240184
rect 219544 240106 219572 240586
rect 219532 240100 219584 240106
rect 219532 240042 219584 240048
rect 219544 233374 219572 240042
rect 219532 233368 219584 233374
rect 219532 233310 219584 233316
rect 219728 233034 219756 315250
rect 219808 308576 219860 308582
rect 219808 308518 219860 308524
rect 219820 233238 219848 308518
rect 219912 290766 219940 372574
rect 220174 307048 220230 307057
rect 220174 306983 220230 306992
rect 219992 292324 220044 292330
rect 219992 292266 220044 292272
rect 219900 290760 219952 290766
rect 219900 290702 219952 290708
rect 219900 290284 219952 290290
rect 219900 290226 219952 290232
rect 219808 233232 219860 233238
rect 219808 233174 219860 233180
rect 219716 233028 219768 233034
rect 219716 232970 219768 232976
rect 219912 212498 219940 290226
rect 220004 280838 220032 292266
rect 220084 291576 220136 291582
rect 220084 291518 220136 291524
rect 219992 280832 220044 280838
rect 219992 280774 220044 280780
rect 219992 241460 220044 241466
rect 219992 241402 220044 241408
rect 220004 236570 220032 241402
rect 220096 239630 220124 291518
rect 220188 241466 220216 306983
rect 220372 293282 220400 373186
rect 220360 293276 220412 293282
rect 220360 293218 220412 293224
rect 220266 291952 220322 291961
rect 220266 291887 220322 291896
rect 220176 241460 220228 241466
rect 220176 241402 220228 241408
rect 220280 241346 220308 291887
rect 220464 291854 220492 373215
rect 220636 304564 220688 304570
rect 220636 304506 220688 304512
rect 220452 291848 220504 291854
rect 220452 291790 220504 291796
rect 220360 291644 220412 291650
rect 220360 291586 220412 291592
rect 220372 273970 220400 291586
rect 220544 289808 220596 289814
rect 220544 289750 220596 289756
rect 220360 273964 220412 273970
rect 220360 273906 220412 273912
rect 220188 241318 220308 241346
rect 220188 240786 220216 241318
rect 220358 240952 220414 240961
rect 220268 240916 220320 240922
rect 220358 240887 220414 240896
rect 220268 240858 220320 240864
rect 220176 240780 220228 240786
rect 220176 240722 220228 240728
rect 220280 240134 220308 240858
rect 220372 240786 220400 240887
rect 220360 240780 220412 240786
rect 220360 240722 220412 240728
rect 220188 240106 220308 240134
rect 220084 239624 220136 239630
rect 220084 239566 220136 239572
rect 220188 239476 220216 240106
rect 220556 239494 220584 289750
rect 220648 284322 220676 304506
rect 220740 291938 220768 375362
rect 222106 374096 222162 374105
rect 222106 374031 222162 374040
rect 222014 369880 222070 369889
rect 222014 369815 222070 369824
rect 221646 305688 221702 305697
rect 221646 305623 221702 305632
rect 220740 291910 220860 291938
rect 220832 291854 220860 291910
rect 220728 291848 220780 291854
rect 220728 291790 220780 291796
rect 220820 291848 220872 291854
rect 220820 291790 220872 291796
rect 220740 291689 220768 291790
rect 221004 291780 221056 291786
rect 221004 291722 221056 291728
rect 220726 291680 220782 291689
rect 220726 291615 220782 291624
rect 220820 291508 220872 291514
rect 220820 291450 220872 291456
rect 220728 290352 220780 290358
rect 220726 290320 220728 290329
rect 220780 290320 220782 290329
rect 220726 290255 220782 290264
rect 220832 285122 220860 291450
rect 220912 291440 220964 291446
rect 220912 291382 220964 291388
rect 220924 286414 220952 291382
rect 220912 286408 220964 286414
rect 220912 286350 220964 286356
rect 220912 286272 220964 286278
rect 221016 286226 221044 291722
rect 221280 291372 221332 291378
rect 221280 291314 221332 291320
rect 221292 287054 221320 291314
rect 221372 291236 221424 291242
rect 221372 291178 221424 291184
rect 220964 286220 221044 286226
rect 220912 286214 221044 286220
rect 220924 286198 221044 286214
rect 221108 287026 221320 287054
rect 220912 285184 220964 285190
rect 220910 285152 220912 285161
rect 220964 285152 220966 285161
rect 220820 285116 220872 285122
rect 220910 285087 220966 285096
rect 220820 285058 220872 285064
rect 220648 284294 220860 284322
rect 220832 277394 220860 284294
rect 221108 283642 221136 287026
rect 220924 283626 221136 283642
rect 220912 283620 221136 283626
rect 220964 283614 221136 283620
rect 220912 283562 220964 283568
rect 221384 279562 221412 291178
rect 221554 285152 221610 285161
rect 221554 285087 221610 285096
rect 220924 279534 221412 279562
rect 220924 279478 220952 279534
rect 220912 279472 220964 279478
rect 220912 279414 220964 279420
rect 220832 277366 221504 277394
rect 220910 276720 220966 276729
rect 220910 276655 220912 276664
rect 220964 276655 220966 276664
rect 220912 276626 220964 276632
rect 221188 241664 221240 241670
rect 221188 241606 221240 241612
rect 220820 241120 220872 241126
rect 220820 241062 220872 241068
rect 220832 240689 220860 241062
rect 220818 240680 220874 240689
rect 220818 240615 220874 240624
rect 221094 240136 221150 240145
rect 221094 240071 221150 240080
rect 221108 239630 221136 240071
rect 221200 239748 221228 241606
rect 221372 241460 221424 241466
rect 221372 241402 221424 241408
rect 221384 241330 221412 241402
rect 221372 241324 221424 241330
rect 221372 241266 221424 241272
rect 221278 240952 221334 240961
rect 221278 240887 221334 240896
rect 221292 239902 221320 240887
rect 221280 239896 221332 239902
rect 221280 239838 221332 239844
rect 221200 239720 221412 239748
rect 221096 239624 221148 239630
rect 221096 239566 221148 239572
rect 221384 239494 221412 239720
rect 220096 239448 220216 239476
rect 220544 239488 220596 239494
rect 219992 236564 220044 236570
rect 219992 236506 220044 236512
rect 219992 234184 220044 234190
rect 219992 234126 220044 234132
rect 219900 212492 219952 212498
rect 219900 212434 219952 212440
rect 219256 209772 219308 209778
rect 219256 209714 219308 209720
rect 219268 209098 219296 209714
rect 219256 209092 219308 209098
rect 219256 209034 219308 209040
rect 220004 155689 220032 234126
rect 219990 155680 220046 155689
rect 219990 155615 220046 155624
rect 220096 152454 220124 239448
rect 220544 239430 220596 239436
rect 221280 239488 221332 239494
rect 221280 239430 221332 239436
rect 221372 239488 221424 239494
rect 221372 239430 221424 239436
rect 220268 238944 220320 238950
rect 220268 238886 220320 238892
rect 220176 235340 220228 235346
rect 220176 235282 220228 235288
rect 220084 152448 220136 152454
rect 220084 152390 220136 152396
rect 220084 149048 220136 149054
rect 220084 148990 220136 148996
rect 218058 145616 218114 145625
rect 218058 145551 218114 145560
rect 218794 145616 218850 145625
rect 218794 145551 218850 145560
rect 217414 144392 217470 144401
rect 217414 144327 217470 144336
rect 219440 137284 219492 137290
rect 219440 137226 219492 137232
rect 219452 16574 219480 137226
rect 219452 16546 220032 16574
rect 217324 3528 217376 3534
rect 217324 3470 217376 3476
rect 218060 3460 218112 3466
rect 218060 3402 218112 3408
rect 218072 480 218100 3402
rect 219256 3188 219308 3194
rect 219256 3130 219308 3136
rect 219268 480 219296 3130
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220096 3670 220124 148990
rect 220188 143138 220216 235282
rect 220280 156670 220308 238886
rect 220728 238876 220780 238882
rect 220728 238818 220780 238824
rect 220360 238808 220412 238814
rect 220360 238750 220412 238756
rect 220372 156738 220400 238750
rect 220740 237153 220768 238818
rect 221292 238241 221320 239430
rect 221278 238232 221334 238241
rect 221278 238167 221334 238176
rect 221476 237998 221504 277366
rect 221568 239902 221596 285087
rect 221556 239896 221608 239902
rect 221556 239838 221608 239844
rect 221464 237992 221516 237998
rect 221464 237934 221516 237940
rect 220726 237144 220782 237153
rect 220726 237079 220782 237088
rect 220450 235240 220506 235249
rect 220450 235175 220506 235184
rect 220360 156732 220412 156738
rect 220360 156674 220412 156680
rect 220268 156664 220320 156670
rect 220268 156606 220320 156612
rect 220464 155281 220492 235175
rect 220450 155272 220506 155281
rect 220450 155207 220506 155216
rect 220740 154018 220768 237079
rect 220728 154012 220780 154018
rect 220728 153954 220780 153960
rect 220176 143132 220228 143138
rect 220176 143074 220228 143080
rect 221476 142769 221504 237934
rect 221660 237318 221688 305623
rect 221924 298852 221976 298858
rect 221924 298794 221976 298800
rect 221740 290420 221792 290426
rect 221740 290362 221792 290368
rect 221648 237312 221700 237318
rect 221648 237254 221700 237260
rect 221556 236768 221608 236774
rect 221556 236710 221608 236716
rect 221568 157962 221596 236710
rect 221646 227080 221702 227089
rect 221646 227015 221702 227024
rect 221556 157956 221608 157962
rect 221556 157898 221608 157904
rect 221462 142760 221518 142769
rect 221462 142695 221518 142704
rect 221660 142633 221688 227015
rect 221752 212022 221780 290362
rect 221936 290358 221964 298794
rect 222028 294642 222056 369815
rect 222016 294636 222068 294642
rect 222016 294578 222068 294584
rect 222028 294030 222056 294578
rect 222016 294024 222068 294030
rect 222016 293966 222068 293972
rect 222120 291990 222148 374031
rect 226984 373312 227036 373318
rect 226984 373254 227036 373260
rect 224224 361616 224276 361622
rect 224224 361558 224276 361564
rect 222200 314084 222252 314090
rect 222200 314026 222252 314032
rect 222108 291984 222160 291990
rect 222108 291926 222160 291932
rect 222016 291712 222068 291718
rect 222016 291654 222068 291660
rect 221924 290352 221976 290358
rect 221924 290294 221976 290300
rect 221830 290184 221886 290193
rect 221830 290119 221886 290128
rect 221844 212158 221872 290119
rect 221936 212294 221964 290294
rect 222028 276729 222056 291654
rect 222014 276720 222070 276729
rect 222014 276655 222070 276664
rect 222016 240712 222068 240718
rect 222016 240654 222068 240660
rect 222028 240145 222056 240654
rect 222014 240136 222070 240145
rect 222014 240071 222070 240080
rect 222108 240032 222160 240038
rect 222108 239974 222160 239980
rect 222120 239476 222148 239974
rect 222212 239698 222240 314026
rect 222292 295996 222344 296002
rect 222292 295938 222344 295944
rect 222304 241602 222332 295938
rect 224236 292913 224264 361558
rect 225602 360904 225658 360913
rect 225602 360839 225658 360848
rect 224316 301504 224368 301510
rect 224316 301446 224368 301452
rect 224222 292904 224278 292913
rect 224222 292839 224278 292848
rect 224328 290170 224356 301446
rect 225616 296714 225644 360839
rect 225694 359408 225750 359417
rect 225694 359343 225750 359352
rect 225524 296686 225644 296714
rect 225052 294024 225104 294030
rect 225052 293966 225104 293972
rect 224682 292904 224738 292913
rect 224682 292839 224738 292848
rect 224590 291952 224646 291961
rect 224590 291887 224646 291896
rect 224604 291689 224632 291887
rect 224406 291680 224462 291689
rect 224590 291680 224646 291689
rect 224462 291638 224540 291666
rect 224406 291615 224462 291624
rect 224236 290142 224356 290170
rect 224236 289898 224264 290142
rect 223592 289870 224264 289898
rect 223592 289814 223620 289870
rect 223580 289808 223632 289814
rect 224512 289762 224540 291638
rect 224590 291615 224646 291624
rect 224696 289884 224724 292839
rect 225064 289884 225092 293966
rect 225524 291281 225552 296686
rect 225708 294506 225736 359343
rect 225786 330440 225842 330449
rect 225786 330375 225842 330384
rect 225696 294500 225748 294506
rect 225696 294442 225748 294448
rect 225708 294030 225736 294442
rect 225696 294024 225748 294030
rect 225696 293966 225748 293972
rect 225800 292641 225828 330375
rect 225878 318744 225934 318753
rect 225878 318679 225934 318688
rect 225892 298081 225920 318679
rect 226064 309936 226116 309942
rect 226064 309878 226116 309884
rect 225878 298072 225934 298081
rect 225878 298007 225934 298016
rect 225972 294024 226024 294030
rect 225972 293966 226024 293972
rect 225786 292632 225842 292641
rect 225786 292567 225842 292576
rect 225510 291272 225566 291281
rect 225510 291207 225566 291216
rect 225800 290170 225828 292567
rect 225708 290142 225828 290170
rect 225708 289898 225736 290142
rect 225446 289870 225736 289898
rect 225984 289762 226012 293966
rect 223580 289750 223632 289756
rect 224342 289734 224540 289762
rect 225814 289734 226012 289762
rect 226076 289649 226104 309878
rect 226524 293276 226576 293282
rect 226524 293218 226576 293224
rect 226154 291272 226210 291281
rect 226154 291207 226210 291216
rect 226168 289884 226196 291207
rect 226536 289884 226564 293218
rect 226996 292738 227024 373254
rect 231768 370660 231820 370666
rect 231768 370602 231820 370608
rect 228364 370524 228416 370530
rect 228364 370466 228416 370472
rect 227074 369200 227130 369209
rect 227074 369135 227130 369144
rect 227088 294574 227116 369135
rect 227996 294704 228048 294710
rect 227996 294646 228048 294652
rect 227076 294568 227128 294574
rect 227076 294510 227128 294516
rect 226984 292732 227036 292738
rect 226984 292674 227036 292680
rect 226996 292534 227024 292674
rect 226984 292528 227036 292534
rect 226984 292470 227036 292476
rect 227088 289898 227116 294510
rect 227720 292664 227772 292670
rect 227720 292606 227772 292612
rect 227732 292466 227760 292606
rect 227720 292460 227772 292466
rect 227720 292402 227772 292408
rect 227720 292120 227772 292126
rect 227720 292062 227772 292068
rect 227260 291984 227312 291990
rect 227260 291926 227312 291932
rect 226918 289870 227116 289898
rect 227272 289884 227300 291926
rect 227732 290766 227760 292062
rect 227720 290760 227772 290766
rect 227720 290702 227772 290708
rect 227626 290320 227682 290329
rect 227626 290255 227682 290264
rect 227640 289884 227668 290255
rect 228008 289884 228036 294646
rect 228376 292466 228404 370466
rect 231124 369164 231176 369170
rect 231124 369106 231176 369112
rect 229742 368928 229798 368937
rect 229742 368863 229798 368872
rect 228456 368552 228508 368558
rect 228456 368494 228508 368500
rect 228468 294710 228496 368494
rect 228546 322280 228602 322289
rect 228546 322215 228602 322224
rect 228456 294704 228508 294710
rect 228456 294646 228508 294652
rect 228364 292460 228416 292466
rect 228364 292402 228416 292408
rect 228560 291310 228588 322215
rect 229756 296714 229784 368863
rect 229836 354000 229888 354006
rect 229836 353942 229888 353948
rect 229388 296686 229784 296714
rect 229388 294234 229416 296686
rect 229848 294438 229876 353942
rect 229926 323640 229982 323649
rect 229926 323575 229982 323584
rect 229836 294432 229888 294438
rect 229836 294374 229888 294380
rect 229100 294228 229152 294234
rect 229100 294170 229152 294176
rect 229376 294228 229428 294234
rect 229376 294170 229428 294176
rect 228732 292528 228784 292534
rect 228732 292470 228784 292476
rect 228548 291304 228600 291310
rect 228548 291246 228600 291252
rect 228560 289898 228588 291246
rect 228390 289870 228588 289898
rect 228744 289884 228772 292470
rect 229112 289884 229140 294170
rect 229836 292460 229888 292466
rect 229836 292402 229888 292408
rect 229466 291816 229522 291825
rect 229466 291751 229522 291760
rect 229480 289884 229508 291751
rect 229848 289884 229876 292402
rect 229940 291825 229968 323575
rect 230202 318608 230258 318617
rect 230202 318543 230258 318552
rect 230216 294681 230244 318543
rect 230756 300076 230808 300082
rect 230756 300018 230808 300024
rect 230572 296200 230624 296206
rect 230572 296142 230624 296148
rect 230584 295934 230612 296142
rect 230572 295928 230624 295934
rect 230572 295870 230624 295876
rect 230202 294672 230258 294681
rect 230202 294607 230258 294616
rect 230204 294432 230256 294438
rect 230204 294374 230256 294380
rect 229926 291816 229982 291825
rect 229926 291751 229982 291760
rect 230216 289884 230244 294374
rect 230584 289884 230612 295870
rect 230768 290018 230796 300018
rect 231136 292806 231164 369106
rect 231216 324964 231268 324970
rect 231216 324906 231268 324912
rect 231228 296206 231256 324906
rect 231780 300082 231808 370602
rect 231768 300076 231820 300082
rect 231768 300018 231820 300024
rect 231780 299538 231808 300018
rect 231768 299532 231820 299538
rect 231768 299474 231820 299480
rect 232516 296714 232544 375770
rect 235264 375760 235316 375766
rect 235264 375702 235316 375708
rect 234620 370864 234672 370870
rect 234620 370806 234672 370812
rect 233148 370728 233200 370734
rect 233148 370670 233200 370676
rect 233160 298790 233188 370670
rect 233884 369232 233936 369238
rect 233884 369174 233936 369180
rect 233148 298784 233200 298790
rect 233148 298726 233200 298732
rect 232424 296686 232544 296714
rect 231216 296200 231268 296206
rect 231216 296142 231268 296148
rect 231306 294672 231362 294681
rect 231306 294607 231362 294616
rect 231320 294409 231348 294607
rect 231306 294400 231362 294409
rect 231306 294335 231362 294344
rect 232424 294302 232452 296686
rect 232412 294296 232464 294302
rect 232412 294238 232464 294244
rect 231952 293344 232004 293350
rect 231952 293286 232004 293292
rect 231964 293078 231992 293286
rect 232044 293208 232096 293214
rect 232044 293150 232096 293156
rect 232056 293078 232084 293150
rect 231952 293072 232004 293078
rect 231952 293014 232004 293020
rect 232044 293072 232096 293078
rect 232044 293014 232096 293020
rect 231124 292800 231176 292806
rect 231124 292742 231176 292748
rect 231308 292800 231360 292806
rect 231308 292742 231360 292748
rect 230756 290012 230808 290018
rect 230756 289954 230808 289960
rect 230768 289898 230796 289954
rect 230768 289870 230966 289898
rect 231320 289884 231348 292742
rect 231676 291848 231728 291854
rect 231676 291790 231728 291796
rect 231688 289884 231716 291790
rect 232056 289884 232084 293014
rect 232424 289884 232452 294238
rect 233160 293078 233188 298726
rect 233700 298104 233752 298110
rect 233700 298046 233752 298052
rect 233712 297090 233740 298046
rect 233700 297084 233752 297090
rect 233700 297026 233752 297032
rect 233516 295520 233568 295526
rect 233516 295462 233568 295468
rect 233148 293072 233200 293078
rect 233148 293014 233200 293020
rect 232780 292868 232832 292874
rect 232780 292810 232832 292816
rect 232792 289884 232820 292810
rect 233148 292120 233200 292126
rect 233148 292062 233200 292068
rect 233160 289884 233188 292062
rect 233528 289884 233556 295462
rect 233712 289898 233740 297026
rect 233896 295526 233924 369174
rect 233976 326392 234028 326398
rect 233976 326334 234028 326340
rect 233988 298110 234016 326334
rect 233976 298104 234028 298110
rect 233976 298046 234028 298052
rect 233884 295520 233936 295526
rect 233884 295462 233936 295468
rect 234252 294772 234304 294778
rect 234252 294714 234304 294720
rect 234264 294166 234292 294714
rect 234252 294160 234304 294166
rect 234252 294102 234304 294108
rect 233712 289870 233910 289898
rect 234264 289884 234292 294102
rect 234632 290170 234660 370806
rect 235276 296714 235304 375702
rect 237380 375692 237432 375698
rect 237380 375634 237432 375640
rect 236644 375488 236696 375494
rect 236644 375430 236696 375436
rect 235356 370184 235408 370190
rect 235356 370126 235408 370132
rect 235368 296954 235396 370126
rect 236656 297430 236684 375430
rect 237392 306374 237420 375634
rect 240140 375624 240192 375630
rect 240140 375566 240192 375572
rect 238116 372768 238168 372774
rect 238116 372710 238168 372716
rect 238024 372224 238076 372230
rect 238024 372166 238076 372172
rect 237392 306346 237788 306374
rect 236644 297424 236696 297430
rect 236644 297366 236696 297372
rect 235356 296948 235408 296954
rect 235356 296890 235408 296896
rect 234908 296686 235304 296714
rect 235368 296714 235396 296890
rect 236656 296714 236684 297366
rect 235368 296686 235488 296714
rect 236656 296686 237052 296714
rect 234908 295798 234936 296686
rect 234896 295792 234948 295798
rect 234896 295734 234948 295740
rect 234540 290142 234660 290170
rect 226062 289640 226118 289649
rect 226062 289575 226118 289584
rect 234540 289406 234568 290142
rect 234908 289898 234936 295734
rect 234988 295520 235040 295526
rect 234988 295462 235040 295468
rect 235000 291922 235028 295462
rect 235356 293276 235408 293282
rect 235356 293218 235408 293224
rect 235368 292602 235396 293218
rect 235356 292596 235408 292602
rect 235356 292538 235408 292544
rect 234988 291916 235040 291922
rect 234988 291858 235040 291864
rect 234646 289870 234936 289898
rect 235000 289884 235028 291858
rect 235368 289884 235396 292538
rect 235460 291242 235488 296686
rect 236460 293344 236512 293350
rect 236460 293286 236512 293292
rect 235448 291236 235500 291242
rect 235448 291178 235500 291184
rect 236092 291236 236144 291242
rect 236092 291178 236144 291184
rect 236104 289884 236132 291178
rect 236472 289884 236500 293286
rect 236828 291848 236880 291854
rect 236828 291790 236880 291796
rect 236840 290154 236868 291790
rect 236828 290148 236880 290154
rect 236828 290090 236880 290096
rect 236840 289884 236868 290090
rect 237024 289898 237052 296686
rect 237380 293684 237432 293690
rect 237380 293626 237432 293632
rect 237392 292262 237420 293626
rect 237472 293412 237524 293418
rect 237472 293354 237524 293360
rect 237484 292942 237512 293354
rect 237472 292936 237524 292942
rect 237472 292878 237524 292884
rect 237380 292256 237432 292262
rect 237380 292198 237432 292204
rect 237484 289898 237512 292878
rect 237760 289898 237788 306346
rect 238036 292874 238064 372166
rect 238128 297226 238156 372710
rect 239404 372292 239456 372298
rect 239404 372234 239456 372240
rect 238116 297220 238168 297226
rect 238116 297162 238168 297168
rect 238024 292868 238076 292874
rect 238024 292810 238076 292816
rect 238128 291242 238156 297162
rect 239036 295588 239088 295594
rect 239036 295530 239088 295536
rect 238392 294636 238444 294642
rect 238392 294578 238444 294584
rect 238404 293622 238432 294578
rect 238392 293616 238444 293622
rect 238392 293558 238444 293564
rect 238404 292574 238432 293558
rect 238404 292546 238524 292574
rect 238300 292256 238352 292262
rect 238300 292198 238352 292204
rect 238116 291236 238168 291242
rect 238116 291178 238168 291184
rect 237024 289870 237222 289898
rect 237484 289870 237590 289898
rect 237760 289870 237880 289898
rect 238312 289884 238340 292198
rect 238496 289898 238524 292546
rect 238496 289870 238694 289898
rect 239048 289884 239076 295530
rect 239416 295526 239444 372234
rect 240152 306374 240180 375566
rect 242164 370116 242216 370122
rect 242164 370058 242216 370064
rect 240152 306346 240456 306374
rect 240048 296132 240100 296138
rect 240048 296074 240100 296080
rect 240060 295594 240088 296074
rect 240048 295588 240100 295594
rect 240048 295530 240100 295536
rect 239404 295520 239456 295526
rect 239404 295462 239456 295468
rect 240048 294704 240100 294710
rect 240048 294646 240100 294652
rect 240060 293010 240088 294646
rect 240048 293004 240100 293010
rect 240048 292946 240100 292952
rect 239404 291236 239456 291242
rect 239404 291178 239456 291184
rect 239416 289884 239444 291178
rect 240060 289898 240088 292946
rect 240428 292574 240456 306346
rect 242176 295662 242204 370058
rect 243268 368620 243320 368626
rect 243268 368562 243320 368568
rect 242440 318164 242492 318170
rect 242440 318106 242492 318112
rect 242452 314090 242480 318106
rect 242440 314084 242492 314090
rect 242440 314026 242492 314032
rect 242808 296064 242860 296070
rect 242808 296006 242860 296012
rect 242164 295656 242216 295662
rect 242164 295598 242216 295604
rect 241980 295452 242032 295458
rect 241980 295394 242032 295400
rect 241612 294364 241664 294370
rect 241612 294306 241664 294312
rect 240428 292546 240548 292574
rect 240140 290760 240192 290766
rect 240140 290702 240192 290708
rect 240152 290494 240180 290702
rect 240140 290488 240192 290494
rect 240140 290430 240192 290436
rect 239798 289870 240088 289898
rect 240152 289884 240180 290430
rect 240520 290426 240548 292546
rect 241624 292398 241652 294306
rect 241888 293140 241940 293146
rect 241888 293082 241940 293088
rect 241900 292534 241928 293082
rect 241888 292528 241940 292534
rect 241888 292470 241940 292476
rect 241612 292392 241664 292398
rect 241612 292334 241664 292340
rect 240876 291304 240928 291310
rect 240876 291246 240928 291252
rect 240508 290420 240560 290426
rect 240508 290362 240560 290368
rect 240520 289884 240548 290362
rect 240888 289884 240916 291246
rect 241624 289884 241652 292334
rect 241900 291310 241928 292470
rect 241888 291304 241940 291310
rect 241888 291246 241940 291252
rect 241992 289884 242020 295394
rect 242176 289898 242204 295598
rect 242820 295458 242848 296006
rect 242808 295452 242860 295458
rect 242808 295394 242860 295400
rect 243084 295316 243136 295322
rect 243084 295258 243136 295264
rect 242716 291984 242768 291990
rect 242716 291926 242768 291932
rect 242728 291242 242756 291926
rect 242716 291236 242768 291242
rect 242716 291178 242768 291184
rect 242176 289870 242374 289898
rect 242728 289884 242756 291178
rect 243096 289884 243124 295258
rect 243280 289898 243308 368562
rect 243556 306374 243584 379578
rect 244924 372836 244976 372842
rect 244924 372778 244976 372784
rect 244280 318300 244332 318306
rect 244280 318242 244332 318248
rect 244292 317121 244320 318242
rect 244278 317112 244334 317121
rect 244278 317047 244334 317056
rect 243556 306346 243676 306374
rect 243360 295860 243412 295866
rect 243360 295802 243412 295808
rect 243372 295322 243400 295802
rect 243360 295316 243412 295322
rect 243360 295258 243412 295264
rect 243648 291786 243676 306346
rect 244556 296812 244608 296818
rect 244556 296754 244608 296760
rect 243636 291780 243688 291786
rect 243636 291722 243688 291728
rect 243648 289898 243676 291722
rect 244188 291712 244240 291718
rect 244240 291660 244320 291666
rect 244188 291654 244320 291660
rect 244200 291638 244320 291654
rect 244292 291242 244320 291638
rect 244280 291236 244332 291242
rect 244280 291178 244332 291184
rect 244188 290488 244240 290494
rect 244188 290430 244240 290436
rect 244200 289898 244228 290430
rect 243280 289882 243478 289898
rect 243268 289876 243478 289882
rect 235552 289462 235750 289490
rect 235552 289406 235580 289462
rect 234528 289400 234580 289406
rect 234528 289342 234580 289348
rect 235540 289400 235592 289406
rect 237852 289388 237880 289870
rect 243320 289870 243478 289876
rect 243648 289870 243846 289898
rect 244016 289884 244228 289898
rect 244568 289884 244596 296754
rect 244936 291242 244964 372778
rect 245016 369912 245068 369918
rect 245016 369854 245068 369860
rect 245028 296818 245056 369854
rect 245660 368688 245712 368694
rect 245660 368630 245712 368636
rect 245016 296812 245068 296818
rect 245016 296754 245068 296760
rect 245292 292052 245344 292058
rect 245292 291994 245344 292000
rect 244924 291236 244976 291242
rect 244924 291178 244976 291184
rect 244936 289884 244964 291178
rect 245304 289898 245332 291994
rect 245672 289898 245700 368630
rect 246316 292194 246344 380938
rect 250536 379908 250588 379914
rect 250536 379850 250588 379856
rect 246396 379772 246448 379778
rect 246396 379714 246448 379720
rect 246408 297022 246436 379714
rect 250444 376916 250496 376922
rect 250444 376858 250496 376864
rect 248418 367704 248474 367713
rect 248418 367639 248474 367648
rect 247682 363624 247738 363633
rect 247682 363559 247738 363568
rect 247040 318232 247092 318238
rect 247040 318174 247092 318180
rect 246948 315444 247000 315450
rect 246948 315386 247000 315392
rect 246396 297016 246448 297022
rect 246396 296958 246448 296964
rect 246408 292574 246436 296958
rect 246408 292546 246620 292574
rect 246304 292188 246356 292194
rect 246304 292130 246356 292136
rect 246316 289898 246344 292130
rect 245212 289884 245332 289898
rect 245488 289884 245700 289898
rect 244016 289870 244214 289884
rect 245212 289870 245318 289884
rect 245488 289870 245686 289884
rect 246054 289870 246344 289898
rect 246592 289898 246620 292546
rect 246592 289870 246790 289898
rect 243268 289818 243320 289824
rect 244016 289406 244044 289870
rect 245212 289474 245240 289870
rect 245200 289468 245252 289474
rect 245200 289410 245252 289416
rect 245488 289406 245516 289870
rect 246394 289640 246450 289649
rect 246394 289575 246450 289584
rect 246960 289490 246988 315386
rect 247052 315217 247080 318174
rect 247038 315208 247094 315217
rect 247038 315143 247094 315152
rect 247040 294092 247092 294098
rect 247040 294034 247092 294040
rect 247052 292466 247080 294034
rect 247696 292574 247724 363559
rect 247774 352608 247830 352617
rect 247774 352543 247830 352552
rect 247420 292546 247724 292574
rect 247040 292460 247092 292466
rect 247040 292402 247092 292408
rect 247420 291582 247448 292546
rect 247500 292460 247552 292466
rect 247500 292402 247552 292408
rect 247408 291576 247460 291582
rect 247408 291518 247460 291524
rect 247420 289898 247448 291518
rect 247158 289870 247448 289898
rect 247512 289884 247540 292402
rect 247788 291650 247816 352543
rect 248144 314696 248196 314702
rect 248144 314638 248196 314644
rect 248052 314084 248104 314090
rect 248052 314026 248104 314032
rect 247868 291916 247920 291922
rect 247868 291858 247920 291864
rect 247776 291644 247828 291650
rect 247776 291586 247828 291592
rect 247788 291242 247816 291586
rect 247776 291236 247828 291242
rect 247776 291178 247828 291184
rect 247682 289912 247738 289921
rect 247880 289898 247908 291858
rect 247738 289884 247908 289898
rect 247738 289870 247894 289884
rect 247682 289847 247738 289856
rect 248064 289513 248092 314026
rect 248156 289649 248184 314638
rect 248432 306374 248460 367639
rect 249064 363656 249116 363662
rect 249064 363598 249116 363604
rect 248432 306346 248644 306374
rect 248616 302234 248644 306346
rect 248616 302206 248828 302234
rect 248604 297220 248656 297226
rect 248604 297162 248656 297168
rect 248616 296886 248644 297162
rect 248604 296880 248656 296886
rect 248604 296822 248656 296828
rect 248236 291236 248288 291242
rect 248236 291178 248288 291184
rect 248328 291236 248380 291242
rect 248328 291178 248380 291184
rect 248248 289884 248276 291178
rect 248340 290737 248368 291178
rect 248326 290728 248382 290737
rect 248326 290663 248382 290672
rect 248616 289884 248644 296822
rect 248800 289762 248828 302206
rect 249076 297226 249104 363598
rect 249156 321156 249208 321162
rect 249156 321098 249208 321104
rect 249064 297220 249116 297226
rect 249064 297162 249116 297168
rect 249168 291689 249196 321098
rect 249340 292256 249392 292262
rect 249340 292198 249392 292204
rect 249352 292126 249380 292198
rect 249340 292120 249392 292126
rect 249340 292062 249392 292068
rect 250456 291990 250484 376858
rect 250548 295390 250576 379850
rect 251822 369064 251878 369073
rect 251822 368999 251878 369008
rect 250626 366344 250682 366353
rect 250626 366279 250682 366288
rect 250536 295384 250588 295390
rect 250536 295326 250588 295332
rect 250444 291984 250496 291990
rect 250444 291926 250496 291932
rect 249154 291680 249210 291689
rect 249154 291615 249210 291624
rect 249168 289898 249196 291615
rect 249706 290728 249762 290737
rect 249706 290663 249762 290672
rect 249720 290193 249748 290663
rect 250548 290306 250576 295326
rect 250640 291553 250668 366279
rect 251178 292088 251234 292097
rect 251178 292023 251234 292032
rect 250810 291952 250866 291961
rect 250810 291887 250866 291896
rect 250626 291544 250682 291553
rect 250626 291479 250682 291488
rect 250364 290278 250576 290306
rect 249706 290184 249762 290193
rect 249706 290119 249762 290128
rect 249168 289870 249366 289898
rect 249720 289884 249748 290119
rect 250364 289898 250392 290278
rect 250640 289898 250668 291479
rect 250824 291242 250852 291887
rect 250812 291236 250864 291242
rect 250812 291178 250864 291184
rect 250102 289870 250392 289898
rect 250470 289870 250668 289898
rect 250824 289884 250852 291178
rect 251192 290329 251220 292023
rect 251546 291408 251602 291417
rect 251546 291343 251602 291352
rect 251178 290320 251234 290329
rect 251178 290255 251234 290264
rect 251192 289884 251220 290255
rect 251560 289884 251588 291343
rect 251836 290329 251864 368999
rect 251914 361040 251970 361049
rect 251914 360975 251970 360984
rect 251928 291417 251956 360975
rect 252468 312656 252520 312662
rect 252468 312598 252520 312604
rect 251914 291408 251970 291417
rect 251914 291343 251970 291352
rect 251914 290456 251970 290465
rect 251914 290391 251970 290400
rect 251822 290320 251878 290329
rect 251822 290255 251878 290264
rect 251730 290048 251786 290057
rect 251730 289983 251786 289992
rect 251744 289898 251772 289983
rect 251928 289898 251956 290391
rect 252098 290320 252154 290329
rect 252098 290255 252154 290264
rect 251744 289884 251956 289898
rect 252112 289898 252140 290255
rect 251744 289870 251942 289884
rect 252112 289870 252310 289898
rect 248970 289776 249026 289785
rect 248800 289734 248970 289762
rect 248970 289711 249026 289720
rect 248142 289640 248198 289649
rect 248142 289575 248198 289584
rect 252480 289513 252508 312598
rect 253216 299742 253244 382366
rect 254584 382288 254636 382294
rect 254584 382230 254636 382236
rect 253848 378276 253900 378282
rect 253848 378218 253900 378224
rect 253296 359508 253348 359514
rect 253296 359450 253348 359456
rect 253204 299736 253256 299742
rect 253204 299678 253256 299684
rect 252558 292224 252614 292233
rect 252558 292159 252614 292168
rect 252572 291990 252600 292159
rect 252836 292120 252888 292126
rect 252836 292062 252888 292068
rect 252560 291984 252612 291990
rect 252560 291926 252612 291932
rect 252572 289898 252600 291926
rect 252848 290601 252876 292062
rect 252834 290592 252890 290601
rect 252834 290527 252890 290536
rect 252848 289898 252876 290527
rect 253216 289898 253244 299678
rect 253308 291514 253336 359450
rect 253756 318776 253808 318782
rect 253756 318718 253808 318724
rect 253768 316985 253796 318718
rect 253754 316976 253810 316985
rect 253754 316911 253810 316920
rect 253664 312724 253716 312730
rect 253664 312666 253716 312672
rect 253296 291508 253348 291514
rect 253296 291450 253348 291456
rect 252572 289870 252678 289898
rect 252848 289870 253046 289898
rect 253216 289870 253414 289898
rect 253676 289513 253704 312666
rect 253756 291508 253808 291514
rect 253756 291450 253808 291456
rect 253768 289884 253796 291450
rect 253860 290562 253888 378218
rect 254492 294840 254544 294846
rect 254492 294782 254544 294788
rect 254504 291718 254532 294782
rect 254492 291712 254544 291718
rect 254492 291654 254544 291660
rect 253848 290556 253900 290562
rect 253848 290498 253900 290504
rect 253860 290170 253888 290498
rect 253860 290142 253980 290170
rect 253952 289898 253980 290142
rect 253952 289870 254150 289898
rect 254504 289884 254532 291654
rect 254596 291446 254624 382230
rect 254768 379840 254820 379846
rect 254768 379782 254820 379788
rect 254676 376780 254728 376786
rect 254676 376722 254728 376728
rect 254584 291440 254636 291446
rect 254584 291382 254636 291388
rect 254596 290170 254624 291382
rect 254688 290630 254716 376722
rect 254780 298178 254808 379782
rect 255332 300830 255360 385018
rect 255964 379704 256016 379710
rect 255964 379646 256016 379652
rect 255320 300824 255372 300830
rect 255320 300766 255372 300772
rect 254768 298172 254820 298178
rect 254768 298114 254820 298120
rect 254780 291650 254808 298114
rect 255976 298110 256004 379646
rect 256056 362228 256108 362234
rect 256056 362170 256108 362176
rect 255964 298104 256016 298110
rect 255964 298046 256016 298052
rect 256068 296714 256096 362170
rect 256620 318782 256648 398103
rect 257988 398074 258040 398080
rect 257804 396636 257856 396642
rect 257804 396578 257856 396584
rect 257344 383716 257396 383722
rect 257344 383658 257396 383664
rect 256700 345704 256752 345710
rect 256700 345646 256752 345652
rect 256712 345098 256740 345646
rect 256700 345092 256752 345098
rect 256700 345034 256752 345040
rect 256608 318776 256660 318782
rect 256608 318718 256660 318724
rect 256712 301374 256740 345034
rect 257066 318472 257122 318481
rect 257066 318407 257122 318416
rect 256792 318368 256844 318374
rect 256792 318310 256844 318316
rect 256804 318238 256832 318310
rect 256792 318232 256844 318238
rect 256792 318174 256844 318180
rect 257080 317898 257108 318407
rect 257068 317892 257120 317898
rect 257068 317834 257120 317840
rect 257158 310448 257214 310457
rect 257158 310383 257214 310392
rect 257172 309505 257200 310383
rect 257158 309496 257214 309505
rect 257158 309431 257214 309440
rect 256700 301368 256752 301374
rect 256700 301310 256752 301316
rect 257252 301368 257304 301374
rect 257252 301310 257304 301316
rect 256712 300966 256740 301310
rect 256700 300960 256752 300966
rect 256700 300902 256752 300908
rect 256148 300824 256200 300830
rect 256148 300766 256200 300772
rect 256160 299674 256188 300766
rect 256148 299668 256200 299674
rect 256148 299610 256200 299616
rect 255976 296686 256096 296714
rect 254768 291644 254820 291650
rect 254768 291586 254820 291592
rect 255596 291644 255648 291650
rect 255596 291586 255648 291592
rect 254676 290624 254728 290630
rect 254676 290566 254728 290572
rect 254688 290306 254716 290566
rect 254688 290278 255084 290306
rect 254596 290142 254716 290170
rect 254688 289898 254716 290142
rect 255056 289898 255084 290278
rect 254688 289870 254886 289898
rect 255056 289870 255254 289898
rect 255608 289884 255636 291586
rect 255976 291378 256004 296686
rect 256160 291786 256188 299610
rect 256332 298104 256384 298110
rect 256332 298046 256384 298052
rect 256344 297294 256372 298046
rect 256332 297288 256384 297294
rect 256332 297230 256384 297236
rect 256148 291780 256200 291786
rect 256148 291722 256200 291728
rect 255964 291372 256016 291378
rect 255964 291314 256016 291320
rect 255976 289884 256004 291314
rect 256344 289884 256372 297230
rect 256976 293548 257028 293554
rect 256976 293490 257028 293496
rect 256988 292330 257016 293490
rect 256976 292324 257028 292330
rect 256976 292266 257028 292272
rect 257068 292188 257120 292194
rect 257068 292130 257120 292136
rect 256700 291780 256752 291786
rect 256700 291722 256752 291728
rect 256792 291780 256844 291786
rect 256792 291722 256844 291728
rect 256516 290692 256568 290698
rect 256516 290634 256568 290640
rect 256528 290018 256556 290634
rect 256516 290012 256568 290018
rect 256516 289954 256568 289960
rect 256712 289884 256740 291722
rect 256804 290698 256832 291722
rect 256792 290692 256844 290698
rect 256792 290634 256844 290640
rect 257080 289884 257108 292130
rect 257264 290170 257292 301310
rect 257356 293554 257384 383658
rect 257436 351212 257488 351218
rect 257436 351154 257488 351160
rect 257344 293548 257396 293554
rect 257344 293490 257396 293496
rect 257448 292194 257476 351154
rect 257816 318374 257844 396578
rect 257896 388476 257948 388482
rect 257896 388418 257948 388424
rect 257804 318368 257856 318374
rect 257804 318310 257856 318316
rect 257908 310457 257936 388418
rect 258000 317898 258028 398074
rect 259366 398032 259422 398041
rect 259366 397967 259422 397976
rect 259276 389836 259328 389842
rect 259276 389778 259328 389784
rect 258724 382356 258776 382362
rect 258724 382298 258776 382304
rect 258356 319456 258408 319462
rect 258356 319398 258408 319404
rect 257988 317892 258040 317898
rect 257988 317834 258040 317840
rect 257894 310448 257950 310457
rect 257894 310383 257950 310392
rect 257436 292188 257488 292194
rect 257436 292130 257488 292136
rect 258172 292188 258224 292194
rect 258172 292130 258224 292136
rect 257264 290142 257660 290170
rect 257252 290012 257304 290018
rect 257252 289954 257304 289960
rect 257264 289898 257292 289954
rect 257632 289898 257660 290142
rect 257264 289870 257462 289898
rect 257632 289870 257830 289898
rect 258184 289884 258212 292130
rect 258368 289950 258396 319398
rect 258736 297362 258764 382298
rect 259184 378344 259236 378350
rect 259184 378286 259236 378292
rect 258816 375012 258868 375018
rect 258816 374954 258868 374960
rect 258724 297356 258776 297362
rect 258724 297298 258776 297304
rect 258736 292330 258764 297298
rect 258724 292324 258776 292330
rect 258724 292266 258776 292272
rect 258540 292256 258592 292262
rect 258828 292210 258856 374954
rect 259196 372570 259224 378286
rect 259184 372564 259236 372570
rect 259184 372506 259236 372512
rect 259196 371278 259224 372506
rect 259184 371272 259236 371278
rect 259184 371214 259236 371220
rect 258908 370592 258960 370598
rect 258908 370534 258960 370540
rect 258920 319462 258948 370534
rect 258908 319456 258960 319462
rect 258908 319398 258960 319404
rect 259288 310457 259316 389778
rect 259380 310486 259408 397967
rect 260654 389872 260710 389881
rect 260654 389807 260710 389816
rect 260470 388376 260526 388385
rect 260470 388311 260526 388320
rect 259828 379568 259880 379574
rect 259828 379510 259880 379516
rect 259552 374944 259604 374950
rect 259552 374886 259604 374892
rect 259368 310480 259420 310486
rect 259274 310448 259330 310457
rect 259368 310422 259420 310428
rect 259274 310383 259330 310392
rect 259288 309641 259316 310383
rect 259380 309942 259408 310422
rect 259368 309936 259420 309942
rect 259368 309878 259420 309884
rect 259274 309632 259330 309641
rect 259274 309567 259330 309576
rect 259276 298104 259328 298110
rect 259276 298046 259328 298052
rect 258592 292204 258856 292210
rect 258540 292198 258856 292204
rect 258908 292256 258960 292262
rect 258908 292198 258960 292204
rect 258552 292182 258856 292198
rect 258356 289944 258408 289950
rect 258408 289892 258566 289898
rect 258356 289886 258566 289892
rect 258368 289870 258566 289886
rect 258920 289884 258948 292198
rect 259288 290358 259316 298046
rect 259276 290352 259328 290358
rect 259276 290294 259328 290300
rect 259288 289884 259316 290294
rect 259564 290086 259592 374886
rect 259736 371272 259788 371278
rect 259736 371214 259788 371220
rect 259644 308508 259696 308514
rect 259644 308450 259696 308456
rect 259656 305114 259684 308450
rect 259644 305108 259696 305114
rect 259644 305050 259696 305056
rect 259656 293078 259684 305050
rect 259644 293072 259696 293078
rect 259644 293014 259696 293020
rect 259748 291786 259776 371214
rect 259840 306374 259868 379510
rect 260484 322969 260512 388311
rect 260562 387016 260618 387025
rect 260562 386951 260618 386960
rect 260470 322960 260526 322969
rect 260470 322895 260526 322904
rect 260484 322318 260512 322895
rect 260472 322312 260524 322318
rect 260472 322254 260524 322260
rect 260472 314220 260524 314226
rect 260472 314162 260524 314168
rect 260484 309126 260512 314162
rect 260576 313274 260604 386951
rect 260668 314226 260696 389807
rect 260656 314220 260708 314226
rect 260656 314162 260708 314168
rect 260760 314106 260788 398210
rect 262034 391232 262090 391241
rect 262034 391167 262090 391176
rect 261484 381132 261536 381138
rect 261484 381074 261536 381080
rect 260668 314078 260788 314106
rect 260564 313268 260616 313274
rect 260564 313210 260616 313216
rect 260668 310185 260696 314078
rect 260748 313268 260800 313274
rect 260748 313210 260800 313216
rect 260760 312798 260788 313210
rect 260748 312792 260800 312798
rect 260748 312734 260800 312740
rect 260654 310176 260710 310185
rect 260654 310111 260710 310120
rect 260472 309120 260524 309126
rect 260472 309062 260524 309068
rect 260748 309120 260800 309126
rect 260748 309062 260800 309068
rect 260760 308582 260788 309062
rect 260748 308576 260800 308582
rect 260748 308518 260800 308524
rect 259840 306346 260604 306374
rect 260196 293072 260248 293078
rect 260196 293014 260248 293020
rect 260012 292324 260064 292330
rect 260012 292266 260064 292272
rect 259736 291780 259788 291786
rect 259736 291722 259788 291728
rect 259552 290080 259604 290086
rect 259552 290022 259604 290028
rect 259564 289898 259592 290022
rect 259564 289870 259670 289898
rect 260024 289884 260052 292266
rect 260208 289898 260236 293014
rect 260576 290290 260604 306346
rect 261300 304632 261352 304638
rect 261300 304574 261352 304580
rect 261312 303686 261340 304574
rect 261300 303680 261352 303686
rect 261300 303622 261352 303628
rect 260932 302252 260984 302258
rect 260932 302194 260984 302200
rect 260564 290284 260616 290290
rect 260564 290226 260616 290232
rect 260576 289898 260604 290226
rect 260944 289898 260972 302194
rect 261312 289898 261340 303622
rect 261496 292097 261524 381074
rect 261576 376100 261628 376106
rect 261576 376042 261628 376048
rect 261482 292088 261538 292097
rect 261482 292023 261538 292032
rect 261588 290766 261616 376042
rect 261668 375556 261720 375562
rect 261668 375498 261720 375504
rect 261680 295730 261708 375498
rect 261760 349852 261812 349858
rect 261760 349794 261812 349800
rect 261772 304638 261800 349794
rect 262048 311846 262076 391167
rect 262128 388544 262180 388550
rect 262128 388486 262180 388492
rect 262036 311840 262088 311846
rect 262036 311782 262088 311788
rect 262048 311234 262076 311782
rect 262036 311228 262088 311234
rect 262036 311170 262088 311176
rect 261760 304632 261812 304638
rect 261760 304574 261812 304580
rect 262140 302161 262168 388486
rect 262864 386504 262916 386510
rect 262864 386446 262916 386452
rect 262220 378208 262272 378214
rect 262220 378150 262272 378156
rect 262126 302152 262182 302161
rect 262126 302087 262182 302096
rect 262140 301617 262168 302087
rect 262126 301608 262182 301617
rect 262126 301543 262182 301552
rect 261668 295724 261720 295730
rect 261668 295666 261720 295672
rect 261576 290760 261628 290766
rect 261576 290702 261628 290708
rect 261680 289898 261708 295666
rect 262232 290834 262260 378150
rect 262312 301368 262364 301374
rect 262312 301310 262364 301316
rect 262324 300898 262352 301310
rect 262312 300892 262364 300898
rect 262312 300834 262364 300840
rect 262324 293078 262352 300834
rect 262876 300830 262904 386446
rect 262956 383852 263008 383858
rect 262956 383794 263008 383800
rect 262968 301374 262996 383794
rect 263048 376848 263100 376854
rect 263048 376790 263100 376796
rect 262956 301368 263008 301374
rect 262956 301310 263008 301316
rect 262404 300824 262456 300830
rect 262404 300766 262456 300772
rect 262864 300824 262916 300830
rect 262864 300766 262916 300772
rect 262416 299606 262444 300766
rect 262404 299600 262456 299606
rect 262404 299542 262456 299548
rect 262312 293072 262364 293078
rect 262312 293014 262364 293020
rect 262220 290828 262272 290834
rect 262220 290770 262272 290776
rect 262232 290222 262260 290770
rect 262220 290216 262272 290222
rect 262220 290158 262272 290164
rect 262416 289898 262444 299542
rect 263060 298246 263088 376790
rect 263336 322998 263364 401775
rect 265622 401704 265678 401713
rect 265622 401639 265678 401648
rect 264886 398304 264942 398313
rect 264886 398239 264942 398248
rect 264796 394120 264848 394126
rect 264796 394062 264848 394068
rect 263506 391368 263562 391377
rect 263506 391303 263562 391312
rect 263416 387184 263468 387190
rect 263416 387126 263468 387132
rect 263324 322992 263376 322998
rect 263324 322934 263376 322940
rect 263336 322250 263364 322934
rect 263324 322244 263376 322250
rect 263324 322186 263376 322192
rect 263428 307766 263456 387126
rect 263520 308553 263548 391303
rect 264520 385144 264572 385150
rect 264520 385086 264572 385092
rect 264336 380928 264388 380934
rect 264336 380870 264388 380876
rect 264244 375896 264296 375902
rect 264244 375838 264296 375844
rect 263690 318200 263746 318209
rect 263690 318135 263746 318144
rect 263704 317665 263732 318135
rect 263690 317656 263746 317665
rect 263690 317591 263746 317600
rect 263506 308544 263562 308553
rect 263506 308479 263562 308488
rect 263140 307760 263192 307766
rect 263140 307702 263192 307708
rect 263416 307760 263468 307766
rect 263416 307702 263468 307708
rect 263152 307222 263180 307702
rect 263140 307216 263192 307222
rect 263140 307158 263192 307164
rect 264060 303816 264112 303822
rect 264060 303758 264112 303764
rect 263048 298240 263100 298246
rect 263048 298182 263100 298188
rect 263060 292330 263088 298182
rect 264072 297498 264100 303758
rect 264256 302234 264284 375838
rect 264164 302206 264284 302234
rect 264060 297492 264112 297498
rect 264060 297434 264112 297440
rect 263140 293072 263192 293078
rect 263140 293014 263192 293020
rect 263048 292324 263100 292330
rect 263048 292266 263100 292272
rect 262588 291236 262640 291242
rect 262588 291178 262640 291184
rect 260208 289870 260406 289898
rect 260576 289870 260774 289898
rect 260944 289870 261142 289898
rect 261312 289870 261510 289898
rect 261680 289870 261878 289898
rect 262246 289870 262444 289898
rect 262600 289884 262628 291178
rect 262956 290828 263008 290834
rect 262956 290770 263008 290776
rect 262968 289884 262996 290770
rect 263152 289898 263180 293014
rect 264164 292574 264192 302206
rect 264244 297492 264296 297498
rect 264244 297434 264296 297440
rect 263980 292546 264192 292574
rect 263980 292126 264008 292546
rect 264060 292324 264112 292330
rect 264060 292266 264112 292272
rect 263968 292120 264020 292126
rect 263968 292062 264020 292068
rect 263692 291304 263744 291310
rect 263692 291246 263744 291252
rect 263152 289870 263350 289898
rect 263704 289884 263732 291246
rect 264072 289884 264100 292266
rect 264256 289898 264284 297434
rect 264348 297158 264376 380870
rect 264428 374400 264480 374406
rect 264428 374342 264480 374348
rect 264336 297152 264388 297158
rect 264336 297094 264388 297100
rect 264348 292262 264376 297094
rect 264336 292256 264388 292262
rect 264336 292198 264388 292204
rect 264440 291854 264468 374342
rect 264532 303822 264560 385086
rect 264612 374536 264664 374542
rect 264612 374478 264664 374484
rect 264520 303816 264572 303822
rect 264520 303758 264572 303764
rect 264520 302252 264572 302258
rect 264520 302194 264572 302200
rect 264532 292330 264560 302194
rect 264624 294778 264652 374478
rect 264808 316033 264836 394062
rect 264900 317665 264928 398239
rect 264886 317656 264942 317665
rect 264886 317591 264942 317600
rect 264794 316024 264850 316033
rect 264794 315959 264796 315968
rect 264848 315959 264850 315968
rect 264796 315930 264848 315936
rect 264808 315899 264836 315930
rect 264888 308576 264940 308582
rect 264888 308518 264940 308524
rect 264900 302258 264928 308518
rect 264980 304904 265032 304910
rect 264980 304846 265032 304852
rect 264992 304502 265020 304846
rect 264980 304496 265032 304502
rect 264980 304438 265032 304444
rect 264888 302252 264940 302258
rect 264888 302194 264940 302200
rect 265636 298314 265664 401639
rect 265716 382492 265768 382498
rect 265716 382434 265768 382440
rect 265624 298308 265676 298314
rect 265624 298250 265676 298256
rect 265728 298110 265756 382434
rect 265820 321706 265848 402047
rect 266266 401976 266322 401985
rect 266266 401911 266322 401920
rect 266174 390008 266230 390017
rect 266174 389943 266230 389952
rect 265900 383784 265952 383790
rect 265900 383726 265952 383732
rect 265808 321700 265860 321706
rect 265808 321642 265860 321648
rect 265820 317830 265848 321642
rect 265808 317824 265860 317830
rect 265808 317766 265860 317772
rect 265912 305046 265940 383726
rect 265992 370320 266044 370326
rect 265992 370262 266044 370268
rect 265900 305040 265952 305046
rect 265900 304982 265952 304988
rect 265716 298104 265768 298110
rect 265716 298046 265768 298052
rect 264612 294772 264664 294778
rect 264612 294714 264664 294720
rect 265912 292574 265940 304982
rect 266004 296138 266032 370262
rect 266188 304910 266216 389943
rect 266280 307193 266308 401911
rect 271696 400444 271748 400450
rect 271696 400386 271748 400392
rect 267002 400344 267058 400353
rect 267002 400279 267058 400288
rect 266360 311772 266412 311778
rect 266360 311714 266412 311720
rect 266372 311166 266400 311714
rect 266360 311160 266412 311166
rect 266360 311102 266412 311108
rect 266266 307184 266322 307193
rect 266266 307119 266322 307128
rect 267016 306406 267044 400279
rect 270130 396944 270186 396953
rect 270130 396879 270186 396888
rect 270038 396808 270094 396817
rect 270038 396743 270094 396752
rect 267648 395140 267700 395146
rect 267648 395082 267700 395088
rect 267556 391264 267608 391270
rect 267556 391206 267608 391212
rect 267188 376032 267240 376038
rect 267188 375974 267240 375980
rect 267096 375964 267148 375970
rect 267096 375906 267148 375912
rect 267004 306400 267056 306406
rect 267004 306342 267056 306348
rect 266360 306332 266412 306338
rect 266360 306274 266412 306280
rect 266372 305726 266400 306274
rect 266360 305720 266412 305726
rect 266360 305662 266412 305668
rect 266176 304904 266228 304910
rect 266176 304846 266228 304852
rect 267016 304774 267044 306342
rect 267004 304768 267056 304774
rect 267004 304710 267056 304716
rect 265992 296132 266044 296138
rect 265992 296074 266044 296080
rect 265728 292546 265940 292574
rect 264520 292324 264572 292330
rect 264520 292266 264572 292272
rect 265532 292324 265584 292330
rect 265532 292266 265584 292272
rect 265164 292256 265216 292262
rect 265164 292198 265216 292204
rect 264428 291848 264480 291854
rect 264428 291790 264480 291796
rect 264796 291372 264848 291378
rect 264796 291314 264848 291320
rect 264256 289870 264454 289898
rect 264808 289884 264836 291314
rect 265176 289884 265204 292198
rect 265544 289884 265572 292266
rect 265728 289898 265756 292546
rect 267108 290465 267136 375906
rect 267200 291961 267228 375974
rect 267280 374196 267332 374202
rect 267280 374138 267332 374144
rect 267292 292058 267320 374138
rect 267464 372904 267516 372910
rect 267464 372846 267516 372852
rect 267280 292052 267332 292058
rect 267280 291994 267332 292000
rect 267186 291952 267242 291961
rect 267186 291887 267242 291896
rect 267094 290456 267150 290465
rect 267094 290391 267150 290400
rect 265728 289870 265926 289898
rect 258368 289821 258396 289870
rect 247038 289504 247094 289513
rect 246960 289462 247038 289490
rect 247038 289439 247094 289448
rect 248050 289504 248106 289513
rect 248050 289439 248106 289448
rect 252466 289504 252522 289513
rect 252466 289439 252522 289448
rect 253662 289504 253718 289513
rect 253662 289439 253718 289448
rect 244004 289400 244056 289406
rect 237852 289377 237972 289388
rect 237852 289368 237986 289377
rect 237852 289360 237930 289368
rect 235540 289342 235592 289348
rect 237930 289303 237986 289312
rect 241242 289368 241298 289377
rect 244004 289342 244056 289348
rect 245476 289400 245528 289406
rect 245476 289342 245528 289348
rect 241242 289303 241298 289312
rect 267476 288561 267504 372846
rect 267568 311778 267596 391206
rect 267556 311772 267608 311778
rect 267556 311714 267608 311720
rect 267660 306338 267688 395082
rect 269026 391504 269082 391513
rect 269026 391439 269082 391448
rect 268658 390144 268714 390153
rect 268658 390079 268714 390088
rect 268384 381064 268436 381070
rect 268384 381006 268436 381012
rect 267648 306332 267700 306338
rect 267648 306274 267700 306280
rect 268396 291378 268424 381006
rect 268568 358080 268620 358086
rect 268568 358022 268620 358028
rect 268580 357474 268608 358022
rect 268568 357468 268620 357474
rect 268568 357410 268620 357416
rect 268580 354674 268608 357410
rect 268488 354646 268608 354674
rect 268488 292194 268516 354646
rect 268672 321094 268700 390079
rect 268842 388512 268898 388521
rect 268842 388447 268898 388456
rect 268750 385656 268806 385665
rect 268750 385591 268806 385600
rect 268660 321088 268712 321094
rect 268660 321030 268712 321036
rect 268764 316034 268792 385591
rect 268856 317422 268884 388447
rect 268936 385824 268988 385830
rect 268936 385766 268988 385772
rect 268844 317416 268896 317422
rect 268844 317358 268896 317364
rect 268580 316006 268792 316034
rect 268948 316034 268976 385766
rect 269040 318578 269068 391439
rect 269856 389904 269908 389910
rect 269856 389846 269908 389852
rect 269486 320512 269542 320521
rect 269486 320447 269542 320456
rect 269500 319802 269528 320447
rect 269488 319796 269540 319802
rect 269488 319738 269540 319744
rect 269764 319252 269816 319258
rect 269764 319194 269816 319200
rect 269028 318572 269080 318578
rect 269028 318514 269080 318520
rect 269040 318102 269068 318514
rect 269028 318096 269080 318102
rect 269028 318038 269080 318044
rect 269580 317416 269632 317422
rect 269580 317358 269632 317364
rect 268948 316006 269068 316034
rect 269592 316033 269620 317358
rect 268580 315761 268608 316006
rect 268566 315752 268622 315761
rect 268566 315687 268622 315696
rect 268580 315217 268608 315687
rect 268566 315208 268622 315217
rect 268566 315143 268622 315152
rect 269040 314537 269068 316006
rect 269578 316024 269634 316033
rect 269578 315959 269634 315968
rect 269026 314528 269082 314537
rect 269026 314463 269082 314472
rect 269040 313721 269068 314463
rect 269026 313712 269082 313721
rect 269026 313647 269082 313656
rect 268476 292188 268528 292194
rect 268476 292130 268528 292136
rect 268384 291372 268436 291378
rect 268384 291314 268436 291320
rect 269028 291372 269080 291378
rect 269028 291314 269080 291320
rect 269040 291174 269068 291314
rect 269028 291168 269080 291174
rect 269028 291110 269080 291116
rect 267462 288552 267518 288561
rect 267462 288487 267518 288496
rect 268384 287700 268436 287706
rect 268384 287642 268436 287648
rect 267554 257272 267610 257281
rect 267554 257207 267610 257216
rect 267568 252554 267596 257207
rect 267568 252526 267688 252554
rect 267554 249248 267610 249257
rect 267554 249183 267610 249192
rect 222292 241596 222344 241602
rect 222292 241538 222344 241544
rect 222304 240106 222332 241538
rect 267568 240530 267596 249183
rect 267660 248414 267688 252526
rect 268014 250608 268070 250617
rect 268014 250543 268070 250552
rect 267660 248386 267872 248414
rect 267738 247616 267794 247625
rect 267738 247551 267794 247560
rect 267398 240502 267596 240530
rect 267568 240428 267596 240502
rect 267568 240400 267688 240428
rect 267660 240156 267688 240400
rect 267752 240310 267780 247551
rect 267740 240304 267792 240310
rect 267740 240246 267792 240252
rect 267660 240128 267780 240156
rect 222292 240100 222344 240106
rect 222292 240042 222344 240048
rect 222534 239970 222562 240108
rect 222626 239970 222654 240108
rect 222718 239970 222746 240108
rect 222522 239964 222574 239970
rect 222522 239906 222574 239912
rect 222614 239964 222666 239970
rect 222614 239906 222666 239912
rect 222706 239964 222758 239970
rect 222706 239906 222758 239912
rect 222384 239896 222436 239902
rect 222810 239850 222838 240108
rect 222902 239902 222930 240108
rect 222994 239907 223022 240108
rect 223086 239970 223114 240108
rect 223178 239970 223206 240108
rect 223074 239964 223126 239970
rect 222384 239838 222436 239844
rect 222200 239692 222252 239698
rect 222200 239634 222252 239640
rect 222120 239448 222240 239476
rect 222108 238876 222160 238882
rect 222108 238818 222160 238824
rect 222014 236464 222070 236473
rect 222014 236399 222070 236408
rect 222028 224942 222056 236399
rect 222016 224936 222068 224942
rect 222016 224878 222068 224884
rect 221924 212288 221976 212294
rect 221924 212230 221976 212236
rect 221832 212152 221884 212158
rect 221832 212094 221884 212100
rect 221740 212016 221792 212022
rect 221740 211958 221792 211964
rect 222028 150113 222056 224878
rect 222120 155650 222148 238818
rect 222212 214606 222240 239448
rect 222396 223574 222424 239838
rect 222764 239822 222838 239850
rect 222890 239896 222942 239902
rect 222890 239838 222942 239844
rect 222980 239898 223036 239907
rect 223074 239906 223126 239912
rect 223166 239964 223218 239970
rect 223166 239906 223218 239912
rect 222980 239833 223036 239842
rect 223270 239850 223298 240108
rect 223362 239970 223390 240108
rect 223454 239970 223482 240108
rect 223546 239970 223574 240108
rect 223638 239970 223666 240108
rect 223730 239970 223758 240108
rect 223350 239964 223402 239970
rect 223350 239906 223402 239912
rect 223442 239964 223494 239970
rect 223442 239906 223494 239912
rect 223534 239964 223586 239970
rect 223534 239906 223586 239912
rect 223626 239964 223678 239970
rect 223626 239906 223678 239912
rect 223718 239964 223770 239970
rect 223718 239906 223770 239912
rect 223670 239864 223726 239873
rect 223120 239828 223172 239834
rect 222764 239737 222792 239822
rect 223270 239822 223344 239850
rect 223120 239770 223172 239776
rect 222844 239760 222896 239766
rect 222750 239728 222806 239737
rect 222844 239702 222896 239708
rect 222750 239663 222806 239672
rect 222568 238468 222620 238474
rect 222568 238410 222620 238416
rect 222580 238202 222608 238410
rect 222764 238338 222792 239663
rect 222856 238678 222884 239702
rect 223132 239465 223160 239770
rect 223316 239612 223344 239822
rect 223822 239850 223850 240108
rect 223914 239970 223942 240108
rect 223902 239964 223954 239970
rect 223902 239906 223954 239912
rect 224006 239850 224034 240108
rect 224098 239902 224126 240108
rect 224190 239970 224218 240108
rect 224282 239970 224310 240108
rect 224374 239970 224402 240108
rect 224178 239964 224230 239970
rect 224178 239906 224230 239912
rect 224270 239964 224322 239970
rect 224270 239906 224322 239912
rect 224362 239964 224414 239970
rect 224362 239906 224414 239912
rect 223592 239808 223670 239816
rect 223592 239788 223672 239808
rect 223396 239760 223448 239766
rect 223394 239728 223396 239737
rect 223488 239760 223540 239766
rect 223448 239728 223450 239737
rect 223488 239702 223540 239708
rect 223394 239663 223450 239672
rect 223316 239584 223436 239612
rect 223118 239456 223174 239465
rect 223118 239391 223174 239400
rect 223304 239420 223356 239426
rect 222844 238672 222896 238678
rect 222844 238614 222896 238620
rect 222844 238468 222896 238474
rect 222844 238410 222896 238416
rect 222752 238332 222804 238338
rect 222752 238274 222804 238280
rect 222568 238196 222620 238202
rect 222568 238138 222620 238144
rect 222568 235068 222620 235074
rect 222568 235010 222620 235016
rect 222580 233170 222608 235010
rect 222568 233164 222620 233170
rect 222568 233106 222620 233112
rect 222304 223546 222424 223574
rect 222304 215966 222332 223546
rect 222580 219434 222608 233106
rect 222396 219406 222608 219434
rect 222292 215960 222344 215966
rect 222292 215902 222344 215908
rect 222200 214600 222252 214606
rect 222200 214542 222252 214548
rect 222396 159254 222424 219406
rect 222384 159248 222436 159254
rect 222384 159190 222436 159196
rect 222108 155644 222160 155650
rect 222108 155586 222160 155592
rect 222014 150104 222070 150113
rect 222014 150039 222070 150048
rect 222200 146872 222252 146878
rect 222200 146814 222252 146820
rect 221646 142624 221702 142633
rect 221646 142559 221702 142568
rect 222212 16574 222240 146814
rect 222856 145518 222884 238410
rect 223132 231266 223160 239391
rect 223304 239362 223356 239368
rect 223120 231260 223172 231266
rect 223120 231202 223172 231208
rect 223212 230240 223264 230246
rect 223212 230182 223264 230188
rect 222936 229220 222988 229226
rect 222936 229162 222988 229168
rect 222844 145512 222896 145518
rect 222844 145454 222896 145460
rect 222948 144158 222976 229162
rect 223028 227316 223080 227322
rect 223028 227258 223080 227264
rect 223040 146878 223068 227258
rect 223120 221740 223172 221746
rect 223120 221682 223172 221688
rect 223028 146872 223080 146878
rect 223028 146814 223080 146820
rect 222936 144152 222988 144158
rect 222936 144094 222988 144100
rect 223132 141273 223160 221682
rect 223224 150958 223252 230182
rect 223316 159186 223344 239362
rect 223408 238785 223436 239584
rect 223500 239494 223528 239702
rect 223488 239488 223540 239494
rect 223488 239430 223540 239436
rect 223394 238776 223450 238785
rect 223394 238711 223450 238720
rect 223408 192506 223436 238711
rect 223592 238406 223620 239788
rect 223724 239799 223726 239808
rect 223776 239822 223850 239850
rect 223960 239822 224034 239850
rect 224086 239896 224138 239902
rect 224086 239838 224138 239844
rect 224224 239828 224276 239834
rect 223672 239770 223724 239776
rect 223672 239692 223724 239698
rect 223672 239634 223724 239640
rect 223580 238400 223632 238406
rect 223580 238342 223632 238348
rect 223684 236638 223712 239634
rect 223776 238746 223804 239822
rect 223960 239737 223988 239822
rect 224224 239770 224276 239776
rect 224316 239828 224368 239834
rect 224316 239770 224368 239776
rect 223946 239728 224002 239737
rect 223946 239663 224002 239672
rect 224132 239624 224184 239630
rect 224132 239566 224184 239572
rect 224038 239456 224094 239465
rect 224038 239391 224094 239400
rect 223946 238776 224002 238785
rect 223764 238740 223816 238746
rect 223946 238711 224002 238720
rect 223764 238682 223816 238688
rect 223672 236632 223724 236638
rect 223672 236574 223724 236580
rect 223578 220688 223634 220697
rect 223578 220623 223634 220632
rect 223592 218006 223620 220623
rect 223684 220153 223712 236574
rect 223764 234388 223816 234394
rect 223764 234330 223816 234336
rect 223776 233102 223804 234330
rect 223856 233368 223908 233374
rect 223856 233310 223908 233316
rect 223764 233096 223816 233102
rect 223764 233038 223816 233044
rect 223670 220144 223726 220153
rect 223670 220079 223726 220088
rect 223580 218000 223632 218006
rect 223580 217942 223632 217948
rect 223396 192500 223448 192506
rect 223396 192442 223448 192448
rect 223304 159180 223356 159186
rect 223304 159122 223356 159128
rect 223212 150952 223264 150958
rect 223212 150894 223264 150900
rect 223118 141264 223174 141273
rect 223118 141199 223174 141208
rect 223776 137834 223804 233038
rect 223868 141778 223896 233310
rect 223960 184249 223988 238711
rect 224052 186998 224080 239391
rect 224144 239057 224172 239566
rect 224236 239222 224264 239770
rect 224224 239216 224276 239222
rect 224224 239158 224276 239164
rect 224130 239048 224186 239057
rect 224130 238983 224186 238992
rect 224224 238740 224276 238746
rect 224224 238682 224276 238688
rect 224130 238504 224186 238513
rect 224130 238439 224186 238448
rect 224144 196654 224172 238439
rect 224236 235890 224264 238682
rect 224328 237250 224356 239770
rect 224466 239714 224494 240108
rect 224558 239902 224586 240108
rect 224650 239970 224678 240108
rect 224638 239964 224690 239970
rect 224638 239906 224690 239912
rect 224742 239902 224770 240108
rect 224834 239970 224862 240108
rect 224926 239970 224954 240108
rect 225018 239970 225046 240108
rect 224822 239964 224874 239970
rect 224822 239906 224874 239912
rect 224914 239964 224966 239970
rect 224914 239906 224966 239912
rect 225006 239964 225058 239970
rect 225006 239906 225058 239912
rect 224546 239896 224598 239902
rect 224546 239838 224598 239844
rect 224730 239896 224782 239902
rect 224730 239838 224782 239844
rect 224868 239828 224920 239834
rect 224868 239770 224920 239776
rect 224420 239686 224494 239714
rect 224592 239760 224644 239766
rect 224592 239702 224644 239708
rect 224684 239760 224736 239766
rect 224684 239702 224736 239708
rect 224420 239494 224448 239686
rect 224500 239624 224552 239630
rect 224500 239566 224552 239572
rect 224408 239488 224460 239494
rect 224512 239465 224540 239566
rect 224408 239430 224460 239436
rect 224498 239456 224554 239465
rect 224498 239391 224554 239400
rect 224500 239352 224552 239358
rect 224500 239294 224552 239300
rect 224408 239216 224460 239222
rect 224408 239158 224460 239164
rect 224420 238377 224448 239158
rect 224406 238368 224462 238377
rect 224406 238303 224462 238312
rect 224512 237658 224540 239294
rect 224500 237652 224552 237658
rect 224500 237594 224552 237600
rect 224316 237244 224368 237250
rect 224316 237186 224368 237192
rect 224408 235952 224460 235958
rect 224408 235894 224460 235900
rect 224224 235884 224276 235890
rect 224224 235826 224276 235832
rect 224222 223000 224278 223009
rect 224222 222935 224278 222944
rect 224132 196648 224184 196654
rect 224132 196590 224184 196596
rect 224040 186992 224092 186998
rect 224040 186934 224092 186940
rect 223946 184240 224002 184249
rect 223946 184175 224002 184184
rect 224236 143002 224264 222935
rect 224314 221640 224370 221649
rect 224314 221575 224370 221584
rect 224224 142996 224276 143002
rect 224224 142938 224276 142944
rect 223856 141772 223908 141778
rect 223856 141714 223908 141720
rect 224328 141409 224356 221575
rect 224420 213926 224448 235894
rect 224604 219337 224632 239702
rect 224696 239426 224724 239702
rect 224776 239692 224828 239698
rect 224776 239634 224828 239640
rect 224684 239420 224736 239426
rect 224684 239362 224736 239368
rect 224684 239148 224736 239154
rect 224684 239090 224736 239096
rect 224696 224913 224724 239090
rect 224788 236065 224816 239634
rect 224774 236056 224830 236065
rect 224774 235991 224830 236000
rect 224880 235958 224908 239770
rect 224958 239728 225014 239737
rect 225110 239714 225138 240108
rect 225202 239902 225230 240108
rect 225190 239896 225242 239902
rect 225294 239873 225322 240108
rect 225190 239838 225242 239844
rect 225280 239864 225336 239873
rect 225280 239799 225336 239808
rect 225236 239760 225288 239766
rect 225110 239686 225184 239714
rect 225386 239748 225414 240108
rect 225478 239902 225506 240108
rect 225570 239970 225598 240108
rect 225558 239964 225610 239970
rect 225558 239906 225610 239912
rect 225466 239896 225518 239902
rect 225464 239864 225466 239873
rect 225518 239864 225520 239873
rect 225464 239799 225520 239808
rect 225662 239816 225690 240108
rect 225754 239970 225782 240108
rect 225846 239970 225874 240108
rect 225742 239964 225794 239970
rect 225742 239906 225794 239912
rect 225834 239964 225886 239970
rect 225834 239906 225886 239912
rect 225788 239828 225840 239834
rect 225662 239788 225736 239816
rect 225386 239720 225644 239748
rect 225708 239737 225736 239788
rect 225938 239816 225966 240108
rect 225788 239770 225840 239776
rect 225892 239788 225966 239816
rect 226030 239816 226058 240108
rect 226122 239970 226150 240108
rect 226110 239964 226162 239970
rect 226110 239906 226162 239912
rect 226030 239788 226104 239816
rect 225236 239702 225288 239708
rect 224958 239663 224960 239672
rect 225012 239663 225014 239672
rect 224960 239634 225012 239640
rect 225156 239612 225184 239686
rect 225064 239584 225184 239612
rect 225248 239612 225276 239702
rect 225420 239624 225472 239630
rect 225248 239584 225368 239612
rect 224960 239284 225012 239290
rect 224960 239226 225012 239232
rect 224868 235952 224920 235958
rect 224868 235894 224920 235900
rect 224866 235104 224922 235113
rect 224866 235039 224922 235048
rect 224880 233986 224908 235039
rect 224868 233980 224920 233986
rect 224868 233922 224920 233928
rect 224682 224904 224738 224913
rect 224682 224839 224738 224848
rect 224972 219434 225000 239226
rect 225064 239057 225092 239584
rect 225144 239488 225196 239494
rect 225236 239488 225288 239494
rect 225144 239430 225196 239436
rect 225234 239456 225236 239465
rect 225288 239456 225290 239465
rect 225156 239358 225184 239430
rect 225234 239391 225290 239400
rect 225144 239352 225196 239358
rect 225144 239294 225196 239300
rect 225248 239290 225276 239391
rect 225236 239284 225288 239290
rect 225236 239226 225288 239232
rect 225050 239048 225106 239057
rect 225050 238983 225106 238992
rect 225144 239012 225196 239018
rect 225144 238954 225196 238960
rect 225156 237930 225184 238954
rect 225234 238504 225290 238513
rect 225234 238439 225290 238448
rect 225144 237924 225196 237930
rect 225144 237866 225196 237872
rect 225248 228546 225276 238439
rect 225340 238406 225368 239584
rect 225420 239566 225472 239572
rect 225328 238400 225380 238406
rect 225328 238342 225380 238348
rect 225432 238338 225460 239566
rect 225512 239488 225564 239494
rect 225512 239430 225564 239436
rect 225420 238332 225472 238338
rect 225420 238274 225472 238280
rect 225328 238264 225380 238270
rect 225328 238206 225380 238212
rect 225236 228540 225288 228546
rect 225236 228482 225288 228488
rect 224972 219406 225092 219434
rect 224590 219328 224646 219337
rect 224590 219263 224646 219272
rect 225064 215294 225092 219406
rect 225340 216306 225368 238206
rect 225420 229900 225472 229906
rect 225420 229842 225472 229848
rect 225432 218657 225460 229842
rect 225524 220318 225552 239430
rect 225616 238134 225644 239720
rect 225694 239728 225750 239737
rect 225694 239663 225750 239672
rect 225696 239420 225748 239426
rect 225696 239362 225748 239368
rect 225708 238202 225736 239362
rect 225800 239034 225828 239770
rect 225892 239154 225920 239788
rect 225972 239692 226024 239698
rect 225972 239634 226024 239640
rect 225880 239148 225932 239154
rect 225880 239090 225932 239096
rect 225800 239006 225920 239034
rect 225786 238776 225842 238785
rect 225786 238711 225842 238720
rect 225800 238406 225828 238711
rect 225892 238513 225920 239006
rect 225878 238504 225934 238513
rect 225878 238439 225934 238448
rect 225788 238400 225840 238406
rect 225788 238342 225840 238348
rect 225696 238196 225748 238202
rect 225696 238138 225748 238144
rect 225604 238128 225656 238134
rect 225604 238070 225656 238076
rect 225616 228682 225644 238070
rect 225696 232484 225748 232490
rect 225696 232426 225748 232432
rect 225604 228676 225656 228682
rect 225604 228618 225656 228624
rect 225512 220312 225564 220318
rect 225512 220254 225564 220260
rect 225418 218648 225474 218657
rect 225418 218583 225474 218592
rect 225328 216300 225380 216306
rect 225328 216242 225380 216248
rect 224972 215266 225092 215294
rect 224408 213920 224460 213926
rect 224408 213862 224460 213868
rect 224972 169017 225000 215266
rect 225340 209774 225368 216242
rect 225340 209746 225644 209774
rect 224958 169008 225014 169017
rect 224958 168943 225014 168952
rect 225616 161090 225644 209746
rect 225604 161084 225656 161090
rect 225604 161026 225656 161032
rect 225604 155644 225656 155650
rect 225604 155586 225656 155592
rect 224314 141400 224370 141409
rect 224314 141335 224370 141344
rect 223764 137828 223816 137834
rect 223764 137770 223816 137776
rect 223578 135960 223634 135969
rect 223578 135895 223634 135904
rect 222212 16546 222792 16574
rect 221556 3732 221608 3738
rect 221556 3674 221608 3680
rect 220084 3664 220136 3670
rect 220084 3606 220136 3612
rect 221568 480 221596 3674
rect 222764 480 222792 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 135895
rect 225144 3800 225196 3806
rect 225144 3742 225196 3748
rect 225156 480 225184 3742
rect 225616 3602 225644 155586
rect 225708 139126 225736 232426
rect 225800 229906 225828 238342
rect 225880 238196 225932 238202
rect 225880 238138 225932 238144
rect 225892 238105 225920 238138
rect 225878 238096 225934 238105
rect 225878 238031 225934 238040
rect 225984 235414 226012 239634
rect 226076 239494 226104 239788
rect 226214 239748 226242 240108
rect 226306 239873 226334 240108
rect 226398 239970 226426 240108
rect 226490 239970 226518 240108
rect 226386 239964 226438 239970
rect 226386 239906 226438 239912
rect 226478 239964 226530 239970
rect 226478 239906 226530 239912
rect 226292 239864 226348 239873
rect 226292 239799 226348 239808
rect 226430 239864 226486 239873
rect 226582 239850 226610 240108
rect 226486 239822 226610 239850
rect 226430 239799 226486 239808
rect 226168 239720 226242 239748
rect 226064 239488 226116 239494
rect 226064 239430 226116 239436
rect 226064 239012 226116 239018
rect 226064 238954 226116 238960
rect 225972 235408 226024 235414
rect 225972 235350 226024 235356
rect 226076 234394 226104 238954
rect 226168 235074 226196 239720
rect 226306 239680 226334 239799
rect 226524 239760 226576 239766
rect 226674 239748 226702 240108
rect 226766 239902 226794 240108
rect 226858 239970 226886 240108
rect 226846 239964 226898 239970
rect 226846 239906 226898 239912
rect 226754 239896 226806 239902
rect 226754 239838 226806 239844
rect 226950 239850 226978 240108
rect 227042 239970 227070 240108
rect 227030 239964 227082 239970
rect 227030 239906 227082 239912
rect 227134 239873 227162 240108
rect 227226 239902 227254 240108
rect 227318 239970 227346 240108
rect 227306 239964 227358 239970
rect 227306 239906 227358 239912
rect 227214 239896 227266 239902
rect 227120 239864 227176 239873
rect 226950 239822 227024 239850
rect 226800 239760 226852 239766
rect 226674 239720 226748 239748
rect 226524 239702 226576 239708
rect 226260 239652 226334 239680
rect 226432 239692 226484 239698
rect 226156 235068 226208 235074
rect 226156 235010 226208 235016
rect 226064 234388 226116 234394
rect 226064 234330 226116 234336
rect 226260 231577 226288 239652
rect 226432 239634 226484 239640
rect 226338 239456 226394 239465
rect 226338 239391 226394 239400
rect 226352 238105 226380 239391
rect 226444 239329 226472 239634
rect 226430 239320 226486 239329
rect 226430 239255 226486 239264
rect 226536 239136 226564 239702
rect 226616 239488 226668 239494
rect 226616 239430 226668 239436
rect 226628 239290 226656 239430
rect 226616 239284 226668 239290
rect 226616 239226 226668 239232
rect 226536 239108 226656 239136
rect 226522 239048 226578 239057
rect 226522 238983 226578 238992
rect 226536 238542 226564 238983
rect 226524 238536 226576 238542
rect 226524 238478 226576 238484
rect 226628 238456 226656 239108
rect 226720 238746 226748 239720
rect 226800 239702 226852 239708
rect 226890 239728 226946 239737
rect 226812 239465 226840 239702
rect 226890 239663 226946 239672
rect 226798 239456 226854 239465
rect 226798 239391 226854 239400
rect 226708 238740 226760 238746
rect 226708 238682 226760 238688
rect 226628 238428 226748 238456
rect 226524 238400 226576 238406
rect 226524 238342 226576 238348
rect 226338 238096 226394 238105
rect 226338 238031 226394 238040
rect 226246 231568 226302 231577
rect 226246 231503 226302 231512
rect 226352 231305 226380 238031
rect 226432 233232 226484 233238
rect 226432 233174 226484 233180
rect 226338 231296 226394 231305
rect 226338 231231 226394 231240
rect 225788 229900 225840 229906
rect 225788 229842 225840 229848
rect 225972 229900 226024 229906
rect 225972 229842 226024 229848
rect 225984 224954 226012 229842
rect 225800 224926 226012 224954
rect 225800 144226 225828 224926
rect 225880 224732 225932 224738
rect 225880 224674 225932 224680
rect 225788 144220 225840 144226
rect 225788 144162 225840 144168
rect 225892 141710 225920 224674
rect 225970 220688 226026 220697
rect 225970 220623 226026 220632
rect 226064 220652 226116 220658
rect 225880 141704 225932 141710
rect 225880 141646 225932 141652
rect 225984 140418 226012 220623
rect 226064 220594 226116 220600
rect 226076 220318 226104 220594
rect 226064 220312 226116 220318
rect 226064 220254 226116 220260
rect 226076 164898 226104 220254
rect 226064 164892 226116 164898
rect 226064 164834 226116 164840
rect 226338 145616 226394 145625
rect 226338 145551 226394 145560
rect 225972 140412 226024 140418
rect 225972 140354 226024 140360
rect 225696 139120 225748 139126
rect 225696 139062 225748 139068
rect 225604 3596 225656 3602
rect 225604 3538 225656 3544
rect 226352 480 226380 145551
rect 226444 138961 226472 233174
rect 226536 231169 226564 238342
rect 226720 231854 226748 238428
rect 226812 232490 226840 239391
rect 226800 232484 226852 232490
rect 226800 232426 226852 232432
rect 226720 231826 226840 231854
rect 226522 231160 226578 231169
rect 226522 231095 226578 231104
rect 226616 230988 226668 230994
rect 226616 230930 226668 230936
rect 226628 223038 226656 230930
rect 226616 223032 226668 223038
rect 226616 222974 226668 222980
rect 226812 216646 226840 231826
rect 226800 216640 226852 216646
rect 226800 216582 226852 216588
rect 226904 215218 226932 239663
rect 226996 238202 227024 239822
rect 227214 239838 227266 239844
rect 227120 239799 227176 239808
rect 227168 239760 227220 239766
rect 227166 239728 227168 239737
rect 227410 239748 227438 240108
rect 227220 239728 227222 239737
rect 227076 239692 227128 239698
rect 227166 239663 227222 239672
rect 227272 239720 227438 239748
rect 227502 239748 227530 240108
rect 227594 239873 227622 240108
rect 227686 239970 227714 240108
rect 227674 239964 227726 239970
rect 227674 239906 227726 239912
rect 227580 239864 227636 239873
rect 227778 239850 227806 240108
rect 227580 239799 227636 239808
rect 227732 239822 227806 239850
rect 227870 239850 227898 240108
rect 227962 239970 227990 240108
rect 228054 239970 228082 240108
rect 227950 239964 228002 239970
rect 227950 239906 228002 239912
rect 228042 239964 228094 239970
rect 228042 239906 228094 239912
rect 227994 239864 228050 239873
rect 227870 239822 227944 239850
rect 227628 239760 227680 239766
rect 227502 239720 227576 239748
rect 227076 239634 227128 239640
rect 226984 238196 227036 238202
rect 226984 238138 227036 238144
rect 226984 227248 227036 227254
rect 226984 227190 227036 227196
rect 226892 215212 226944 215218
rect 226892 215154 226944 215160
rect 226996 145382 227024 227190
rect 227088 226302 227116 239634
rect 227168 239284 227220 239290
rect 227168 239226 227220 239232
rect 227180 233238 227208 239226
rect 227272 238649 227300 239720
rect 227352 239624 227404 239630
rect 227352 239566 227404 239572
rect 227444 239624 227496 239630
rect 227444 239566 227496 239572
rect 227364 239329 227392 239566
rect 227456 239358 227484 239566
rect 227444 239352 227496 239358
rect 227350 239320 227406 239329
rect 227444 239294 227496 239300
rect 227350 239255 227406 239264
rect 227258 238640 227314 238649
rect 227258 238575 227314 238584
rect 227364 238406 227392 239255
rect 227352 238400 227404 238406
rect 227352 238342 227404 238348
rect 227444 238332 227496 238338
rect 227444 238274 227496 238280
rect 227350 236328 227406 236337
rect 227350 236263 227406 236272
rect 227168 233232 227220 233238
rect 227168 233174 227220 233180
rect 227364 231418 227392 236263
rect 227180 231390 227392 231418
rect 227076 226296 227128 226302
rect 227076 226238 227128 226244
rect 227076 221876 227128 221882
rect 227076 221818 227128 221824
rect 226984 145376 227036 145382
rect 226984 145318 227036 145324
rect 227088 141642 227116 221818
rect 227180 218006 227208 231390
rect 227352 231260 227404 231266
rect 227352 231202 227404 231208
rect 227258 226264 227314 226273
rect 227258 226199 227314 226208
rect 227168 218000 227220 218006
rect 227168 217942 227220 217948
rect 227168 216640 227220 216646
rect 227168 216582 227220 216588
rect 227076 141636 227128 141642
rect 227076 141578 227128 141584
rect 226430 138952 226486 138961
rect 226430 138887 226486 138896
rect 227180 138009 227208 216582
rect 227272 147121 227300 226199
rect 227364 158137 227392 231202
rect 227456 231033 227484 238274
rect 227442 231024 227498 231033
rect 227548 230994 227576 239720
rect 227628 239702 227680 239708
rect 227640 239465 227668 239702
rect 227626 239456 227682 239465
rect 227626 239391 227682 239400
rect 227442 230959 227498 230968
rect 227536 230988 227588 230994
rect 227536 230930 227588 230936
rect 227536 229152 227588 229158
rect 227536 229094 227588 229100
rect 227548 215294 227576 229094
rect 227640 218793 227668 239391
rect 227732 235210 227760 239822
rect 227812 239760 227864 239766
rect 227812 239702 227864 239708
rect 227824 238202 227852 239702
rect 227916 238270 227944 239822
rect 228146 239850 228174 240108
rect 228238 239902 228266 240108
rect 228330 239902 228358 240108
rect 227994 239799 227996 239808
rect 228048 239799 228050 239808
rect 228100 239822 228174 239850
rect 228226 239896 228278 239902
rect 228226 239838 228278 239844
rect 228318 239896 228370 239902
rect 228318 239838 228370 239844
rect 227996 239770 228048 239776
rect 227994 239728 228050 239737
rect 227994 239663 228050 239672
rect 228008 239426 228036 239663
rect 227996 239420 228048 239426
rect 227996 239362 228048 239368
rect 227996 239216 228048 239222
rect 227996 239158 228048 239164
rect 228008 238377 228036 239158
rect 228100 239018 228128 239822
rect 228238 239748 228266 239838
rect 228422 239748 228450 240108
rect 228514 239970 228542 240108
rect 228502 239964 228554 239970
rect 228502 239906 228554 239912
rect 228238 239720 228312 239748
rect 228180 239624 228232 239630
rect 228180 239566 228232 239572
rect 228088 239012 228140 239018
rect 228088 238954 228140 238960
rect 228086 238640 228142 238649
rect 228192 238626 228220 239566
rect 228142 238598 228220 238626
rect 228086 238575 228142 238584
rect 227994 238368 228050 238377
rect 227994 238303 228050 238312
rect 227904 238264 227956 238270
rect 227904 238206 227956 238212
rect 227812 238196 227864 238202
rect 227812 238138 227864 238144
rect 227720 235204 227772 235210
rect 227720 235146 227772 235152
rect 227824 234614 227852 238138
rect 227732 234586 227852 234614
rect 227732 231441 227760 234586
rect 227996 231872 228048 231878
rect 227996 231814 228048 231820
rect 227718 231432 227774 231441
rect 227718 231367 227774 231376
rect 227626 218784 227682 218793
rect 227626 218719 227682 218728
rect 227720 218000 227772 218006
rect 227720 217942 227772 217948
rect 227732 217394 227760 217942
rect 227720 217388 227772 217394
rect 227720 217330 227772 217336
rect 227456 215266 227576 215294
rect 227456 158302 227484 215266
rect 227444 158296 227496 158302
rect 227444 158238 227496 158244
rect 227350 158128 227406 158137
rect 227350 158063 227406 158072
rect 227258 147112 227314 147121
rect 227258 147047 227314 147056
rect 227732 139194 227760 217330
rect 228008 216510 228036 231814
rect 228100 224233 228128 238575
rect 228178 238504 228234 238513
rect 228178 238439 228234 238448
rect 228192 234394 228220 238439
rect 228180 234388 228232 234394
rect 228180 234330 228232 234336
rect 228284 229809 228312 239720
rect 228376 239720 228450 239748
rect 228606 239748 228634 240108
rect 228698 239902 228726 240108
rect 228686 239896 228738 239902
rect 228686 239838 228738 239844
rect 228790 239850 228818 240108
rect 228882 239970 228910 240108
rect 228870 239964 228922 239970
rect 228870 239906 228922 239912
rect 228974 239873 229002 240108
rect 228960 239864 229016 239873
rect 228790 239822 228864 239850
rect 228836 239748 228864 239822
rect 229066 239850 229094 240108
rect 229158 239970 229186 240108
rect 229250 239970 229278 240108
rect 229342 239970 229370 240108
rect 229434 239970 229462 240108
rect 229146 239964 229198 239970
rect 229146 239906 229198 239912
rect 229238 239964 229290 239970
rect 229238 239906 229290 239912
rect 229330 239964 229382 239970
rect 229330 239906 229382 239912
rect 229422 239964 229474 239970
rect 229422 239906 229474 239912
rect 229526 239850 229554 240108
rect 229066 239822 229140 239850
rect 228960 239799 229016 239808
rect 229112 239748 229140 239822
rect 229376 239828 229428 239834
rect 229376 239770 229428 239776
rect 229480 239822 229554 239850
rect 228606 239720 228680 239748
rect 228744 239737 228864 239748
rect 228376 238762 228404 239720
rect 228456 239624 228508 239630
rect 228456 239566 228508 239572
rect 228548 239624 228600 239630
rect 228548 239566 228600 239572
rect 228468 238921 228496 239566
rect 228560 239290 228588 239566
rect 228548 239284 228600 239290
rect 228548 239226 228600 239232
rect 228454 238912 228510 238921
rect 228454 238847 228510 238856
rect 228376 238734 228588 238762
rect 228456 238400 228508 238406
rect 228456 238342 228508 238348
rect 228468 237289 228496 238342
rect 228454 237280 228510 237289
rect 228454 237215 228510 237224
rect 228456 234388 228508 234394
rect 228456 234330 228508 234336
rect 228364 229832 228416 229838
rect 228270 229800 228326 229809
rect 228364 229774 228416 229780
rect 228270 229735 228326 229744
rect 228180 227520 228232 227526
rect 228180 227462 228232 227468
rect 228086 224224 228142 224233
rect 228086 224159 228142 224168
rect 227996 216504 228048 216510
rect 227996 216446 228048 216452
rect 228192 215286 228220 227462
rect 228180 215280 228232 215286
rect 228180 215222 228232 215228
rect 228376 159390 228404 229774
rect 228468 220289 228496 234330
rect 228560 224954 228588 238734
rect 228652 227526 228680 239720
rect 228730 239728 228864 239737
rect 228786 239720 228864 239728
rect 229020 239720 229140 239748
rect 228730 239663 228786 239672
rect 228732 239624 228784 239630
rect 228732 239566 228784 239572
rect 228824 239624 228876 239630
rect 228824 239566 228876 239572
rect 228744 239465 228772 239566
rect 228730 239456 228786 239465
rect 228730 239391 228786 239400
rect 228836 239154 228864 239566
rect 228824 239148 228876 239154
rect 228824 239090 228876 239096
rect 228730 238912 228786 238921
rect 228730 238847 228786 238856
rect 228744 229838 228772 238847
rect 228824 238536 228876 238542
rect 229020 238513 229048 239720
rect 229284 239624 229336 239630
rect 229284 239566 229336 239572
rect 229100 239556 229152 239562
rect 229100 239498 229152 239504
rect 228824 238478 228876 238484
rect 229006 238504 229062 238513
rect 228836 231849 228864 238478
rect 229006 238439 229062 238448
rect 229112 238406 229140 239498
rect 229296 239290 229324 239566
rect 229284 239284 229336 239290
rect 229284 239226 229336 239232
rect 229282 239184 229338 239193
rect 229282 239119 229338 239128
rect 229100 238400 229152 238406
rect 229100 238342 229152 238348
rect 229192 238264 229244 238270
rect 229192 238206 229244 238212
rect 229100 237856 229152 237862
rect 229100 237798 229152 237804
rect 229112 237697 229140 237798
rect 229098 237688 229154 237697
rect 229098 237623 229154 237632
rect 228822 231840 228878 231849
rect 228822 231775 228878 231784
rect 229006 231296 229062 231305
rect 229006 231231 229062 231240
rect 228916 230444 228968 230450
rect 228916 230386 228968 230392
rect 228732 229832 228784 229838
rect 228732 229774 228784 229780
rect 228640 227520 228692 227526
rect 228640 227462 228692 227468
rect 228560 224926 228680 224954
rect 228546 224224 228602 224233
rect 228546 224159 228602 224168
rect 228454 220280 228510 220289
rect 228454 220215 228510 220224
rect 228456 216640 228508 216646
rect 228456 216582 228508 216588
rect 228468 216442 228496 216582
rect 228456 216436 228508 216442
rect 228456 216378 228508 216384
rect 228364 159384 228416 159390
rect 228364 159326 228416 159332
rect 227812 154148 227864 154154
rect 227812 154090 227864 154096
rect 227824 153270 227852 154090
rect 228364 154012 228416 154018
rect 228364 153954 228416 153960
rect 227812 153264 227864 153270
rect 227812 153206 227864 153212
rect 227720 139188 227772 139194
rect 227720 139130 227772 139136
rect 227166 138000 227222 138009
rect 227166 137935 227222 137944
rect 226430 130384 226486 130393
rect 226430 130319 226486 130328
rect 226444 16574 226472 130319
rect 226444 16546 227576 16574
rect 227548 480 227576 16546
rect 228376 3738 228404 153954
rect 228468 139058 228496 216378
rect 228560 147626 228588 224159
rect 228652 216646 228680 224926
rect 228640 216640 228692 216646
rect 228640 216582 228692 216588
rect 228732 216640 228784 216646
rect 228732 216582 228784 216588
rect 228640 216504 228692 216510
rect 228640 216446 228692 216452
rect 228652 216374 228680 216446
rect 228640 216368 228692 216374
rect 228640 216310 228692 216316
rect 228548 147620 228600 147626
rect 228548 147562 228600 147568
rect 228652 144537 228680 216310
rect 228744 216306 228772 216582
rect 228732 216300 228784 216306
rect 228732 216242 228784 216248
rect 228928 153270 228956 230386
rect 228916 153264 228968 153270
rect 228916 153206 228968 153212
rect 228638 144528 228694 144537
rect 228638 144463 228694 144472
rect 228456 139052 228508 139058
rect 228456 138994 228508 139000
rect 229020 124137 229048 231231
rect 229204 159050 229232 238206
rect 229296 217025 229324 239119
rect 229388 237454 229416 239770
rect 229376 237448 229428 237454
rect 229376 237390 229428 237396
rect 229480 231946 229508 239822
rect 229618 239748 229646 240108
rect 229710 239873 229738 240108
rect 229802 239902 229830 240108
rect 229894 239970 229922 240108
rect 229882 239964 229934 239970
rect 229882 239906 229934 239912
rect 229790 239896 229842 239902
rect 229696 239864 229752 239873
rect 229986 239850 230014 240108
rect 230078 239970 230106 240108
rect 230066 239964 230118 239970
rect 230066 239906 230118 239912
rect 229790 239838 229842 239844
rect 229696 239799 229752 239808
rect 229940 239822 230014 239850
rect 229572 239720 229646 239748
rect 229836 239760 229888 239766
rect 229572 237561 229600 239720
rect 229836 239702 229888 239708
rect 229652 239624 229704 239630
rect 229652 239566 229704 239572
rect 229664 239465 229692 239566
rect 229744 239488 229796 239494
rect 229650 239456 229706 239465
rect 229744 239430 229796 239436
rect 229650 239391 229706 239400
rect 229664 238270 229692 239391
rect 229756 239018 229784 239430
rect 229744 239012 229796 239018
rect 229744 238954 229796 238960
rect 229848 238649 229876 239702
rect 229834 238640 229890 238649
rect 229834 238575 229890 238584
rect 229848 238338 229876 238575
rect 229836 238332 229888 238338
rect 229836 238274 229888 238280
rect 229652 238264 229704 238270
rect 229652 238206 229704 238212
rect 229940 237912 229968 239822
rect 230020 239760 230072 239766
rect 230170 239737 230198 240108
rect 230262 239748 230290 240108
rect 230354 239873 230382 240108
rect 230340 239864 230396 239873
rect 230446 239850 230474 240108
rect 230538 239970 230566 240108
rect 230526 239964 230578 239970
rect 230526 239906 230578 239912
rect 230630 239873 230658 240108
rect 230616 239864 230672 239873
rect 230446 239822 230566 239850
rect 230340 239799 230396 239808
rect 230538 239748 230566 239822
rect 230616 239799 230672 239808
rect 230020 239702 230072 239708
rect 230156 239728 230212 239737
rect 230032 238746 230060 239702
rect 230262 239720 230336 239748
rect 230156 239663 230212 239672
rect 230112 239420 230164 239426
rect 230112 239362 230164 239368
rect 230124 239193 230152 239362
rect 230110 239184 230166 239193
rect 230166 239142 230244 239170
rect 230110 239119 230166 239128
rect 230020 238740 230072 238746
rect 230020 238682 230072 238688
rect 230216 238474 230244 239142
rect 230204 238468 230256 238474
rect 230204 238410 230256 238416
rect 229664 237884 229968 237912
rect 229558 237552 229614 237561
rect 229558 237487 229614 237496
rect 229560 237448 229612 237454
rect 229560 237390 229612 237396
rect 229468 231940 229520 231946
rect 229468 231882 229520 231888
rect 229572 229945 229600 237390
rect 229664 231810 229692 237884
rect 229928 237788 229980 237794
rect 229928 237730 229980 237736
rect 229940 237454 229968 237730
rect 229928 237448 229980 237454
rect 229928 237390 229980 237396
rect 229834 235648 229890 235657
rect 229834 235583 229890 235592
rect 229744 235408 229796 235414
rect 229744 235350 229796 235356
rect 229652 231804 229704 231810
rect 229652 231746 229704 231752
rect 229558 229936 229614 229945
rect 229558 229871 229614 229880
rect 229650 217968 229706 217977
rect 229650 217903 229706 217912
rect 229664 217705 229692 217903
rect 229650 217696 229706 217705
rect 229650 217631 229706 217640
rect 229282 217016 229338 217025
rect 229282 216951 229338 216960
rect 229756 160954 229784 235350
rect 229744 160948 229796 160954
rect 229744 160890 229796 160896
rect 229192 159044 229244 159050
rect 229192 158986 229244 158992
rect 229744 153264 229796 153270
rect 229744 153206 229796 153212
rect 229100 151360 229152 151366
rect 229100 151302 229152 151308
rect 229006 124128 229062 124137
rect 229006 124063 229062 124072
rect 229020 122913 229048 124063
rect 229006 122904 229062 122913
rect 229006 122839 229062 122848
rect 229112 16574 229140 151302
rect 229112 16546 229416 16574
rect 228364 3732 228416 3738
rect 228364 3674 228416 3680
rect 228732 3596 228784 3602
rect 228732 3538 228784 3544
rect 228744 480 228772 3538
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 229756 3126 229784 153206
rect 229848 142934 229876 235583
rect 230020 230376 230072 230382
rect 230020 230318 230072 230324
rect 229926 220280 229982 220289
rect 229926 220215 229982 220224
rect 229836 142928 229888 142934
rect 229836 142870 229888 142876
rect 229940 140049 229968 220215
rect 230032 151366 230060 230318
rect 230308 229090 230336 239720
rect 230400 239720 230566 239748
rect 230722 239748 230750 240108
rect 230814 239902 230842 240108
rect 230802 239896 230854 239902
rect 230906 239873 230934 240108
rect 230998 239970 231026 240108
rect 230986 239964 231038 239970
rect 230986 239906 231038 239912
rect 230802 239838 230854 239844
rect 230892 239864 230948 239873
rect 231090 239850 231118 240108
rect 230892 239799 230948 239808
rect 231044 239822 231118 239850
rect 231182 239850 231210 240108
rect 231274 239970 231302 240108
rect 231262 239964 231314 239970
rect 231262 239906 231314 239912
rect 231366 239850 231394 240108
rect 231458 239902 231486 240108
rect 231182 239822 231256 239850
rect 230722 239720 230888 239748
rect 230400 238338 230428 239720
rect 230664 239624 230716 239630
rect 230492 239584 230664 239612
rect 230492 238626 230520 239584
rect 230664 239566 230716 239572
rect 230756 239624 230808 239630
rect 230756 239566 230808 239572
rect 230664 239420 230716 239426
rect 230664 239362 230716 239368
rect 230676 238950 230704 239362
rect 230664 238944 230716 238950
rect 230664 238886 230716 238892
rect 230662 238640 230718 238649
rect 230492 238598 230612 238626
rect 230388 238332 230440 238338
rect 230388 238274 230440 238280
rect 230400 235414 230428 238274
rect 230584 237522 230612 238598
rect 230662 238575 230718 238584
rect 230676 238474 230704 238575
rect 230664 238468 230716 238474
rect 230664 238410 230716 238416
rect 230572 237516 230624 237522
rect 230572 237458 230624 237464
rect 230478 237416 230534 237425
rect 230478 237351 230534 237360
rect 230388 235408 230440 235414
rect 230388 235350 230440 235356
rect 230388 231940 230440 231946
rect 230388 231882 230440 231888
rect 230296 229084 230348 229090
rect 230296 229026 230348 229032
rect 230204 224188 230256 224194
rect 230204 224130 230256 224136
rect 230112 221808 230164 221814
rect 230112 221750 230164 221756
rect 230124 160585 230152 221750
rect 230216 214577 230244 224130
rect 230400 217977 230428 231882
rect 230386 217968 230442 217977
rect 230386 217903 230442 217912
rect 230492 217161 230520 237351
rect 230584 229022 230612 237458
rect 230572 229016 230624 229022
rect 230572 228958 230624 228964
rect 230676 224194 230704 238410
rect 230768 231878 230796 239566
rect 230860 238950 230888 239720
rect 230938 239728 230994 239737
rect 230938 239663 230994 239672
rect 230848 238944 230900 238950
rect 230848 238886 230900 238892
rect 230756 231872 230808 231878
rect 230756 231814 230808 231820
rect 230846 231840 230902 231849
rect 230846 231775 230902 231784
rect 230756 231736 230808 231742
rect 230756 231678 230808 231684
rect 230664 224188 230716 224194
rect 230664 224130 230716 224136
rect 230572 218068 230624 218074
rect 230572 218010 230624 218016
rect 230478 217152 230534 217161
rect 230478 217087 230534 217096
rect 230584 216306 230612 218010
rect 230572 216300 230624 216306
rect 230572 216242 230624 216248
rect 230202 214568 230258 214577
rect 230202 214503 230258 214512
rect 230204 184204 230256 184210
rect 230204 184146 230256 184152
rect 230110 160576 230166 160585
rect 230110 160511 230166 160520
rect 230020 151360 230072 151366
rect 230020 151302 230072 151308
rect 230216 148306 230244 184146
rect 230768 160886 230796 231678
rect 230860 217841 230888 231775
rect 230952 231742 230980 239663
rect 231044 238377 231072 239822
rect 231124 239760 231176 239766
rect 231122 239728 231124 239737
rect 231176 239728 231178 239737
rect 231122 239663 231178 239672
rect 231124 239624 231176 239630
rect 231124 239566 231176 239572
rect 231030 238368 231086 238377
rect 231030 238303 231086 238312
rect 231136 237538 231164 239566
rect 231228 239465 231256 239822
rect 231320 239822 231394 239850
rect 231446 239896 231498 239902
rect 231446 239838 231498 239844
rect 231214 239456 231270 239465
rect 231320 239442 231348 239822
rect 231550 239748 231578 240108
rect 231642 239850 231670 240108
rect 231734 239970 231762 240108
rect 231722 239964 231774 239970
rect 231722 239906 231774 239912
rect 231826 239850 231854 240108
rect 231918 239902 231946 240108
rect 231642 239822 231716 239850
rect 231398 239728 231454 239737
rect 231550 239720 231624 239748
rect 231398 239663 231400 239672
rect 231452 239663 231454 239672
rect 231400 239634 231452 239640
rect 231320 239414 231440 239442
rect 231214 239391 231270 239400
rect 231228 238542 231256 239391
rect 231308 239284 231360 239290
rect 231308 239226 231360 239232
rect 231320 238649 231348 239226
rect 231306 238640 231362 238649
rect 231306 238575 231362 238584
rect 231216 238536 231268 238542
rect 231216 238478 231268 238484
rect 231214 237552 231270 237561
rect 231136 237510 231214 237538
rect 231214 237487 231270 237496
rect 231228 233918 231256 237487
rect 231308 237448 231360 237454
rect 231308 237390 231360 237396
rect 231216 233912 231268 233918
rect 231216 233854 231268 233860
rect 230940 231736 230992 231742
rect 230940 231678 230992 231684
rect 231320 229094 231348 237390
rect 231412 234614 231440 239414
rect 231492 238944 231544 238950
rect 231492 238886 231544 238892
rect 231504 238270 231532 238886
rect 231492 238264 231544 238270
rect 231492 238206 231544 238212
rect 231504 237454 231532 238206
rect 231596 237969 231624 239720
rect 231688 239544 231716 239822
rect 231780 239822 231854 239850
rect 231906 239896 231958 239902
rect 232010 239873 232038 240108
rect 231906 239838 231958 239844
rect 231996 239864 232052 239873
rect 231780 239612 231808 239822
rect 231996 239799 232052 239808
rect 231860 239760 231912 239766
rect 231858 239728 231860 239737
rect 232102 239748 232130 240108
rect 232194 239850 232222 240108
rect 232286 239970 232314 240108
rect 232274 239964 232326 239970
rect 232274 239906 232326 239912
rect 232194 239822 232268 239850
rect 231912 239728 231914 239737
rect 232102 239720 232176 239748
rect 231858 239663 231914 239672
rect 231780 239584 231900 239612
rect 231688 239516 231808 239544
rect 231676 239284 231728 239290
rect 231676 239226 231728 239232
rect 231688 239154 231716 239226
rect 231676 239148 231728 239154
rect 231676 239090 231728 239096
rect 231780 238134 231808 239516
rect 231872 238610 231900 239584
rect 231952 239556 232004 239562
rect 231952 239498 232004 239504
rect 231964 239465 231992 239498
rect 231950 239456 232006 239465
rect 231950 239391 232006 239400
rect 232042 239184 232098 239193
rect 232042 239119 232098 239128
rect 231860 238604 231912 238610
rect 231860 238546 231912 238552
rect 231676 238128 231728 238134
rect 231674 238096 231676 238105
rect 231768 238128 231820 238134
rect 231728 238096 231730 238105
rect 231768 238070 231820 238076
rect 231674 238031 231730 238040
rect 231582 237960 231638 237969
rect 231638 237918 231716 237946
rect 231582 237895 231638 237904
rect 231596 237835 231624 237895
rect 231688 237590 231716 237918
rect 231584 237584 231636 237590
rect 231584 237526 231636 237532
rect 231676 237584 231728 237590
rect 231676 237526 231728 237532
rect 231596 237454 231624 237526
rect 231492 237448 231544 237454
rect 231492 237390 231544 237396
rect 231584 237448 231636 237454
rect 231584 237390 231636 237396
rect 231780 237374 231808 238070
rect 231872 237726 231900 238546
rect 231952 238400 232004 238406
rect 231952 238342 232004 238348
rect 231964 238202 231992 238342
rect 231952 238196 232004 238202
rect 231952 238138 232004 238144
rect 231860 237720 231912 237726
rect 231860 237662 231912 237668
rect 231688 237346 231808 237374
rect 231952 237380 232004 237386
rect 231412 234586 231532 234614
rect 231320 229066 231440 229094
rect 231308 229016 231360 229022
rect 231308 228958 231360 228964
rect 231124 228948 231176 228954
rect 231124 228890 231176 228896
rect 230846 217832 230902 217841
rect 230846 217767 230902 217776
rect 230756 160880 230808 160886
rect 230756 160822 230808 160828
rect 230204 148300 230256 148306
rect 230204 148242 230256 148248
rect 231136 144294 231164 228890
rect 231214 221776 231270 221785
rect 231214 221711 231270 221720
rect 231124 144288 231176 144294
rect 231124 144230 231176 144236
rect 231228 140486 231256 221711
rect 231320 188329 231348 228958
rect 231412 217433 231440 229066
rect 231504 218074 231532 234586
rect 231688 232626 231716 237346
rect 231952 237322 232004 237328
rect 231964 236706 231992 237322
rect 231952 236700 232004 236706
rect 231952 236642 232004 236648
rect 231858 234152 231914 234161
rect 231858 234087 231914 234096
rect 231872 233306 231900 234087
rect 231860 233300 231912 233306
rect 231860 233242 231912 233248
rect 231676 232620 231728 232626
rect 231676 232562 231728 232568
rect 232056 223574 232084 239119
rect 232148 238542 232176 239720
rect 232240 239358 232268 239822
rect 232378 239816 232406 240108
rect 232470 239970 232498 240108
rect 232458 239964 232510 239970
rect 232458 239906 232510 239912
rect 232562 239816 232590 240108
rect 232654 239970 232682 240108
rect 232642 239964 232694 239970
rect 232642 239906 232694 239912
rect 232746 239850 232774 240108
rect 232332 239788 232406 239816
rect 232516 239788 232590 239816
rect 232700 239822 232774 239850
rect 232838 239850 232866 240108
rect 232930 239970 232958 240108
rect 232918 239964 232970 239970
rect 232918 239906 232970 239912
rect 232838 239822 232912 239850
rect 232228 239352 232280 239358
rect 232228 239294 232280 239300
rect 232136 238536 232188 238542
rect 232136 238478 232188 238484
rect 232240 237386 232268 239294
rect 232332 237998 232360 239788
rect 232412 239692 232464 239698
rect 232412 239634 232464 239640
rect 232424 238950 232452 239634
rect 232412 238944 232464 238950
rect 232412 238886 232464 238892
rect 232424 238678 232452 238886
rect 232412 238672 232464 238678
rect 232412 238614 232464 238620
rect 232320 237992 232372 237998
rect 232320 237934 232372 237940
rect 232228 237380 232280 237386
rect 232228 237322 232280 237328
rect 232516 236978 232544 239788
rect 232596 239692 232648 239698
rect 232596 239634 232648 239640
rect 232504 236972 232556 236978
rect 232504 236914 232556 236920
rect 232608 232914 232636 239634
rect 232700 238377 232728 239822
rect 232884 239748 232912 239822
rect 233022 239748 233050 240108
rect 232792 239720 232912 239748
rect 232976 239720 233050 239748
rect 233114 239748 233142 240108
rect 233206 239873 233234 240108
rect 233298 239902 233326 240108
rect 233390 239970 233418 240108
rect 233482 239970 233510 240108
rect 233574 239970 233602 240108
rect 233666 239970 233694 240108
rect 233758 239970 233786 240108
rect 233850 239970 233878 240108
rect 233942 239970 233970 240108
rect 233378 239964 233430 239970
rect 233378 239906 233430 239912
rect 233470 239964 233522 239970
rect 233470 239906 233522 239912
rect 233562 239964 233614 239970
rect 233562 239906 233614 239912
rect 233654 239964 233706 239970
rect 233654 239906 233706 239912
rect 233746 239964 233798 239970
rect 233746 239906 233798 239912
rect 233838 239964 233890 239970
rect 233838 239906 233890 239912
rect 233930 239964 233982 239970
rect 233930 239906 233982 239912
rect 233286 239896 233338 239902
rect 233192 239864 233248 239873
rect 233286 239838 233338 239844
rect 233514 239864 233570 239873
rect 233192 239799 233248 239808
rect 233424 239828 233476 239834
rect 233514 239799 233516 239808
rect 233424 239770 233476 239776
rect 233568 239799 233570 239808
rect 233790 239864 233846 239873
rect 234034 239850 234062 240108
rect 233790 239799 233792 239808
rect 233516 239770 233568 239776
rect 233844 239799 233846 239808
rect 233884 239828 233936 239834
rect 233792 239770 233844 239776
rect 233884 239770 233936 239776
rect 233988 239822 234062 239850
rect 233332 239760 233384 239766
rect 233114 239720 233188 239748
rect 232792 239494 232820 239720
rect 232780 239488 232832 239494
rect 232780 239430 232832 239436
rect 232872 239488 232924 239494
rect 232872 239430 232924 239436
rect 232792 238610 232820 239430
rect 232780 238604 232832 238610
rect 232780 238546 232832 238552
rect 232884 238490 232912 239430
rect 232792 238462 232912 238490
rect 232686 238368 232742 238377
rect 232686 238303 232742 238312
rect 232688 236972 232740 236978
rect 232688 236914 232740 236920
rect 231964 223546 232084 223574
rect 232332 232886 232636 232914
rect 231860 219428 231912 219434
rect 231860 219370 231912 219376
rect 231872 218754 231900 219370
rect 231860 218748 231912 218754
rect 231860 218690 231912 218696
rect 231492 218068 231544 218074
rect 231492 218010 231544 218016
rect 231964 217569 231992 223546
rect 232332 219434 232360 232886
rect 232504 232756 232556 232762
rect 232504 232698 232556 232704
rect 232320 219428 232372 219434
rect 232320 219370 232372 219376
rect 231950 217560 232006 217569
rect 231950 217495 232006 217504
rect 231398 217424 231454 217433
rect 231398 217359 231454 217368
rect 231306 188320 231362 188329
rect 231306 188255 231362 188264
rect 232516 151434 232544 232698
rect 232596 230988 232648 230994
rect 232596 230930 232648 230936
rect 232504 151428 232556 151434
rect 232504 151370 232556 151376
rect 231216 140480 231268 140486
rect 231216 140422 231268 140428
rect 229926 140040 229982 140049
rect 229926 139975 229982 139984
rect 230478 122904 230534 122913
rect 230478 122839 230534 122848
rect 230492 16574 230520 122839
rect 230492 16546 231072 16574
rect 229744 3120 229796 3126
rect 229744 3062 229796 3068
rect 231044 480 231072 16546
rect 232516 3670 232544 151370
rect 232608 147257 232636 230930
rect 232700 228342 232728 236914
rect 232688 228336 232740 228342
rect 232688 228278 232740 228284
rect 232594 147248 232650 147257
rect 232594 147183 232650 147192
rect 232700 143177 232728 228278
rect 232792 226273 232820 238462
rect 232872 234796 232924 234802
rect 232872 234738 232924 234744
rect 232778 226264 232834 226273
rect 232778 226199 232834 226208
rect 232884 224466 232912 234738
rect 232976 229906 233004 239720
rect 233160 239680 233188 239720
rect 233068 239652 233188 239680
rect 233238 239728 233294 239737
rect 233332 239702 233384 239708
rect 233238 239663 233240 239672
rect 233068 239494 233096 239652
rect 233292 239663 233294 239672
rect 233240 239634 233292 239640
rect 233240 239556 233292 239562
rect 233240 239498 233292 239504
rect 233056 239488 233108 239494
rect 233148 239488 233200 239494
rect 233056 239430 233108 239436
rect 233146 239456 233148 239465
rect 233200 239456 233202 239465
rect 233146 239391 233202 239400
rect 233056 239148 233108 239154
rect 233056 239090 233108 239096
rect 233068 238814 233096 239090
rect 233252 238814 233280 239498
rect 233344 239329 233372 239702
rect 233436 239562 233464 239770
rect 233424 239556 233476 239562
rect 233424 239498 233476 239504
rect 233330 239320 233386 239329
rect 233330 239255 233386 239264
rect 233528 239170 233556 239770
rect 233700 239760 233752 239766
rect 233606 239728 233662 239737
rect 233700 239702 233752 239708
rect 233606 239663 233662 239672
rect 233344 239142 233556 239170
rect 233056 238808 233108 238814
rect 233240 238808 233292 238814
rect 233056 238750 233108 238756
rect 233160 238756 233240 238762
rect 233160 238750 233292 238756
rect 233160 238734 233280 238750
rect 233056 238536 233108 238542
rect 233056 238478 233108 238484
rect 233068 238202 233096 238478
rect 233056 238196 233108 238202
rect 233056 238138 233108 238144
rect 232964 229900 233016 229906
rect 232964 229842 233016 229848
rect 232872 224460 232924 224466
rect 232872 224402 232924 224408
rect 232780 220108 232832 220114
rect 232780 220050 232832 220056
rect 232686 143168 232742 143177
rect 232686 143103 232742 143112
rect 232792 141681 232820 220050
rect 232884 149734 232912 224402
rect 232976 156466 233004 229842
rect 233068 217297 233096 238138
rect 233160 235278 233188 238734
rect 233252 238685 233280 238734
rect 233240 238536 233292 238542
rect 233240 238478 233292 238484
rect 233252 238338 233280 238478
rect 233240 238332 233292 238338
rect 233240 238274 233292 238280
rect 233148 235272 233200 235278
rect 233148 235214 233200 235220
rect 233344 229022 233372 239142
rect 233516 238740 233568 238746
rect 233516 238682 233568 238688
rect 233424 238332 233476 238338
rect 233424 238274 233476 238280
rect 233436 237794 233464 238274
rect 233424 237788 233476 237794
rect 233424 237730 233476 237736
rect 233528 236609 233556 238682
rect 233514 236600 233570 236609
rect 233514 236535 233570 236544
rect 233620 230994 233648 239663
rect 233712 232490 233740 239702
rect 233804 238746 233832 239770
rect 233896 239737 233924 239770
rect 233882 239728 233938 239737
rect 233882 239663 233938 239672
rect 233988 239329 234016 239822
rect 234126 239748 234154 240108
rect 234218 239970 234246 240108
rect 234310 239970 234338 240108
rect 234206 239964 234258 239970
rect 234206 239906 234258 239912
rect 234298 239964 234350 239970
rect 234298 239906 234350 239912
rect 234250 239864 234306 239873
rect 234250 239799 234252 239808
rect 234304 239799 234306 239808
rect 234252 239770 234304 239776
rect 234080 239720 234154 239748
rect 233974 239320 234030 239329
rect 233974 239255 234030 239264
rect 233792 238740 233844 238746
rect 233792 238682 233844 238688
rect 233988 237374 234016 239255
rect 233896 237346 234016 237374
rect 233790 235512 233846 235521
rect 233790 235447 233846 235456
rect 233700 232484 233752 232490
rect 233700 232426 233752 232432
rect 233608 230988 233660 230994
rect 233608 230930 233660 230936
rect 233804 229094 233832 235447
rect 233896 232665 233924 237346
rect 233976 236156 234028 236162
rect 233976 236098 234028 236104
rect 233882 232656 233938 232665
rect 233882 232591 233938 232600
rect 233804 229066 233924 229094
rect 233332 229016 233384 229022
rect 233332 228958 233384 228964
rect 233792 229016 233844 229022
rect 233792 228958 233844 228964
rect 233700 228268 233752 228274
rect 233700 228210 233752 228216
rect 233712 221678 233740 228210
rect 233700 221672 233752 221678
rect 233700 221614 233752 221620
rect 233804 221513 233832 228958
rect 233790 221504 233846 221513
rect 233790 221439 233846 221448
rect 233054 217288 233110 217297
rect 233054 217223 233110 217232
rect 232964 156460 233016 156466
rect 232964 156402 233016 156408
rect 233240 151020 233292 151026
rect 233240 150962 233292 150968
rect 233252 150550 233280 150962
rect 233240 150544 233292 150550
rect 233240 150486 233292 150492
rect 232872 149728 232924 149734
rect 232872 149670 232924 149676
rect 232778 141672 232834 141681
rect 232778 141607 232834 141616
rect 233252 16574 233280 150486
rect 233896 126993 233924 229066
rect 233988 151298 234016 236098
rect 234080 231402 234108 239720
rect 234264 239630 234292 239770
rect 234402 239748 234430 240108
rect 234494 239907 234522 240108
rect 234480 239898 234536 239907
rect 234586 239902 234614 240108
rect 234480 239833 234536 239842
rect 234574 239896 234626 239902
rect 234574 239838 234626 239844
rect 234678 239850 234706 240108
rect 234770 239970 234798 240108
rect 234862 239970 234890 240108
rect 234758 239964 234810 239970
rect 234758 239906 234810 239912
rect 234850 239964 234902 239970
rect 234850 239906 234902 239912
rect 234678 239822 234752 239850
rect 234620 239760 234672 239766
rect 234402 239720 234568 239748
rect 234252 239624 234304 239630
rect 234252 239566 234304 239572
rect 234436 239624 234488 239630
rect 234436 239566 234488 239572
rect 234344 239488 234396 239494
rect 234344 239430 234396 239436
rect 234250 239320 234306 239329
rect 234250 239255 234306 239264
rect 234264 237374 234292 239255
rect 234172 237346 234292 237374
rect 234068 231396 234120 231402
rect 234068 231338 234120 231344
rect 234066 231160 234122 231169
rect 234066 231095 234122 231104
rect 233976 151292 234028 151298
rect 233976 151234 234028 151240
rect 234080 149802 234108 231095
rect 234172 228274 234200 237346
rect 234252 232484 234304 232490
rect 234252 232426 234304 232432
rect 234160 228268 234212 228274
rect 234160 228210 234212 228216
rect 234264 228154 234292 232426
rect 234172 228126 234292 228154
rect 234172 224806 234200 228126
rect 234356 227118 234384 239430
rect 234448 232801 234476 239566
rect 234540 239494 234568 239720
rect 234618 239728 234620 239737
rect 234672 239728 234674 239737
rect 234618 239663 234674 239672
rect 234620 239624 234672 239630
rect 234620 239566 234672 239572
rect 234528 239488 234580 239494
rect 234632 239465 234660 239566
rect 234528 239430 234580 239436
rect 234618 239456 234674 239465
rect 234618 239391 234674 239400
rect 234724 239086 234752 239822
rect 234862 239816 234890 239906
rect 234816 239788 234890 239816
rect 234712 239080 234764 239086
rect 234712 239022 234764 239028
rect 234816 238932 234844 239788
rect 234954 239748 234982 240108
rect 235046 239970 235074 240108
rect 235034 239964 235086 239970
rect 235034 239906 235086 239912
rect 235138 239850 235166 240108
rect 234632 238904 234844 238932
rect 234908 239720 234982 239748
rect 235092 239822 235166 239850
rect 234434 232792 234490 232801
rect 234434 232727 234490 232736
rect 234632 232558 234660 238904
rect 234908 237250 234936 239720
rect 234988 239148 235040 239154
rect 234988 239090 235040 239096
rect 235000 238950 235028 239090
rect 234988 238944 235040 238950
rect 234988 238886 235040 238892
rect 234988 238672 235040 238678
rect 234988 238614 235040 238620
rect 234896 237244 234948 237250
rect 234896 237186 234948 237192
rect 234804 237108 234856 237114
rect 234804 237050 234856 237056
rect 234712 235272 234764 235278
rect 234712 235214 234764 235220
rect 234620 232552 234672 232558
rect 234620 232494 234672 232500
rect 234528 231532 234580 231538
rect 234528 231474 234580 231480
rect 234436 231396 234488 231402
rect 234436 231338 234488 231344
rect 234448 228546 234476 231338
rect 234436 228540 234488 228546
rect 234436 228482 234488 228488
rect 234344 227112 234396 227118
rect 234344 227054 234396 227060
rect 234252 225684 234304 225690
rect 234252 225626 234304 225632
rect 234160 224800 234212 224806
rect 234160 224742 234212 224748
rect 234068 149796 234120 149802
rect 234068 149738 234120 149744
rect 234172 147529 234200 224742
rect 234264 150550 234292 225626
rect 234342 224904 234398 224913
rect 234342 224839 234398 224848
rect 234356 151201 234384 224839
rect 234448 155038 234476 228482
rect 234540 158642 234568 231474
rect 234724 227458 234752 235214
rect 234816 227798 234844 237050
rect 234908 234054 234936 237186
rect 235000 237153 235028 238614
rect 234986 237144 235042 237153
rect 234986 237079 235042 237088
rect 234896 234048 234948 234054
rect 234896 233990 234948 233996
rect 235092 229094 235120 239822
rect 235230 239748 235258 240108
rect 235322 239850 235350 240108
rect 235414 239970 235442 240108
rect 235402 239964 235454 239970
rect 235402 239906 235454 239912
rect 235506 239850 235534 240108
rect 235598 239970 235626 240108
rect 235690 239970 235718 240108
rect 235586 239964 235638 239970
rect 235586 239906 235638 239912
rect 235678 239964 235730 239970
rect 235678 239906 235730 239912
rect 235782 239850 235810 240108
rect 235874 239902 235902 240108
rect 235322 239822 235396 239850
rect 235506 239822 235580 239850
rect 235184 239720 235258 239748
rect 235184 237658 235212 239720
rect 235264 239624 235316 239630
rect 235264 239566 235316 239572
rect 235276 239465 235304 239566
rect 235262 239456 235318 239465
rect 235262 239391 235318 239400
rect 235172 237652 235224 237658
rect 235172 237594 235224 237600
rect 235368 236065 235396 239822
rect 235448 239760 235500 239766
rect 235448 239702 235500 239708
rect 235460 236337 235488 239702
rect 235446 236328 235502 236337
rect 235446 236263 235502 236272
rect 235354 236056 235410 236065
rect 235354 235991 235410 236000
rect 235552 232830 235580 239822
rect 235736 239822 235810 239850
rect 235862 239896 235914 239902
rect 235862 239838 235914 239844
rect 235966 239850 235994 240108
rect 236058 239970 236086 240108
rect 236046 239964 236098 239970
rect 236046 239906 236098 239912
rect 236150 239850 236178 240108
rect 235966 239822 236040 239850
rect 235632 239760 235684 239766
rect 235632 239702 235684 239708
rect 235644 237114 235672 239702
rect 235736 237862 235764 239822
rect 235908 239760 235960 239766
rect 235908 239702 235960 239708
rect 235816 239488 235868 239494
rect 235816 239430 235868 239436
rect 235724 237856 235776 237862
rect 235724 237798 235776 237804
rect 235828 237374 235856 239430
rect 235736 237346 235856 237374
rect 235632 237108 235684 237114
rect 235632 237050 235684 237056
rect 235632 236972 235684 236978
rect 235632 236914 235684 236920
rect 235540 232824 235592 232830
rect 235540 232766 235592 232772
rect 235552 232370 235580 232766
rect 235000 229066 235120 229094
rect 235184 232342 235580 232370
rect 234804 227792 234856 227798
rect 234804 227734 234856 227740
rect 234712 227452 234764 227458
rect 234712 227394 234764 227400
rect 234724 226574 234752 227394
rect 234712 226568 234764 226574
rect 234712 226510 234764 226516
rect 235000 221610 235028 229066
rect 234988 221604 235040 221610
rect 234988 221546 235040 221552
rect 235000 213217 235028 221546
rect 234986 213208 235042 213217
rect 234986 213143 235042 213152
rect 234528 158636 234580 158642
rect 234528 158578 234580 158584
rect 235184 156398 235212 232342
rect 235264 229696 235316 229702
rect 235264 229638 235316 229644
rect 235172 156392 235224 156398
rect 235172 156334 235224 156340
rect 234436 155032 234488 155038
rect 234436 154974 234488 154980
rect 234342 151192 234398 151201
rect 234342 151127 234398 151136
rect 234252 150544 234304 150550
rect 234252 150486 234304 150492
rect 235276 149938 235304 229638
rect 235540 228268 235592 228274
rect 235540 228210 235592 228216
rect 235552 227798 235580 228210
rect 235540 227792 235592 227798
rect 235540 227734 235592 227740
rect 235448 226568 235500 226574
rect 235448 226510 235500 226516
rect 235354 220416 235410 220425
rect 235354 220351 235410 220360
rect 235264 149932 235316 149938
rect 235264 149874 235316 149880
rect 234158 147520 234214 147529
rect 234158 147455 234214 147464
rect 233882 126984 233938 126993
rect 233882 126919 233938 126928
rect 233896 126313 233924 126919
rect 233882 126304 233938 126313
rect 233882 126239 233938 126248
rect 234712 93220 234764 93226
rect 234712 93162 234764 93168
rect 233252 16546 233464 16574
rect 232504 3664 232556 3670
rect 232504 3606 232556 3612
rect 232228 3120 232280 3126
rect 232228 3062 232280 3068
rect 232240 480 232268 3062
rect 233436 480 233464 16546
rect 234724 6914 234752 93162
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235276 3942 235304 149874
rect 235368 141545 235396 220351
rect 235460 150142 235488 226510
rect 235552 151638 235580 227734
rect 235644 159526 235672 236914
rect 235736 235278 235764 237346
rect 235920 237046 235948 239702
rect 235908 237040 235960 237046
rect 235908 236982 235960 236988
rect 236012 235929 236040 239822
rect 236104 239822 236178 239850
rect 236242 239850 236270 240108
rect 236334 239970 236362 240108
rect 236426 239970 236454 240108
rect 236322 239964 236374 239970
rect 236322 239906 236374 239912
rect 236414 239964 236466 239970
rect 236414 239906 236466 239912
rect 236518 239850 236546 240108
rect 236610 239970 236638 240108
rect 236598 239964 236650 239970
rect 236598 239906 236650 239912
rect 236702 239850 236730 240108
rect 236794 239907 236822 240108
rect 236242 239822 236408 239850
rect 236518 239822 236592 239850
rect 235998 235920 236054 235929
rect 235998 235855 236054 235864
rect 235724 235272 235776 235278
rect 235724 235214 235776 235220
rect 236104 234614 236132 239822
rect 236184 239760 236236 239766
rect 236182 239728 236184 239737
rect 236276 239760 236328 239766
rect 236236 239728 236238 239737
rect 236276 239702 236328 239708
rect 236182 239663 236238 239672
rect 236184 239624 236236 239630
rect 236184 239566 236236 239572
rect 236196 238746 236224 239566
rect 236184 238740 236236 238746
rect 236184 238682 236236 238688
rect 236288 237998 236316 239702
rect 236276 237992 236328 237998
rect 236276 237934 236328 237940
rect 236276 237856 236328 237862
rect 236276 237798 236328 237804
rect 235920 234586 236132 234614
rect 235920 230110 235948 234586
rect 236288 234054 236316 237798
rect 236380 237374 236408 239822
rect 236460 239692 236512 239698
rect 236460 239634 236512 239640
rect 236472 237862 236500 239634
rect 236460 237856 236512 237862
rect 236460 237798 236512 237804
rect 236380 237346 236500 237374
rect 236276 234048 236328 234054
rect 236276 233990 236328 233996
rect 236090 232792 236146 232801
rect 236090 232727 236146 232736
rect 236000 230444 236052 230450
rect 236000 230386 236052 230392
rect 235908 230104 235960 230110
rect 235908 230046 235960 230052
rect 236012 230042 236040 230386
rect 236000 230036 236052 230042
rect 236000 229978 236052 229984
rect 236104 229770 236132 232727
rect 236092 229764 236144 229770
rect 236092 229706 236144 229712
rect 236472 229226 236500 237346
rect 236564 229770 236592 239822
rect 236656 239822 236730 239850
rect 236780 239898 236836 239907
rect 236886 239902 236914 240108
rect 236978 239970 237006 240108
rect 237070 239970 237098 240108
rect 236966 239964 237018 239970
rect 236966 239906 237018 239912
rect 237058 239964 237110 239970
rect 237058 239906 237110 239912
rect 236780 239833 236836 239842
rect 236874 239896 236926 239902
rect 236874 239838 236926 239844
rect 236966 239828 237018 239834
rect 236656 237697 236684 239822
rect 237018 239788 237098 239816
rect 236966 239770 237018 239776
rect 236828 239760 236880 239766
rect 236826 239728 236828 239737
rect 236880 239728 236882 239737
rect 237070 239714 237098 239788
rect 237162 239748 237190 240108
rect 237254 239816 237282 240108
rect 237346 239970 237374 240108
rect 237334 239964 237386 239970
rect 237334 239906 237386 239912
rect 237254 239788 237328 239816
rect 237162 239720 237236 239748
rect 236826 239663 236882 239672
rect 236920 239692 236972 239698
rect 236736 239420 236788 239426
rect 236736 239362 236788 239368
rect 236642 237688 236698 237697
rect 236642 237623 236698 237632
rect 236748 237017 236776 239362
rect 236734 237008 236790 237017
rect 236734 236943 236790 236952
rect 236644 235204 236696 235210
rect 236644 235146 236696 235152
rect 236552 229764 236604 229770
rect 236552 229706 236604 229712
rect 236460 229220 236512 229226
rect 236460 229162 236512 229168
rect 236472 228206 236500 229162
rect 236460 228200 236512 228206
rect 236460 228142 236512 228148
rect 236000 227112 236052 227118
rect 236000 227054 236052 227060
rect 235816 199436 235868 199442
rect 235816 199378 235868 199384
rect 235632 159520 235684 159526
rect 235632 159462 235684 159468
rect 235540 151632 235592 151638
rect 235540 151574 235592 151580
rect 235448 150136 235500 150142
rect 235448 150078 235500 150084
rect 235828 146946 235856 199378
rect 236012 153678 236040 227054
rect 236656 153921 236684 235146
rect 236736 232348 236788 232354
rect 236736 232290 236788 232296
rect 236748 229566 236776 232290
rect 236736 229560 236788 229566
rect 236736 229502 236788 229508
rect 236840 228954 236868 239663
rect 236920 239634 236972 239640
rect 237024 239686 237098 239714
rect 236932 239306 236960 239634
rect 237024 239426 237052 239686
rect 237104 239556 237156 239562
rect 237104 239498 237156 239504
rect 237116 239465 237144 239498
rect 237102 239456 237158 239465
rect 237012 239420 237064 239426
rect 237102 239391 237158 239400
rect 237012 239362 237064 239368
rect 236932 239278 237052 239306
rect 237024 239086 237052 239278
rect 237012 239080 237064 239086
rect 237012 239022 237064 239028
rect 236920 237992 236972 237998
rect 236920 237934 236972 237940
rect 236932 237454 236960 237934
rect 236920 237448 236972 237454
rect 236920 237390 236972 237396
rect 236932 235958 236960 237390
rect 236920 235952 236972 235958
rect 236920 235894 236972 235900
rect 237024 234394 237052 239022
rect 237116 238660 237144 239391
rect 237208 238785 237236 239720
rect 237194 238776 237250 238785
rect 237194 238711 237250 238720
rect 237116 238632 237236 238660
rect 237102 238504 237158 238513
rect 237102 238439 237158 238448
rect 237116 238406 237144 238439
rect 237104 238400 237156 238406
rect 237104 238342 237156 238348
rect 237208 238252 237236 238632
rect 237116 238224 237236 238252
rect 237116 235346 237144 238224
rect 237300 237232 237328 239788
rect 237438 239737 237466 240108
rect 237530 239970 237558 240108
rect 237518 239964 237570 239970
rect 237518 239906 237570 239912
rect 237622 239873 237650 240108
rect 237714 239970 237742 240108
rect 237702 239964 237754 239970
rect 237702 239906 237754 239912
rect 237608 239864 237664 239873
rect 237608 239799 237664 239808
rect 237564 239760 237616 239766
rect 237424 239728 237480 239737
rect 237806 239748 237834 240108
rect 237898 239970 237926 240108
rect 237886 239964 237938 239970
rect 237886 239906 237938 239912
rect 237990 239816 238018 240108
rect 238082 239902 238110 240108
rect 238070 239896 238122 239902
rect 238070 239838 238122 239844
rect 238174 239850 238202 240108
rect 238266 239970 238294 240108
rect 238358 239970 238386 240108
rect 238450 239970 238478 240108
rect 238254 239964 238306 239970
rect 238254 239906 238306 239912
rect 238346 239964 238398 239970
rect 238346 239906 238398 239912
rect 238438 239964 238490 239970
rect 238438 239906 238490 239912
rect 238542 239902 238570 240108
rect 238634 239902 238662 240108
rect 238726 239907 238754 240108
rect 238530 239896 238582 239902
rect 238174 239822 238248 239850
rect 238530 239838 238582 239844
rect 238622 239896 238674 239902
rect 238622 239838 238674 239844
rect 238712 239898 238768 239907
rect 238818 239902 238846 240108
rect 238910 239902 238938 240108
rect 237564 239702 237616 239708
rect 237654 239728 237710 239737
rect 237424 239663 237480 239672
rect 237472 239624 237524 239630
rect 237472 239566 237524 239572
rect 237484 239465 237512 239566
rect 237470 239456 237526 239465
rect 237208 237204 237328 237232
rect 237392 239414 237470 239442
rect 237208 236745 237236 237204
rect 237288 237108 237340 237114
rect 237288 237050 237340 237056
rect 237194 236736 237250 236745
rect 237194 236671 237250 236680
rect 237104 235340 237156 235346
rect 237104 235282 237156 235288
rect 237196 234932 237248 234938
rect 237196 234874 237248 234880
rect 237012 234388 237064 234394
rect 237012 234330 237064 234336
rect 237104 234184 237156 234190
rect 237104 234126 237156 234132
rect 237116 230314 237144 234126
rect 237104 230308 237156 230314
rect 237104 230250 237156 230256
rect 237208 230042 237236 234874
rect 237196 230036 237248 230042
rect 237196 229978 237248 229984
rect 236828 228948 236880 228954
rect 236828 228890 236880 228896
rect 236826 227488 236882 227497
rect 236826 227423 236882 227432
rect 236736 224868 236788 224874
rect 236736 224810 236788 224816
rect 236642 153912 236698 153921
rect 236642 153847 236698 153856
rect 236000 153672 236052 153678
rect 236000 153614 236052 153620
rect 236748 151814 236776 224810
rect 236840 155553 236868 227423
rect 237300 224874 237328 237050
rect 237288 224868 237340 224874
rect 237288 224810 237340 224816
rect 236920 218068 236972 218074
rect 236920 218010 236972 218016
rect 236826 155544 236882 155553
rect 236826 155479 236882 155488
rect 236656 151786 236776 151814
rect 236656 151502 236684 151786
rect 236644 151496 236696 151502
rect 236644 151438 236696 151444
rect 236000 151088 236052 151094
rect 236000 151030 236052 151036
rect 236012 150482 236040 151030
rect 236000 150476 236052 150482
rect 236000 150418 236052 150424
rect 235816 146940 235868 146946
rect 235816 146882 235868 146888
rect 235354 141536 235410 141545
rect 235354 141471 235410 141480
rect 236012 16574 236040 150418
rect 236012 16546 236592 16574
rect 235264 3936 235316 3942
rect 235264 3878 235316 3884
rect 235816 3732 235868 3738
rect 235816 3674 235868 3680
rect 235828 480 235856 3674
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236656 3806 236684 151438
rect 236932 150482 236960 218010
rect 237392 213897 237420 239414
rect 237470 239391 237526 239400
rect 237576 239018 237604 239702
rect 237654 239663 237710 239672
rect 237760 239720 237834 239748
rect 237944 239788 238018 239816
rect 237564 239012 237616 239018
rect 237564 238954 237616 238960
rect 237472 236088 237524 236094
rect 237472 236030 237524 236036
rect 237484 220833 237512 236030
rect 237576 234258 237604 238954
rect 237668 234462 237696 239663
rect 237760 236473 237788 239720
rect 237944 239680 237972 239788
rect 238220 239737 238248 239822
rect 238300 239828 238352 239834
rect 238712 239833 238768 239842
rect 238806 239896 238858 239902
rect 238806 239838 238858 239844
rect 238898 239896 238950 239902
rect 238898 239838 238950 239844
rect 239002 239816 239030 240108
rect 239094 239970 239122 240108
rect 239082 239964 239134 239970
rect 239082 239906 239134 239912
rect 239186 239816 239214 240108
rect 239278 239907 239306 240108
rect 239264 239898 239320 239907
rect 239264 239833 239320 239842
rect 239002 239788 239076 239816
rect 238300 239770 238352 239776
rect 238206 239728 238262 239737
rect 237852 239652 237972 239680
rect 238116 239692 238168 239698
rect 237852 239086 237880 239652
rect 238206 239663 238262 239672
rect 238116 239634 238168 239640
rect 237932 239556 237984 239562
rect 237932 239498 237984 239504
rect 237840 239080 237892 239086
rect 237840 239022 237892 239028
rect 237746 236464 237802 236473
rect 237746 236399 237802 236408
rect 237656 234456 237708 234462
rect 237656 234398 237708 234404
rect 237564 234252 237616 234258
rect 237564 234194 237616 234200
rect 237668 224262 237696 234398
rect 237852 228410 237880 239022
rect 237944 231849 237972 239498
rect 238024 239488 238076 239494
rect 238024 239430 238076 239436
rect 237930 231840 237986 231849
rect 237930 231775 237986 231784
rect 238036 229242 238064 239430
rect 238128 236910 238156 239634
rect 238208 239624 238260 239630
rect 238208 239566 238260 239572
rect 238116 236904 238168 236910
rect 238116 236846 238168 236852
rect 238220 234122 238248 239566
rect 238312 234802 238340 239770
rect 238484 239760 238536 239766
rect 238390 239728 238446 239737
rect 238484 239702 238536 239708
rect 238576 239760 238628 239766
rect 238760 239760 238812 239766
rect 238576 239702 238628 239708
rect 238666 239728 238722 239737
rect 238390 239663 238446 239672
rect 238404 237946 238432 239663
rect 238496 238066 238524 239702
rect 238484 238060 238536 238066
rect 238484 238002 238536 238008
rect 238404 237918 238524 237946
rect 238390 237824 238446 237833
rect 238390 237759 238446 237768
rect 238300 234796 238352 234802
rect 238300 234738 238352 234744
rect 238300 234252 238352 234258
rect 238300 234194 238352 234200
rect 238208 234116 238260 234122
rect 238208 234058 238260 234064
rect 238036 229214 238248 229242
rect 237840 228404 237892 228410
rect 237840 228346 237892 228352
rect 237656 224256 237708 224262
rect 237656 224198 237708 224204
rect 238220 224194 238248 229214
rect 238208 224188 238260 224194
rect 238208 224130 238260 224136
rect 238024 224052 238076 224058
rect 238024 223994 238076 224000
rect 237470 220824 237526 220833
rect 237470 220759 237526 220768
rect 237378 213888 237434 213897
rect 237378 213823 237434 213832
rect 237012 203584 237064 203590
rect 237012 203526 237064 203532
rect 236920 150476 236972 150482
rect 236920 150418 236972 150424
rect 237024 148374 237052 203526
rect 237012 148368 237064 148374
rect 237012 148310 237064 148316
rect 238036 141817 238064 223994
rect 238116 218136 238168 218142
rect 238116 218078 238168 218084
rect 238128 144566 238156 218078
rect 238220 151337 238248 224130
rect 238312 221474 238340 234194
rect 238300 221468 238352 221474
rect 238300 221410 238352 221416
rect 238404 219230 238432 237759
rect 238392 219224 238444 219230
rect 238392 219166 238444 219172
rect 238404 218142 238432 219166
rect 238392 218136 238444 218142
rect 238392 218078 238444 218084
rect 238496 213761 238524 237918
rect 238588 224670 238616 239702
rect 238760 239702 238812 239708
rect 238666 239663 238722 239672
rect 238680 236094 238708 239663
rect 238772 239578 238800 239702
rect 238772 239550 238984 239578
rect 238760 239488 238812 239494
rect 238760 239430 238812 239436
rect 238850 239456 238906 239465
rect 238772 238950 238800 239430
rect 238850 239391 238852 239400
rect 238904 239391 238906 239400
rect 238852 239362 238904 239368
rect 238760 238944 238812 238950
rect 238760 238886 238812 238892
rect 238758 238776 238814 238785
rect 238758 238711 238814 238720
rect 238668 236088 238720 236094
rect 238668 236030 238720 236036
rect 238576 224664 238628 224670
rect 238576 224606 238628 224612
rect 238482 213752 238538 213761
rect 238482 213687 238538 213696
rect 238772 211857 238800 238711
rect 238864 213081 238892 239362
rect 238956 237930 238984 239550
rect 238944 237924 238996 237930
rect 238944 237866 238996 237872
rect 239048 235385 239076 239788
rect 239140 239788 239214 239816
rect 239034 235376 239090 235385
rect 239034 235311 239090 235320
rect 239140 235260 239168 239788
rect 239370 239748 239398 240108
rect 239462 239850 239490 240108
rect 239554 239970 239582 240108
rect 239542 239964 239594 239970
rect 239542 239906 239594 239912
rect 239646 239907 239674 240108
rect 239632 239898 239688 239907
rect 239738 239902 239766 240108
rect 239462 239822 239536 239850
rect 239632 239833 239688 239842
rect 239726 239896 239778 239902
rect 239726 239838 239778 239844
rect 239232 239737 239398 239748
rect 239218 239728 239398 239737
rect 239274 239720 239398 239728
rect 239218 239663 239274 239672
rect 239232 238406 239260 239663
rect 239508 239578 239536 239822
rect 239830 239771 239858 240108
rect 239922 239970 239950 240108
rect 239910 239964 239962 239970
rect 239910 239906 239962 239912
rect 240014 239816 240042 240108
rect 240106 239970 240134 240108
rect 240094 239964 240146 239970
rect 240094 239906 240146 239912
rect 240198 239816 240226 240108
rect 240290 239907 240318 240108
rect 240382 239970 240410 240108
rect 240370 239964 240422 239970
rect 240276 239898 240332 239907
rect 240370 239906 240422 239912
rect 240276 239833 240332 239842
rect 240474 239816 240502 240108
rect 240566 239902 240594 240108
rect 240658 239907 240686 240108
rect 240554 239896 240606 239902
rect 240554 239838 240606 239844
rect 240644 239898 240700 239907
rect 240644 239833 240700 239842
rect 240750 239850 240778 240108
rect 240842 239970 240870 240108
rect 240934 239970 240962 240108
rect 241026 239970 241054 240108
rect 240830 239964 240882 239970
rect 240830 239906 240882 239912
rect 240922 239964 240974 239970
rect 240922 239906 240974 239912
rect 241014 239964 241066 239970
rect 241014 239906 241066 239912
rect 241118 239850 241146 240108
rect 241210 239970 241238 240108
rect 241198 239964 241250 239970
rect 241198 239906 241250 239912
rect 241302 239902 241330 240108
rect 241290 239896 241342 239902
rect 240750 239822 241008 239850
rect 241118 239822 241238 239850
rect 241290 239838 241342 239844
rect 239968 239788 240042 239816
rect 240152 239788 240226 239816
rect 240428 239788 240502 239816
rect 239588 239760 239640 239766
rect 239588 239702 239640 239708
rect 239816 239762 239872 239771
rect 239324 239550 239536 239578
rect 239220 238400 239272 238406
rect 239220 238342 239272 238348
rect 239220 238060 239272 238066
rect 239220 238002 239272 238008
rect 239048 235232 239168 235260
rect 239048 228818 239076 235232
rect 239232 234025 239260 238002
rect 239218 234016 239274 234025
rect 239218 233951 239274 233960
rect 239324 230586 239352 239550
rect 239496 239488 239548 239494
rect 239496 239430 239548 239436
rect 239404 239420 239456 239426
rect 239404 239362 239456 239368
rect 239416 238066 239444 239362
rect 239404 238060 239456 238066
rect 239404 238002 239456 238008
rect 239404 235612 239456 235618
rect 239404 235554 239456 235560
rect 239416 235142 239444 235554
rect 239404 235136 239456 235142
rect 239404 235078 239456 235084
rect 239312 230580 239364 230586
rect 239312 230522 239364 230528
rect 239508 230474 239536 239430
rect 239600 238610 239628 239702
rect 239816 239697 239872 239706
rect 239864 239624 239916 239630
rect 239784 239584 239864 239612
rect 239678 239048 239734 239057
rect 239678 238983 239734 238992
rect 239588 238604 239640 238610
rect 239588 238546 239640 238552
rect 239588 238400 239640 238406
rect 239588 238342 239640 238348
rect 239600 234258 239628 238342
rect 239692 235521 239720 238983
rect 239678 235512 239734 235521
rect 239678 235447 239734 235456
rect 239678 235104 239734 235113
rect 239678 235039 239734 235048
rect 239588 234252 239640 234258
rect 239588 234194 239640 234200
rect 239692 232354 239720 235039
rect 239680 232348 239732 232354
rect 239680 232290 239732 232296
rect 239588 230580 239640 230586
rect 239588 230522 239640 230528
rect 239324 230446 239536 230474
rect 239128 230240 239180 230246
rect 239128 230182 239180 230188
rect 239140 229974 239168 230182
rect 239128 229968 239180 229974
rect 239128 229910 239180 229916
rect 239036 228812 239088 228818
rect 239036 228754 239088 228760
rect 239324 227390 239352 230446
rect 239404 230240 239456 230246
rect 239404 230182 239456 230188
rect 239312 227384 239364 227390
rect 239312 227326 239364 227332
rect 238850 213072 238906 213081
rect 238850 213007 238906 213016
rect 238758 211848 238814 211857
rect 238758 211783 238814 211792
rect 239416 152862 239444 230182
rect 239600 224602 239628 230522
rect 239784 230474 239812 239584
rect 239864 239566 239916 239572
rect 239864 237924 239916 237930
rect 239864 237866 239916 237872
rect 239876 237182 239904 237866
rect 239864 237176 239916 237182
rect 239864 237118 239916 237124
rect 239864 237040 239916 237046
rect 239864 236982 239916 236988
rect 239876 231305 239904 236982
rect 239968 236881 239996 239788
rect 240152 239748 240180 239788
rect 240152 239720 240272 239748
rect 240140 239624 240192 239630
rect 240140 239566 240192 239572
rect 240152 239465 240180 239566
rect 240138 239456 240194 239465
rect 240138 239391 240194 239400
rect 240048 237176 240100 237182
rect 240048 237118 240100 237124
rect 239954 236872 240010 236881
rect 239954 236807 240010 236816
rect 239862 231296 239918 231305
rect 239862 231231 239918 231240
rect 239784 230446 239996 230474
rect 239864 230172 239916 230178
rect 239968 230160 239996 230446
rect 240060 230246 240088 237118
rect 240152 234433 240180 239391
rect 240244 238882 240272 239720
rect 240322 239728 240378 239737
rect 240322 239663 240378 239672
rect 240232 238876 240284 238882
rect 240232 238818 240284 238824
rect 240244 238678 240272 238818
rect 240232 238672 240284 238678
rect 240232 238614 240284 238620
rect 240138 234424 240194 234433
rect 240138 234359 240194 234368
rect 240336 232626 240364 239663
rect 240428 234938 240456 239788
rect 240782 239728 240838 239737
rect 240508 239692 240560 239698
rect 240782 239663 240838 239672
rect 240508 239634 240560 239640
rect 240416 234932 240468 234938
rect 240416 234874 240468 234880
rect 240324 232620 240376 232626
rect 240324 232562 240376 232568
rect 240048 230240 240100 230246
rect 240048 230182 240100 230188
rect 239916 230132 239996 230160
rect 239864 230114 239916 230120
rect 239876 229566 239904 230114
rect 239864 229560 239916 229566
rect 239864 229502 239916 229508
rect 239680 228676 239732 228682
rect 239680 228618 239732 228624
rect 239588 224596 239640 224602
rect 239588 224538 239640 224544
rect 239494 220144 239550 220153
rect 239494 220079 239550 220088
rect 239404 152856 239456 152862
rect 239404 152798 239456 152804
rect 238206 151328 238262 151337
rect 238206 151263 238262 151272
rect 238116 144560 238168 144566
rect 238116 144502 238168 144508
rect 238022 141808 238078 141817
rect 238022 141743 238078 141752
rect 237380 129056 237432 129062
rect 237380 128998 237432 129004
rect 237392 16574 237420 128998
rect 237392 16546 237696 16574
rect 236644 3800 236696 3806
rect 236644 3742 236696 3748
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239416 4010 239444 152798
rect 239508 137329 239536 220079
rect 239600 146810 239628 224538
rect 239692 152561 239720 228618
rect 239772 228404 239824 228410
rect 239772 228346 239824 228352
rect 239784 156777 239812 228346
rect 239864 226908 239916 226914
rect 239864 226850 239916 226856
rect 239876 156942 239904 226850
rect 240520 225690 240548 239634
rect 240692 239624 240744 239630
rect 240692 239566 240744 239572
rect 240600 238944 240652 238950
rect 240600 238886 240652 238892
rect 240612 233986 240640 238886
rect 240704 237046 240732 239566
rect 240796 239494 240824 239663
rect 240876 239556 240928 239562
rect 240876 239498 240928 239504
rect 240784 239488 240836 239494
rect 240784 239430 240836 239436
rect 240692 237040 240744 237046
rect 240692 236982 240744 236988
rect 240784 237040 240836 237046
rect 240784 236982 240836 236988
rect 240692 236904 240744 236910
rect 240692 236846 240744 236852
rect 240600 233980 240652 233986
rect 240600 233922 240652 233928
rect 240508 225684 240560 225690
rect 240508 225626 240560 225632
rect 240704 224330 240732 236846
rect 240796 234190 240824 236982
rect 240888 234938 240916 239498
rect 240980 238746 241008 239822
rect 241210 239714 241238 239822
rect 241394 239816 241422 240108
rect 241486 239970 241514 240108
rect 241474 239964 241526 239970
rect 241474 239906 241526 239912
rect 241578 239873 241606 240108
rect 241564 239864 241620 239873
rect 241394 239788 241468 239816
rect 241564 239799 241620 239808
rect 241060 239692 241112 239698
rect 241060 239634 241112 239640
rect 241164 239686 241238 239714
rect 240968 238740 241020 238746
rect 240968 238682 241020 238688
rect 241072 237046 241100 239634
rect 241164 237114 241192 239686
rect 241244 239624 241296 239630
rect 241244 239566 241296 239572
rect 241152 237108 241204 237114
rect 241152 237050 241204 237056
rect 241060 237040 241112 237046
rect 241060 236982 241112 236988
rect 241256 236858 241284 239566
rect 241336 239488 241388 239494
rect 241334 239456 241336 239465
rect 241388 239456 241390 239465
rect 241334 239391 241390 239400
rect 241440 236910 241468 239788
rect 241670 239748 241698 240108
rect 241624 239720 241698 239748
rect 241520 239692 241572 239698
rect 241520 239634 241572 239640
rect 241532 239057 241560 239634
rect 241518 239048 241574 239057
rect 241518 238983 241574 238992
rect 241624 238048 241652 239720
rect 241762 239680 241790 240108
rect 241854 239902 241882 240108
rect 241946 239970 241974 240108
rect 242038 239970 242066 240108
rect 241934 239964 241986 239970
rect 241934 239906 241986 239912
rect 242026 239964 242078 239970
rect 242026 239906 242078 239912
rect 242130 239907 242158 240108
rect 241842 239896 241894 239902
rect 241842 239838 241894 239844
rect 242116 239898 242172 239907
rect 242116 239833 242172 239842
rect 241888 239760 241940 239766
rect 242072 239760 242124 239766
rect 241888 239702 241940 239708
rect 241978 239728 242034 239737
rect 241532 238020 241652 238048
rect 241716 239652 241790 239680
rect 240980 236830 241284 236858
rect 241428 236904 241480 236910
rect 241428 236846 241480 236852
rect 240876 234932 240928 234938
rect 240876 234874 240928 234880
rect 240874 234832 240930 234841
rect 240874 234767 240930 234776
rect 240784 234184 240836 234190
rect 240784 234126 240836 234132
rect 240888 229838 240916 234767
rect 240980 232762 241008 236830
rect 241532 236722 241560 238020
rect 241610 237960 241666 237969
rect 241610 237895 241612 237904
rect 241664 237895 241666 237904
rect 241612 237866 241664 237872
rect 241256 236694 241560 236722
rect 241150 235920 241206 235929
rect 241150 235855 241206 235864
rect 241060 234932 241112 234938
rect 241060 234874 241112 234880
rect 240968 232756 241020 232762
rect 240968 232698 241020 232704
rect 240968 232620 241020 232626
rect 240968 232562 241020 232568
rect 240980 231742 241008 232562
rect 240968 231736 241020 231742
rect 240968 231678 241020 231684
rect 240980 230382 241008 231678
rect 240968 230376 241020 230382
rect 240968 230318 241020 230324
rect 240876 229832 240928 229838
rect 240876 229774 240928 229780
rect 240888 229702 240916 229774
rect 240876 229696 240928 229702
rect 240876 229638 240928 229644
rect 241072 229094 241100 234874
rect 240980 229066 241100 229094
rect 240876 225004 240928 225010
rect 240876 224946 240928 224952
rect 240692 224324 240744 224330
rect 240692 224266 240744 224272
rect 240784 224256 240836 224262
rect 240784 224198 240836 224204
rect 239954 218104 240010 218113
rect 239954 218039 240010 218048
rect 239968 211993 239996 218039
rect 239954 211984 240010 211993
rect 239954 211919 240010 211928
rect 239864 156936 239916 156942
rect 239864 156878 239916 156884
rect 239770 156768 239826 156777
rect 239770 156703 239826 156712
rect 240796 154358 240824 224198
rect 240784 154352 240836 154358
rect 240784 154294 240836 154300
rect 239678 152552 239734 152561
rect 239678 152487 239734 152496
rect 239588 146804 239640 146810
rect 239588 146746 239640 146752
rect 239494 137320 239550 137329
rect 239494 137255 239550 137264
rect 239404 4004 239456 4010
rect 239404 3946 239456 3952
rect 240508 3800 240560 3806
rect 240508 3742 240560 3748
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 239324 480 239352 3470
rect 240520 480 240548 3742
rect 240796 3534 240824 154294
rect 240888 151230 240916 224946
rect 240980 224534 241008 229066
rect 241164 226166 241192 235855
rect 241152 226160 241204 226166
rect 241152 226102 241204 226108
rect 241164 225010 241192 226102
rect 241152 225004 241204 225010
rect 241152 224946 241204 224952
rect 240968 224528 241020 224534
rect 240968 224470 241020 224476
rect 240980 218074 241008 224470
rect 241256 224262 241284 236694
rect 241336 236632 241388 236638
rect 241336 236574 241388 236580
rect 241348 230314 241376 236574
rect 241716 236065 241744 239652
rect 241796 239488 241848 239494
rect 241796 239430 241848 239436
rect 241702 236056 241758 236065
rect 241702 235991 241758 236000
rect 241808 234546 241836 239430
rect 241900 235929 241928 239702
rect 242222 239748 242250 240108
rect 242072 239702 242124 239708
rect 242176 239720 242250 239748
rect 241978 239663 241980 239672
rect 242032 239663 242034 239672
rect 241980 239634 242032 239640
rect 241978 239456 242034 239465
rect 242084 239442 242112 239702
rect 242034 239414 242112 239442
rect 241978 239391 242034 239400
rect 241886 235920 241942 235929
rect 241886 235855 241942 235864
rect 241886 235784 241942 235793
rect 241886 235719 241942 235728
rect 241440 234518 241836 234546
rect 241440 233646 241468 234518
rect 241428 233640 241480 233646
rect 241428 233582 241480 233588
rect 241336 230308 241388 230314
rect 241336 230250 241388 230256
rect 241244 224256 241296 224262
rect 241244 224198 241296 224204
rect 241256 224126 241284 224198
rect 241244 224120 241296 224126
rect 241244 224062 241296 224068
rect 240968 218068 241020 218074
rect 240968 218010 241020 218016
rect 241348 153882 241376 230250
rect 241336 153876 241388 153882
rect 241336 153818 241388 153824
rect 241440 152930 241468 233582
rect 241704 232620 241756 232626
rect 241704 232562 241756 232568
rect 241716 225554 241744 232562
rect 241704 225548 241756 225554
rect 241704 225490 241756 225496
rect 241900 219434 241928 235719
rect 241992 230081 242020 239391
rect 242072 236088 242124 236094
rect 242072 236030 242124 236036
rect 242084 235958 242112 236030
rect 242072 235952 242124 235958
rect 242072 235894 242124 235900
rect 242176 235890 242204 239720
rect 242314 239680 242342 240108
rect 242406 239970 242434 240108
rect 242394 239964 242446 239970
rect 242394 239906 242446 239912
rect 242498 239816 242526 240108
rect 242268 239652 242342 239680
rect 242452 239788 242526 239816
rect 242164 235884 242216 235890
rect 242164 235826 242216 235832
rect 242072 232212 242124 232218
rect 242072 232154 242124 232160
rect 241978 230072 242034 230081
rect 241978 230007 242034 230016
rect 242084 224262 242112 232154
rect 242164 225004 242216 225010
rect 242164 224946 242216 224952
rect 242072 224256 242124 224262
rect 242072 224198 242124 224204
rect 241808 219406 241928 219434
rect 241428 152924 241480 152930
rect 241428 152866 241480 152872
rect 240876 151224 240928 151230
rect 240876 151166 240928 151172
rect 240888 4078 240916 151166
rect 241808 140554 241836 219406
rect 242176 157146 242204 224946
rect 242268 219065 242296 239652
rect 242452 232218 242480 239788
rect 242590 239748 242618 240108
rect 242682 239816 242710 240108
rect 242774 239970 242802 240108
rect 242866 239970 242894 240108
rect 242958 239970 242986 240108
rect 242762 239964 242814 239970
rect 242762 239906 242814 239912
rect 242854 239964 242906 239970
rect 242854 239906 242906 239912
rect 242946 239964 242998 239970
rect 242946 239906 242998 239912
rect 243050 239902 243078 240108
rect 243142 239970 243170 240108
rect 243130 239964 243182 239970
rect 243130 239906 243182 239912
rect 243038 239896 243090 239902
rect 243038 239838 243090 239844
rect 243234 239816 243262 240108
rect 243326 239970 243354 240108
rect 243418 239970 243446 240108
rect 243314 239964 243366 239970
rect 243314 239906 243366 239912
rect 243406 239964 243458 239970
rect 243406 239906 243458 239912
rect 242682 239788 242940 239816
rect 242590 239720 242664 239748
rect 242532 236700 242584 236706
rect 242532 236642 242584 236648
rect 242440 232212 242492 232218
rect 242440 232154 242492 232160
rect 242544 225486 242572 236642
rect 242636 234569 242664 239720
rect 242806 239728 242862 239737
rect 242716 239692 242768 239698
rect 242806 239663 242808 239672
rect 242716 239634 242768 239640
rect 242860 239663 242862 239672
rect 242808 239634 242860 239640
rect 242622 234560 242678 234569
rect 242622 234495 242678 234504
rect 242728 232626 242756 239634
rect 242912 239034 242940 239788
rect 243188 239788 243262 239816
rect 242992 239692 243044 239698
rect 242992 239634 243044 239640
rect 243084 239692 243136 239698
rect 243084 239634 243136 239640
rect 242820 239006 242940 239034
rect 242820 235822 242848 239006
rect 242900 238060 242952 238066
rect 242900 238002 242952 238008
rect 242808 235816 242860 235822
rect 242808 235758 242860 235764
rect 242716 232620 242768 232626
rect 242716 232562 242768 232568
rect 242912 231854 242940 238002
rect 243004 236638 243032 239634
rect 243096 236706 243124 239634
rect 243084 236700 243136 236706
rect 243084 236642 243136 236648
rect 242992 236632 243044 236638
rect 242992 236574 243044 236580
rect 243188 232422 243216 239788
rect 243510 239748 243538 240108
rect 243602 239816 243630 240108
rect 243694 239970 243722 240108
rect 243682 239964 243734 239970
rect 243682 239906 243734 239912
rect 243786 239850 243814 240108
rect 243878 239970 243906 240108
rect 243866 239964 243918 239970
rect 243866 239906 243918 239912
rect 243740 239822 243814 239850
rect 243602 239788 243676 239816
rect 243510 239720 243584 239748
rect 243268 239692 243320 239698
rect 243268 239634 243320 239640
rect 243280 235657 243308 239634
rect 243452 239624 243504 239630
rect 243452 239566 243504 239572
rect 243360 239556 243412 239562
rect 243360 239498 243412 239504
rect 243266 235648 243322 235657
rect 243266 235583 243322 235592
rect 243372 234598 243400 239498
rect 243464 235346 243492 239566
rect 243452 235340 243504 235346
rect 243452 235282 243504 235288
rect 243450 235104 243506 235113
rect 243450 235039 243506 235048
rect 243360 234592 243412 234598
rect 243360 234534 243412 234540
rect 243176 232416 243228 232422
rect 243176 232358 243228 232364
rect 242820 231826 242940 231854
rect 242624 231804 242676 231810
rect 242624 231746 242676 231752
rect 242532 225480 242584 225486
rect 242532 225422 242584 225428
rect 242544 225010 242572 225422
rect 242532 225004 242584 225010
rect 242532 224946 242584 224952
rect 242636 221542 242664 231746
rect 242716 225548 242768 225554
rect 242716 225490 242768 225496
rect 242624 221536 242676 221542
rect 242624 221478 242676 221484
rect 242254 219056 242310 219065
rect 242254 218991 242310 219000
rect 242268 218793 242296 218991
rect 242254 218784 242310 218793
rect 242254 218719 242310 218728
rect 242728 186998 242756 225490
rect 242716 186992 242768 186998
rect 242716 186934 242768 186940
rect 242164 157140 242216 157146
rect 242164 157082 242216 157088
rect 241796 140548 241848 140554
rect 241796 140490 241848 140496
rect 241520 134564 241572 134570
rect 241520 134506 241572 134512
rect 241532 16574 241560 134506
rect 241532 16546 241744 16574
rect 240876 4072 240928 4078
rect 240876 4014 240928 4020
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 241716 480 241744 16546
rect 242176 3806 242204 157082
rect 242820 151570 242848 231826
rect 243464 226953 243492 235039
rect 243556 234598 243584 239720
rect 243544 234592 243596 234598
rect 243544 234534 243596 234540
rect 243556 233850 243584 234534
rect 243544 233844 243596 233850
rect 243544 233786 243596 233792
rect 243648 231810 243676 239788
rect 243740 237930 243768 239822
rect 243970 239816 243998 240108
rect 244062 239873 244090 240108
rect 244154 239902 244182 240108
rect 244246 239902 244274 240108
rect 244142 239896 244194 239902
rect 243924 239788 243998 239816
rect 244048 239864 244104 239873
rect 244142 239838 244194 239844
rect 244234 239896 244286 239902
rect 244234 239838 244286 239844
rect 244048 239799 244104 239808
rect 244338 239816 244366 240108
rect 244430 239970 244458 240108
rect 244418 239964 244470 239970
rect 244418 239906 244470 239912
rect 244522 239902 244550 240108
rect 244510 239896 244562 239902
rect 244510 239838 244562 239844
rect 244614 239816 244642 240108
rect 244706 239970 244734 240108
rect 244694 239964 244746 239970
rect 244694 239906 244746 239912
rect 244798 239873 244826 240108
rect 244784 239864 244840 239873
rect 244338 239788 244412 239816
rect 244614 239788 244688 239816
rect 244890 239850 244918 240108
rect 244982 239970 245010 240108
rect 244970 239964 245022 239970
rect 244970 239906 245022 239912
rect 245074 239850 245102 240108
rect 244890 239822 244964 239850
rect 244784 239799 244840 239808
rect 243820 239760 243872 239766
rect 243820 239702 243872 239708
rect 243728 237924 243780 237930
rect 243728 237866 243780 237872
rect 243728 235884 243780 235890
rect 243728 235826 243780 235832
rect 243636 231804 243688 231810
rect 243636 231746 243688 231752
rect 243450 226944 243506 226953
rect 243450 226879 243506 226888
rect 243544 225072 243596 225078
rect 243544 225014 243596 225020
rect 242900 224324 242952 224330
rect 242900 224266 242952 224272
rect 242912 171134 242940 224266
rect 242912 171106 243032 171134
rect 242808 151564 242860 151570
rect 242808 151506 242860 151512
rect 242820 151094 242848 151506
rect 243004 151162 243032 171106
rect 243556 154290 243584 225014
rect 243636 225004 243688 225010
rect 243636 224946 243688 224952
rect 243544 154284 243596 154290
rect 243544 154226 243596 154232
rect 242992 151156 243044 151162
rect 242992 151098 243044 151104
rect 242808 151088 242860 151094
rect 242808 151030 242860 151036
rect 243004 16574 243032 151098
rect 243004 16546 243492 16574
rect 242164 3800 242216 3806
rect 242164 3742 242216 3748
rect 242900 3664 242952 3670
rect 242900 3606 242952 3612
rect 242912 480 242940 3606
rect 243464 3482 243492 16546
rect 243556 3670 243584 154226
rect 243648 148714 243676 224946
rect 243740 224398 243768 235826
rect 243832 225418 243860 239702
rect 243924 235521 243952 239788
rect 244096 239760 244148 239766
rect 244002 239728 244058 239737
rect 244096 239702 244148 239708
rect 244002 239663 244004 239672
rect 244056 239663 244058 239672
rect 244004 239634 244056 239640
rect 244004 239556 244056 239562
rect 244004 239498 244056 239504
rect 243910 235512 243966 235521
rect 243910 235447 243966 235456
rect 243912 235340 243964 235346
rect 243912 235282 243964 235288
rect 243924 225758 243952 235282
rect 244016 230382 244044 239498
rect 244108 236774 244136 239702
rect 244188 239692 244240 239698
rect 244188 239634 244240 239640
rect 244096 236768 244148 236774
rect 244096 236710 244148 236716
rect 244200 234297 244228 239634
rect 244384 239562 244412 239788
rect 244556 239692 244608 239698
rect 244556 239634 244608 239640
rect 244464 239624 244516 239630
rect 244464 239566 244516 239572
rect 244372 239556 244424 239562
rect 244372 239498 244424 239504
rect 244370 239456 244426 239465
rect 244370 239391 244372 239400
rect 244424 239391 244426 239400
rect 244372 239362 244424 239368
rect 244384 238785 244412 239362
rect 244370 238776 244426 238785
rect 244370 238711 244426 238720
rect 244476 238649 244504 239566
rect 244462 238640 244518 238649
rect 244462 238575 244518 238584
rect 244186 234288 244242 234297
rect 244186 234223 244242 234232
rect 244188 233844 244240 233850
rect 244188 233786 244240 233792
rect 244096 230444 244148 230450
rect 244096 230386 244148 230392
rect 244004 230376 244056 230382
rect 244004 230318 244056 230324
rect 243912 225752 243964 225758
rect 243912 225694 243964 225700
rect 243820 225412 243872 225418
rect 243820 225354 243872 225360
rect 243832 225078 243860 225354
rect 243820 225072 243872 225078
rect 243820 225014 243872 225020
rect 243924 225010 243952 225694
rect 243912 225004 243964 225010
rect 243912 224946 243964 224952
rect 243728 224392 243780 224398
rect 243728 224334 243780 224340
rect 243740 148850 243768 224334
rect 244016 219434 244044 230318
rect 244108 229158 244136 230386
rect 244096 229152 244148 229158
rect 244096 229094 244148 229100
rect 244108 225622 244136 229094
rect 244096 225616 244148 225622
rect 244096 225558 244148 225564
rect 244016 219406 244136 219434
rect 244002 218240 244058 218249
rect 244002 218175 244058 218184
rect 243818 218104 243874 218113
rect 243818 218039 243874 218048
rect 243832 213353 243860 218039
rect 243818 213344 243874 213353
rect 243818 213279 243874 213288
rect 244016 213246 244044 218175
rect 244004 213240 244056 213246
rect 244004 213182 244056 213188
rect 243728 148844 243780 148850
rect 243728 148786 243780 148792
rect 243636 148708 243688 148714
rect 243636 148650 243688 148656
rect 243648 3738 243676 148650
rect 243740 4146 243768 148786
rect 244108 148782 244136 219406
rect 244096 148776 244148 148782
rect 244096 148718 244148 148724
rect 244108 148374 244136 148718
rect 244096 148368 244148 148374
rect 244096 148310 244148 148316
rect 244200 143206 244228 233786
rect 244476 230217 244504 238575
rect 244568 236910 244596 239634
rect 244556 236904 244608 236910
rect 244556 236846 244608 236852
rect 244556 236428 244608 236434
rect 244556 236370 244608 236376
rect 244568 235686 244596 236370
rect 244556 235680 244608 235686
rect 244556 235622 244608 235628
rect 244660 235006 244688 239788
rect 244740 239760 244792 239766
rect 244936 239714 244964 239822
rect 245028 239822 245102 239850
rect 245028 239766 245056 239822
rect 244740 239702 244792 239708
rect 244752 235550 244780 239702
rect 244844 239686 244964 239714
rect 245016 239760 245068 239766
rect 245166 239748 245194 240108
rect 245258 239816 245286 240108
rect 245350 239970 245378 240108
rect 245338 239964 245390 239970
rect 245338 239906 245390 239912
rect 245442 239816 245470 240108
rect 245534 239970 245562 240108
rect 245626 239970 245654 240108
rect 245522 239964 245574 239970
rect 245522 239906 245574 239912
rect 245614 239964 245666 239970
rect 245614 239906 245666 239912
rect 245718 239902 245746 240108
rect 245706 239896 245758 239902
rect 245706 239838 245758 239844
rect 245258 239788 245332 239816
rect 245442 239788 245608 239816
rect 245016 239702 245068 239708
rect 245120 239720 245194 239748
rect 244844 236638 244872 239686
rect 244924 239624 244976 239630
rect 244924 239566 244976 239572
rect 244832 236632 244884 236638
rect 244832 236574 244884 236580
rect 244832 236496 244884 236502
rect 244832 236438 244884 236444
rect 244740 235544 244792 235550
rect 244740 235486 244792 235492
rect 244648 235000 244700 235006
rect 244648 234942 244700 234948
rect 244844 230450 244872 236438
rect 244936 236162 244964 239566
rect 245016 239420 245068 239426
rect 245016 239362 245068 239368
rect 245028 238066 245056 239362
rect 245016 238060 245068 238066
rect 245016 238002 245068 238008
rect 245120 237776 245148 239720
rect 245200 239624 245252 239630
rect 245200 239566 245252 239572
rect 245212 238746 245240 239566
rect 245304 238898 245332 239788
rect 245580 239714 245608 239788
rect 245810 239748 245838 240108
rect 245902 239907 245930 240108
rect 245994 239970 246022 240108
rect 245982 239964 246034 239970
rect 245888 239898 245944 239907
rect 245982 239906 246034 239912
rect 246086 239902 246114 240108
rect 246178 239902 246206 240108
rect 246270 239902 246298 240108
rect 246362 239902 246390 240108
rect 245888 239833 245944 239842
rect 246074 239896 246126 239902
rect 246074 239838 246126 239844
rect 246166 239896 246218 239902
rect 246166 239838 246218 239844
rect 246258 239896 246310 239902
rect 246258 239838 246310 239844
rect 246350 239896 246402 239902
rect 246350 239838 246402 239844
rect 246454 239816 246482 240108
rect 246546 239970 246574 240108
rect 246638 239970 246666 240108
rect 246534 239964 246586 239970
rect 246534 239906 246586 239912
rect 246626 239964 246678 239970
rect 246626 239906 246678 239912
rect 246578 239864 246634 239873
rect 246454 239808 246578 239816
rect 246730 239850 246758 240108
rect 246822 239970 246850 240108
rect 246810 239964 246862 239970
rect 246810 239906 246862 239912
rect 246914 239850 246942 240108
rect 247006 239970 247034 240108
rect 247098 239970 247126 240108
rect 246994 239964 247046 239970
rect 246994 239906 247046 239912
rect 247086 239964 247138 239970
rect 247086 239906 247138 239912
rect 247190 239873 247218 240108
rect 247282 239970 247310 240108
rect 247374 239970 247402 240108
rect 247270 239964 247322 239970
rect 247270 239906 247322 239912
rect 247362 239964 247414 239970
rect 247362 239906 247414 239912
rect 247176 239864 247232 239873
rect 246730 239822 246804 239850
rect 246914 239822 246988 239850
rect 246454 239799 246634 239808
rect 246454 239788 246620 239799
rect 246028 239760 246080 239766
rect 245810 239720 245884 239748
rect 245580 239686 245700 239714
rect 245476 239624 245528 239630
rect 245476 239566 245528 239572
rect 245568 239624 245620 239630
rect 245568 239566 245620 239572
rect 245304 238870 245424 238898
rect 245292 238808 245344 238814
rect 245396 238785 245424 238870
rect 245292 238750 245344 238756
rect 245382 238776 245438 238785
rect 245200 238740 245252 238746
rect 245200 238682 245252 238688
rect 245028 237748 245148 237776
rect 244924 236156 244976 236162
rect 244924 236098 244976 236104
rect 244924 235816 244976 235822
rect 244924 235758 244976 235764
rect 244936 233782 244964 235758
rect 244924 233776 244976 233782
rect 244924 233718 244976 233724
rect 244832 230444 244884 230450
rect 244832 230386 244884 230392
rect 244462 230208 244518 230217
rect 244462 230143 244518 230152
rect 244740 230172 244792 230178
rect 244740 230114 244792 230120
rect 244280 224256 244332 224262
rect 244280 224198 244332 224204
rect 244292 148510 244320 224198
rect 244280 148504 244332 148510
rect 244280 148446 244332 148452
rect 244292 147694 244320 148446
rect 244280 147688 244332 147694
rect 244280 147630 244332 147636
rect 244188 143200 244240 143206
rect 244188 143142 244240 143148
rect 244752 139262 244780 230114
rect 244936 151706 244964 233718
rect 245028 229430 245056 237748
rect 245106 237688 245162 237697
rect 245106 237623 245162 237632
rect 245016 229424 245068 229430
rect 245016 229366 245068 229372
rect 245028 159118 245056 229366
rect 245120 224738 245148 237623
rect 245212 237017 245240 238682
rect 245198 237008 245254 237017
rect 245198 236943 245254 236952
rect 245304 236892 245332 238750
rect 245382 238711 245438 238720
rect 245382 238640 245438 238649
rect 245382 238575 245438 238584
rect 245212 236864 245332 236892
rect 245212 236706 245240 236864
rect 245200 236700 245252 236706
rect 245200 236642 245252 236648
rect 245212 235754 245240 236642
rect 245292 236632 245344 236638
rect 245292 236574 245344 236580
rect 245200 235748 245252 235754
rect 245200 235690 245252 235696
rect 245200 235000 245252 235006
rect 245200 234942 245252 234948
rect 245212 233102 245240 234942
rect 245200 233096 245252 233102
rect 245200 233038 245252 233044
rect 245212 225894 245240 233038
rect 245304 230450 245332 236574
rect 245292 230444 245344 230450
rect 245292 230386 245344 230392
rect 245304 230178 245332 230386
rect 245292 230172 245344 230178
rect 245292 230114 245344 230120
rect 245292 229696 245344 229702
rect 245292 229638 245344 229644
rect 245200 225888 245252 225894
rect 245200 225830 245252 225836
rect 245108 224732 245160 224738
rect 245108 224674 245160 224680
rect 245304 171154 245332 229638
rect 245292 171148 245344 171154
rect 245120 171106 245292 171134
rect 245016 159112 245068 159118
rect 245016 159054 245068 159060
rect 245028 156670 245056 159054
rect 245016 156664 245068 156670
rect 245016 156606 245068 156612
rect 244924 151700 244976 151706
rect 244924 151642 244976 151648
rect 244936 150482 244964 151642
rect 244924 150476 244976 150482
rect 244924 150418 244976 150424
rect 244924 147688 244976 147694
rect 244924 147630 244976 147636
rect 244740 139256 244792 139262
rect 244740 139198 244792 139204
rect 244278 126304 244334 126313
rect 244278 126239 244334 126248
rect 244292 16574 244320 126239
rect 244292 16546 244872 16574
rect 243728 4140 243780 4146
rect 243728 4082 243780 4088
rect 243636 3732 243688 3738
rect 243636 3674 243688 3680
rect 243544 3664 243596 3670
rect 243544 3606 243596 3612
rect 244844 3482 244872 16546
rect 244936 3874 244964 147630
rect 245120 144430 245148 171106
rect 245292 171090 245344 171096
rect 245396 168434 245424 238575
rect 245488 236502 245516 239566
rect 245580 239193 245608 239566
rect 245566 239184 245622 239193
rect 245566 239119 245622 239128
rect 245476 236496 245528 236502
rect 245476 236438 245528 236444
rect 245476 235408 245528 235414
rect 245476 235350 245528 235356
rect 245488 234734 245516 235350
rect 245476 234728 245528 234734
rect 245476 234670 245528 234676
rect 245488 226030 245516 234670
rect 245580 229702 245608 239119
rect 245672 237114 245700 239686
rect 245856 238814 245884 239720
rect 246028 239702 246080 239708
rect 246120 239760 246172 239766
rect 246672 239760 246724 239766
rect 246578 239728 246634 239737
rect 246172 239708 246252 239714
rect 246120 239702 246252 239708
rect 245934 239184 245990 239193
rect 245934 239119 245990 239128
rect 245844 238808 245896 238814
rect 245844 238750 245896 238756
rect 245660 237108 245712 237114
rect 245660 237050 245712 237056
rect 245660 236156 245712 236162
rect 245660 236098 245712 236104
rect 245672 235006 245700 236098
rect 245948 236042 245976 239119
rect 245764 236014 245976 236042
rect 245660 235000 245712 235006
rect 245660 234942 245712 234948
rect 245764 229702 245792 236014
rect 246040 235940 246068 239702
rect 246132 239686 246252 239702
rect 246118 239592 246174 239601
rect 246118 239527 246174 239536
rect 245856 235912 246068 235940
rect 245568 229696 245620 229702
rect 245568 229638 245620 229644
rect 245752 229696 245804 229702
rect 245752 229638 245804 229644
rect 245476 226024 245528 226030
rect 245476 225966 245528 225972
rect 245476 225888 245528 225894
rect 245476 225830 245528 225836
rect 245384 168428 245436 168434
rect 245384 168370 245436 168376
rect 245396 161474 245424 168370
rect 245212 161446 245424 161474
rect 245212 147354 245240 161446
rect 245200 147348 245252 147354
rect 245200 147290 245252 147296
rect 245488 146198 245516 225830
rect 245856 222902 245884 235912
rect 246132 233850 246160 239527
rect 246224 236178 246252 239686
rect 246304 239692 246356 239698
rect 246304 239634 246356 239640
rect 246488 239692 246540 239698
rect 246672 239702 246724 239708
rect 246578 239663 246634 239672
rect 246488 239634 246540 239640
rect 246316 239426 246344 239634
rect 246304 239420 246356 239426
rect 246304 239362 246356 239368
rect 246394 239184 246450 239193
rect 246394 239119 246450 239128
rect 246408 237998 246436 239119
rect 246500 238882 246528 239634
rect 246592 239562 246620 239663
rect 246580 239556 246632 239562
rect 246580 239498 246632 239504
rect 246488 238876 246540 238882
rect 246488 238818 246540 238824
rect 246684 238754 246712 239702
rect 246500 238726 246712 238754
rect 246396 237992 246448 237998
rect 246396 237934 246448 237940
rect 246224 236150 246436 236178
rect 246304 236020 246356 236026
rect 246304 235962 246356 235968
rect 246120 233844 246172 233850
rect 246120 233786 246172 233792
rect 246316 226098 246344 235962
rect 246408 231854 246436 236150
rect 246500 235414 246528 238726
rect 246580 238060 246632 238066
rect 246580 238002 246632 238008
rect 246592 237046 246620 238002
rect 246580 237040 246632 237046
rect 246580 236982 246632 236988
rect 246488 235408 246540 235414
rect 246488 235350 246540 235356
rect 246776 235226 246804 239822
rect 246856 239760 246908 239766
rect 246856 239702 246908 239708
rect 246684 235198 246804 235226
rect 246684 234530 246712 235198
rect 246672 234524 246724 234530
rect 246672 234466 246724 234472
rect 246408 231826 246620 231854
rect 246394 228712 246450 228721
rect 246394 228647 246450 228656
rect 246304 226092 246356 226098
rect 246304 226034 246356 226040
rect 245844 222896 245896 222902
rect 245844 222838 245896 222844
rect 246304 222896 246356 222902
rect 246304 222838 246356 222844
rect 245660 204264 245712 204270
rect 245660 204206 245712 204212
rect 245672 203590 245700 204206
rect 245660 203584 245712 203590
rect 245660 203526 245712 203532
rect 246316 158166 246344 222838
rect 246304 158160 246356 158166
rect 246304 158102 246356 158108
rect 246304 152924 246356 152930
rect 246304 152866 246356 152872
rect 245476 146192 245528 146198
rect 245476 146134 245528 146140
rect 245108 144424 245160 144430
rect 245108 144366 245160 144372
rect 246316 16574 246344 152866
rect 246408 148578 246436 228647
rect 246592 219298 246620 231826
rect 246764 231668 246816 231674
rect 246764 231610 246816 231616
rect 246672 229696 246724 229702
rect 246672 229638 246724 229644
rect 246684 220590 246712 229638
rect 246672 220584 246724 220590
rect 246672 220526 246724 220532
rect 246580 219292 246632 219298
rect 246580 219234 246632 219240
rect 246592 218142 246620 219234
rect 246580 218136 246632 218142
rect 246580 218078 246632 218084
rect 246488 216572 246540 216578
rect 246488 216514 246540 216520
rect 246500 158234 246528 216514
rect 246776 204270 246804 231610
rect 246868 231402 246896 239702
rect 246960 236026 246988 239822
rect 247466 239816 247494 240108
rect 247558 239902 247586 240108
rect 247546 239896 247598 239902
rect 247546 239838 247598 239844
rect 247176 239799 247232 239808
rect 247328 239788 247494 239816
rect 247132 239760 247184 239766
rect 247132 239702 247184 239708
rect 247224 239760 247276 239766
rect 247224 239702 247276 239708
rect 247040 239692 247092 239698
rect 247040 239634 247092 239640
rect 247052 239601 247080 239634
rect 247038 239592 247094 239601
rect 247038 239527 247094 239536
rect 247040 239420 247092 239426
rect 247040 239362 247092 239368
rect 246948 236020 247000 236026
rect 246948 235962 247000 235968
rect 247052 234530 247080 239362
rect 247144 237998 247172 239702
rect 247132 237992 247184 237998
rect 247132 237934 247184 237940
rect 247236 236638 247264 239702
rect 247328 239601 247356 239788
rect 247500 239624 247552 239630
rect 247314 239592 247370 239601
rect 247650 239612 247678 240108
rect 247742 239907 247770 240108
rect 247728 239898 247784 239907
rect 247728 239833 247784 239842
rect 247834 239748 247862 240108
rect 247500 239566 247552 239572
rect 247604 239584 247678 239612
rect 247788 239720 247862 239748
rect 247926 239748 247954 240108
rect 248018 239970 248046 240108
rect 248006 239964 248058 239970
rect 248006 239906 248058 239912
rect 248110 239816 248138 240108
rect 248064 239788 248138 239816
rect 247926 239720 248000 239748
rect 247314 239527 247370 239536
rect 247316 239488 247368 239494
rect 247316 239430 247368 239436
rect 247328 238814 247356 239430
rect 247408 239420 247460 239426
rect 247408 239362 247460 239368
rect 247420 239193 247448 239362
rect 247406 239184 247462 239193
rect 247406 239119 247462 239128
rect 247316 238808 247368 238814
rect 247316 238750 247368 238756
rect 247406 238776 247462 238785
rect 247406 238711 247462 238720
rect 247420 236960 247448 238711
rect 247512 238649 247540 239566
rect 247498 238640 247554 238649
rect 247498 238575 247554 238584
rect 247328 236932 247448 236960
rect 247224 236632 247276 236638
rect 247224 236574 247276 236580
rect 247222 236056 247278 236065
rect 247132 236020 247184 236026
rect 247222 235991 247278 236000
rect 247132 235962 247184 235968
rect 247040 234524 247092 234530
rect 247040 234466 247092 234472
rect 247052 231854 247080 234466
rect 246960 231826 247080 231854
rect 246856 231396 246908 231402
rect 246856 231338 246908 231344
rect 246856 218136 246908 218142
rect 246856 218078 246908 218084
rect 246764 204264 246816 204270
rect 246764 204206 246816 204212
rect 246868 176730 246896 218078
rect 246580 176724 246632 176730
rect 246580 176666 246632 176672
rect 246856 176724 246908 176730
rect 246856 176666 246908 176672
rect 246488 158228 246540 158234
rect 246488 158170 246540 158176
rect 246396 148572 246448 148578
rect 246396 148514 246448 148520
rect 246592 147286 246620 176666
rect 246580 147280 246632 147286
rect 246580 147222 246632 147228
rect 246960 141846 246988 231826
rect 247040 220720 247092 220726
rect 247040 220662 247092 220668
rect 247052 220114 247080 220662
rect 247040 220108 247092 220114
rect 247040 220050 247092 220056
rect 247144 217326 247172 235962
rect 247236 226137 247264 235991
rect 247328 234666 247356 236932
rect 247406 236872 247462 236881
rect 247406 236807 247462 236816
rect 247316 234660 247368 234666
rect 247316 234602 247368 234608
rect 247222 226128 247278 226137
rect 247222 226063 247278 226072
rect 247236 224058 247264 226063
rect 247224 224052 247276 224058
rect 247224 223994 247276 224000
rect 247132 217320 247184 217326
rect 247132 217262 247184 217268
rect 247040 200116 247092 200122
rect 247040 200058 247092 200064
rect 247052 199442 247080 200058
rect 247040 199436 247092 199442
rect 247040 199378 247092 199384
rect 247328 152794 247356 234602
rect 247420 230178 247448 236807
rect 247604 236586 247632 239584
rect 247684 239488 247736 239494
rect 247684 239430 247736 239436
rect 247696 238134 247724 239430
rect 247684 238128 247736 238134
rect 247684 238070 247736 238076
rect 247512 236558 247632 236586
rect 247684 236632 247736 236638
rect 247684 236574 247736 236580
rect 247512 232490 247540 236558
rect 247500 232484 247552 232490
rect 247500 232426 247552 232432
rect 247408 230172 247460 230178
rect 247408 230114 247460 230120
rect 247420 229974 247448 230114
rect 247408 229968 247460 229974
rect 247408 229910 247460 229916
rect 247512 229498 247540 232426
rect 247592 229968 247644 229974
rect 247592 229910 247644 229916
rect 247604 229838 247632 229910
rect 247592 229832 247644 229838
rect 247592 229774 247644 229780
rect 247500 229492 247552 229498
rect 247500 229434 247552 229440
rect 247696 220726 247724 236574
rect 247788 236065 247816 239720
rect 247868 239624 247920 239630
rect 247868 239566 247920 239572
rect 247774 236056 247830 236065
rect 247774 235991 247830 236000
rect 247880 231854 247908 239566
rect 247972 233578 248000 239720
rect 248064 239601 248092 239788
rect 248202 239748 248230 240108
rect 248156 239720 248230 239748
rect 248050 239592 248106 239601
rect 248050 239527 248106 239536
rect 248052 239284 248104 239290
rect 248052 239226 248104 239232
rect 248064 238921 248092 239226
rect 248050 238912 248106 238921
rect 248050 238847 248106 238856
rect 247960 233572 248012 233578
rect 247960 233514 248012 233520
rect 247880 231826 248000 231854
rect 247774 222864 247830 222873
rect 247774 222799 247830 222808
rect 247684 220720 247736 220726
rect 247684 220662 247736 220668
rect 247684 217320 247736 217326
rect 247684 217262 247736 217268
rect 247316 152788 247368 152794
rect 247316 152730 247368 152736
rect 247696 147150 247724 217262
rect 247788 162353 247816 222799
rect 247972 219434 248000 231826
rect 248156 231062 248184 239720
rect 248294 239680 248322 240108
rect 248386 239850 248414 240108
rect 248478 239970 248506 240108
rect 248466 239964 248518 239970
rect 248466 239906 248518 239912
rect 248570 239873 248598 240108
rect 248662 239970 248690 240108
rect 248754 239970 248782 240108
rect 248846 239970 248874 240108
rect 248938 239970 248966 240108
rect 249030 239970 249058 240108
rect 248650 239964 248702 239970
rect 248650 239906 248702 239912
rect 248742 239964 248794 239970
rect 248742 239906 248794 239912
rect 248834 239964 248886 239970
rect 248834 239906 248886 239912
rect 248926 239964 248978 239970
rect 248926 239906 248978 239912
rect 249018 239964 249070 239970
rect 249018 239906 249070 239912
rect 248556 239864 248612 239873
rect 248386 239822 248460 239850
rect 248248 239652 248322 239680
rect 248248 237374 248276 239652
rect 248328 239488 248380 239494
rect 248328 239430 248380 239436
rect 248340 239154 248368 239430
rect 248328 239148 248380 239154
rect 248328 239090 248380 239096
rect 248432 238649 248460 239822
rect 248556 239799 248612 239808
rect 248970 239864 249026 239873
rect 249122 239850 249150 240108
rect 249214 239970 249242 240108
rect 249202 239964 249254 239970
rect 249202 239906 249254 239912
rect 249306 239902 249334 240108
rect 249398 239970 249426 240108
rect 249490 239970 249518 240108
rect 249386 239964 249438 239970
rect 249386 239906 249438 239912
rect 249478 239964 249530 239970
rect 249478 239906 249530 239912
rect 248970 239799 249026 239808
rect 249076 239822 249150 239850
rect 249294 239896 249346 239902
rect 249582 239850 249610 240108
rect 249674 239902 249702 240108
rect 249766 239907 249794 240108
rect 249294 239838 249346 239844
rect 249536 239822 249610 239850
rect 249662 239896 249714 239902
rect 249662 239838 249714 239844
rect 249752 239898 249808 239907
rect 249858 239902 249886 240108
rect 249950 239970 249978 240108
rect 249938 239964 249990 239970
rect 249938 239906 249990 239912
rect 249752 239833 249808 239842
rect 249846 239896 249898 239902
rect 249846 239838 249898 239844
rect 250042 239850 250070 240108
rect 250134 239970 250162 240108
rect 250122 239964 250174 239970
rect 250122 239906 250174 239912
rect 250226 239850 250254 240108
rect 250318 239970 250346 240108
rect 250306 239964 250358 239970
rect 250306 239906 250358 239912
rect 250410 239850 250438 240108
rect 250502 239970 250530 240108
rect 250594 239970 250622 240108
rect 250490 239964 250542 239970
rect 250490 239906 250542 239912
rect 250582 239964 250634 239970
rect 250582 239906 250634 239912
rect 250042 239822 250116 239850
rect 248512 239760 248564 239766
rect 248512 239702 248564 239708
rect 248696 239760 248748 239766
rect 248696 239702 248748 239708
rect 248788 239760 248840 239766
rect 248788 239702 248840 239708
rect 248524 239329 248552 239702
rect 248602 239592 248658 239601
rect 248602 239527 248658 239536
rect 248510 239320 248566 239329
rect 248510 239255 248566 239264
rect 248512 239148 248564 239154
rect 248512 239090 248564 239096
rect 248524 238950 248552 239090
rect 248512 238944 248564 238950
rect 248512 238886 248564 238892
rect 248418 238640 248474 238649
rect 248418 238575 248474 238584
rect 248510 237960 248566 237969
rect 248510 237895 248566 237904
rect 248248 237346 248460 237374
rect 248236 236632 248288 236638
rect 248236 236574 248288 236580
rect 248144 231056 248196 231062
rect 248144 230998 248196 231004
rect 248248 229786 248276 236574
rect 248432 236026 248460 237346
rect 248420 236020 248472 236026
rect 248420 235962 248472 235968
rect 248328 233368 248380 233374
rect 248328 233310 248380 233316
rect 248156 229758 248276 229786
rect 248050 227352 248106 227361
rect 248050 227287 248106 227296
rect 248064 225593 248092 227287
rect 248050 225584 248106 225593
rect 248050 225519 248106 225528
rect 247880 219406 248000 219434
rect 247880 216578 247908 219406
rect 247868 216572 247920 216578
rect 247868 216514 247920 216520
rect 248156 200122 248184 229758
rect 248340 229650 248368 233310
rect 248248 229622 248368 229650
rect 248144 200116 248196 200122
rect 248144 200058 248196 200064
rect 247774 162344 247830 162353
rect 247774 162279 247830 162288
rect 247684 147144 247736 147150
rect 247684 147086 247736 147092
rect 246948 141840 247000 141846
rect 246948 141782 247000 141788
rect 246960 141642 246988 141782
rect 246948 141636 247000 141642
rect 246948 141578 247000 141584
rect 247316 136468 247368 136474
rect 247316 136410 247368 136416
rect 247328 135998 247356 136410
rect 248248 135998 248276 229622
rect 248328 229492 248380 229498
rect 248328 229434 248380 229440
rect 247316 135992 247368 135998
rect 247316 135934 247368 135940
rect 248236 135992 248288 135998
rect 248236 135934 248288 135940
rect 248340 132394 248368 229434
rect 248524 221882 248552 237895
rect 248616 229362 248644 239527
rect 248708 230081 248736 239702
rect 248800 231674 248828 239702
rect 248880 239692 248932 239698
rect 248984 239680 249012 239799
rect 248932 239652 249012 239680
rect 248880 239634 248932 239640
rect 248880 239556 248932 239562
rect 249076 239544 249104 239822
rect 249156 239760 249208 239766
rect 249156 239702 249208 239708
rect 249248 239760 249300 239766
rect 249248 239702 249300 239708
rect 248880 239498 248932 239504
rect 248984 239516 249104 239544
rect 248892 232966 248920 239498
rect 248984 236638 249012 239516
rect 249064 239420 249116 239426
rect 249064 239362 249116 239368
rect 249076 238678 249104 239362
rect 249168 239193 249196 239702
rect 249154 239184 249210 239193
rect 249154 239119 249210 239128
rect 249260 239034 249288 239702
rect 249340 239692 249392 239698
rect 249340 239634 249392 239640
rect 249168 239006 249288 239034
rect 249064 238672 249116 238678
rect 249064 238614 249116 238620
rect 248972 236632 249024 236638
rect 248972 236574 249024 236580
rect 248880 232960 248932 232966
rect 248880 232902 248932 232908
rect 248788 231668 248840 231674
rect 248788 231610 248840 231616
rect 248694 230072 248750 230081
rect 248892 230058 248920 232902
rect 249168 232626 249196 239006
rect 249248 238944 249300 238950
rect 249248 238886 249300 238892
rect 249260 238746 249288 238886
rect 249248 238740 249300 238746
rect 249248 238682 249300 238688
rect 249156 232620 249208 232626
rect 249156 232562 249208 232568
rect 249248 230512 249300 230518
rect 249248 230454 249300 230460
rect 249064 230444 249116 230450
rect 249064 230386 249116 230392
rect 249076 230246 249104 230386
rect 249064 230240 249116 230246
rect 249064 230182 249116 230188
rect 249260 230178 249288 230454
rect 249248 230172 249300 230178
rect 249248 230114 249300 230120
rect 248892 230030 249104 230058
rect 248694 230007 248750 230016
rect 248604 229356 248656 229362
rect 248604 229298 248656 229304
rect 248972 225004 249024 225010
rect 248972 224946 249024 224952
rect 248512 221876 248564 221882
rect 248512 221818 248564 221824
rect 248984 220794 249012 224946
rect 248972 220788 249024 220794
rect 248972 220730 249024 220736
rect 249076 160818 249104 230030
rect 249248 229832 249300 229838
rect 249248 229774 249300 229780
rect 249260 229566 249288 229774
rect 249248 229560 249300 229566
rect 249248 229502 249300 229508
rect 249248 229356 249300 229362
rect 249248 229298 249300 229304
rect 249156 228812 249208 228818
rect 249156 228754 249208 228760
rect 249064 160812 249116 160818
rect 249064 160754 249116 160760
rect 249168 159633 249196 228754
rect 249260 213246 249288 229298
rect 249352 225010 249380 239634
rect 249432 238672 249484 238678
rect 249432 238614 249484 238620
rect 249444 233170 249472 238614
rect 249432 233164 249484 233170
rect 249432 233106 249484 233112
rect 249340 225004 249392 225010
rect 249340 224946 249392 224952
rect 249444 224954 249472 233106
rect 249536 229362 249564 239822
rect 249616 239760 249668 239766
rect 249616 239702 249668 239708
rect 249628 236434 249656 239702
rect 250088 239680 250116 239822
rect 249996 239652 250116 239680
rect 250180 239822 250254 239850
rect 250364 239822 250438 239850
rect 250534 239864 250590 239873
rect 249708 239624 249760 239630
rect 249706 239592 249708 239601
rect 249800 239624 249852 239630
rect 249760 239592 249762 239601
rect 249800 239566 249852 239572
rect 249706 239527 249762 239536
rect 249706 239320 249762 239329
rect 249706 239255 249762 239264
rect 249616 236428 249668 236434
rect 249616 236370 249668 236376
rect 249720 234705 249748 239255
rect 249706 234696 249762 234705
rect 249706 234631 249762 234640
rect 249812 234326 249840 239566
rect 249892 239556 249944 239562
rect 249892 239498 249944 239504
rect 249800 234320 249852 234326
rect 249800 234262 249852 234268
rect 249812 233374 249840 234262
rect 249800 233368 249852 233374
rect 249800 233310 249852 233316
rect 249524 229356 249576 229362
rect 249524 229298 249576 229304
rect 249904 226302 249932 239498
rect 249996 237425 250024 239652
rect 250076 239556 250128 239562
rect 250076 239498 250128 239504
rect 249982 237416 250038 237425
rect 249982 237351 250038 237360
rect 250088 231606 250116 239498
rect 250180 238610 250208 239822
rect 250260 239760 250312 239766
rect 250260 239702 250312 239708
rect 250272 239465 250300 239702
rect 250258 239456 250314 239465
rect 250258 239391 250314 239400
rect 250168 238604 250220 238610
rect 250168 238546 250220 238552
rect 250076 231600 250128 231606
rect 250076 231542 250128 231548
rect 249892 226296 249944 226302
rect 249892 226238 249944 226244
rect 249444 224926 249748 224954
rect 249430 220824 249486 220833
rect 249340 220788 249392 220794
rect 249430 220759 249486 220768
rect 249340 220730 249392 220736
rect 249352 220114 249380 220730
rect 249340 220108 249392 220114
rect 249340 220050 249392 220056
rect 249248 213240 249300 213246
rect 249248 213182 249300 213188
rect 249154 159624 249210 159633
rect 249154 159559 249210 159568
rect 249260 154426 249288 213182
rect 249352 161158 249380 220050
rect 249444 210361 249472 220759
rect 249430 210352 249486 210361
rect 249430 210287 249486 210296
rect 249340 161152 249392 161158
rect 249340 161094 249392 161100
rect 249248 154420 249300 154426
rect 249248 154362 249300 154368
rect 249064 139256 249116 139262
rect 249064 139198 249116 139204
rect 248328 132388 248380 132394
rect 248328 132330 248380 132336
rect 248340 131850 248368 132330
rect 248328 131844 248380 131850
rect 248328 131786 248380 131792
rect 247682 112432 247738 112441
rect 247682 112367 247738 112376
rect 246316 16546 246620 16574
rect 246592 3942 246620 16546
rect 246396 3936 246448 3942
rect 246396 3878 246448 3884
rect 246580 3936 246632 3942
rect 246580 3878 246632 3884
rect 244924 3868 244976 3874
rect 244924 3810 244976 3816
rect 243464 3454 244136 3482
rect 244844 3454 245240 3482
rect 244108 480 244136 3454
rect 245212 480 245240 3454
rect 246408 480 246436 3878
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 247604 480 247632 3470
rect 247696 3126 247724 112367
rect 249076 3534 249104 139198
rect 249720 135182 249748 224926
rect 250272 221746 250300 239391
rect 250364 235822 250392 239822
rect 250686 239850 250714 240108
rect 250778 239970 250806 240108
rect 250766 239964 250818 239970
rect 250766 239906 250818 239912
rect 250870 239850 250898 240108
rect 250962 239970 250990 240108
rect 250950 239964 251002 239970
rect 250950 239906 251002 239912
rect 250686 239822 250760 239850
rect 250870 239822 250944 239850
rect 250534 239799 250590 239808
rect 250444 239760 250496 239766
rect 250444 239702 250496 239708
rect 250352 235816 250404 235822
rect 250352 235758 250404 235764
rect 250456 225962 250484 239702
rect 250548 239698 250576 239799
rect 250628 239760 250680 239766
rect 250628 239702 250680 239708
rect 250536 239692 250588 239698
rect 250536 239634 250588 239640
rect 250640 239601 250668 239702
rect 250626 239592 250682 239601
rect 250626 239527 250682 239536
rect 250536 239284 250588 239290
rect 250536 239226 250588 239232
rect 250548 238921 250576 239226
rect 250534 238912 250590 238921
rect 250534 238847 250590 238856
rect 250534 238776 250590 238785
rect 250534 238711 250590 238720
rect 250548 234161 250576 238711
rect 250640 234614 250668 239527
rect 250732 236065 250760 239822
rect 250812 239760 250864 239766
rect 250812 239702 250864 239708
rect 250718 236056 250774 236065
rect 250718 235991 250774 236000
rect 250824 235142 250852 239702
rect 250916 239601 250944 239822
rect 251054 239816 251082 240108
rect 251146 239970 251174 240108
rect 251134 239964 251186 239970
rect 251134 239906 251186 239912
rect 251238 239902 251266 240108
rect 251226 239896 251278 239902
rect 251226 239838 251278 239844
rect 251008 239788 251082 239816
rect 250902 239592 250958 239601
rect 250902 239527 250958 239536
rect 250916 238921 250944 239527
rect 250902 238912 250958 238921
rect 250902 238847 250958 238856
rect 250904 238740 250956 238746
rect 250904 238682 250956 238688
rect 250812 235136 250864 235142
rect 250812 235078 250864 235084
rect 250640 234586 250760 234614
rect 250534 234152 250590 234161
rect 250534 234087 250590 234096
rect 250628 226772 250680 226778
rect 250628 226714 250680 226720
rect 250536 226296 250588 226302
rect 250536 226238 250588 226244
rect 250444 225956 250496 225962
rect 250444 225898 250496 225904
rect 250260 221740 250312 221746
rect 250260 221682 250312 221688
rect 250456 158098 250484 225898
rect 250548 225894 250576 226238
rect 250536 225888 250588 225894
rect 250536 225830 250588 225836
rect 250444 158092 250496 158098
rect 250444 158034 250496 158040
rect 250444 150476 250496 150482
rect 250444 150418 250496 150424
rect 249708 135176 249760 135182
rect 249708 135118 249760 135124
rect 249720 134706 249748 135118
rect 249708 134700 249760 134706
rect 249708 134642 249760 134648
rect 250456 4010 250484 150418
rect 250548 147014 250576 225830
rect 250640 161022 250668 226714
rect 250732 184210 250760 234586
rect 250812 231600 250864 231606
rect 250812 231542 250864 231548
rect 250824 226642 250852 231542
rect 250916 230994 250944 238682
rect 251008 231146 251036 239788
rect 251330 239714 251358 240108
rect 251422 239748 251450 240108
rect 251514 239902 251542 240108
rect 251606 239902 251634 240108
rect 251502 239896 251554 239902
rect 251502 239838 251554 239844
rect 251594 239896 251646 239902
rect 251594 239838 251646 239844
rect 251698 239748 251726 240108
rect 251790 239850 251818 240108
rect 251882 239970 251910 240108
rect 251870 239964 251922 239970
rect 251870 239906 251922 239912
rect 251974 239907 252002 240108
rect 251960 239898 252016 239907
rect 251790 239822 251864 239850
rect 251960 239833 252016 239842
rect 251422 239720 251588 239748
rect 251698 239720 251772 239748
rect 251180 239692 251232 239698
rect 251180 239634 251232 239640
rect 251284 239686 251358 239714
rect 251088 239624 251140 239630
rect 251088 239566 251140 239572
rect 251100 232937 251128 239566
rect 251192 238746 251220 239634
rect 251284 238754 251312 239686
rect 251456 239624 251508 239630
rect 251456 239566 251508 239572
rect 251364 239556 251416 239562
rect 251364 239498 251416 239504
rect 251376 239329 251404 239498
rect 251362 239320 251418 239329
rect 251362 239255 251418 239264
rect 251180 238740 251232 238746
rect 251284 238726 251404 238754
rect 251180 238682 251232 238688
rect 251272 238604 251324 238610
rect 251272 238546 251324 238552
rect 251284 234614 251312 238546
rect 251192 234586 251312 234614
rect 251086 232928 251142 232937
rect 251086 232863 251142 232872
rect 251008 231118 251128 231146
rect 250904 230988 250956 230994
rect 250904 230930 250956 230936
rect 250812 226636 250864 226642
rect 250812 226578 250864 226584
rect 250916 224954 250944 230930
rect 251100 227322 251128 231118
rect 251192 228721 251220 234586
rect 251272 229628 251324 229634
rect 251272 229570 251324 229576
rect 251178 228712 251234 228721
rect 251178 228647 251234 228656
rect 251088 227316 251140 227322
rect 251088 227258 251140 227264
rect 251100 226778 251128 227258
rect 251088 226772 251140 226778
rect 251088 226714 251140 226720
rect 251088 226636 251140 226642
rect 251088 226578 251140 226584
rect 250916 224926 251036 224954
rect 250720 184204 250772 184210
rect 250720 184146 250772 184152
rect 250628 161016 250680 161022
rect 250628 160958 250680 160964
rect 250536 147008 250588 147014
rect 250536 146950 250588 146956
rect 251008 146062 251036 224926
rect 251100 146130 251128 226578
rect 251284 222154 251312 229570
rect 251376 223514 251404 238726
rect 251468 238678 251496 239566
rect 251456 238672 251508 238678
rect 251456 238614 251508 238620
rect 251560 237697 251588 239720
rect 251640 239624 251692 239630
rect 251640 239566 251692 239572
rect 251546 237688 251602 237697
rect 251546 237623 251602 237632
rect 251652 229094 251680 239566
rect 251744 230926 251772 239720
rect 251836 239714 251864 239822
rect 252066 239748 252094 240108
rect 252158 239902 252186 240108
rect 252146 239896 252198 239902
rect 252146 239838 252198 239844
rect 252250 239748 252278 240108
rect 252342 239902 252370 240108
rect 252330 239896 252382 239902
rect 252330 239838 252382 239844
rect 252434 239850 252462 240108
rect 252526 239970 252554 240108
rect 252514 239964 252566 239970
rect 252514 239906 252566 239912
rect 252434 239822 252508 239850
rect 252376 239760 252428 239766
rect 252066 239720 252140 239748
rect 252250 239720 252324 239748
rect 251836 239686 251956 239714
rect 251824 239624 251876 239630
rect 251824 239566 251876 239572
rect 251836 238678 251864 239566
rect 251824 238672 251876 238678
rect 251824 238614 251876 238620
rect 251928 234870 251956 239686
rect 252112 239680 252140 239720
rect 252112 239652 252232 239680
rect 252008 239624 252060 239630
rect 252008 239566 252060 239572
rect 252020 238610 252048 239566
rect 252100 239556 252152 239562
rect 252100 239498 252152 239504
rect 252008 238604 252060 238610
rect 252008 238546 252060 238552
rect 251916 234864 251968 234870
rect 251916 234806 251968 234812
rect 252006 234152 252062 234161
rect 252006 234087 252062 234096
rect 252020 232529 252048 234087
rect 252006 232520 252062 232529
rect 252006 232455 252062 232464
rect 251732 230920 251784 230926
rect 251732 230862 251784 230868
rect 251468 229066 251680 229094
rect 251468 223582 251496 229066
rect 252112 224954 252140 239498
rect 252204 239329 252232 239652
rect 252190 239320 252246 239329
rect 252190 239255 252246 239264
rect 252296 239170 252324 239720
rect 252376 239702 252428 239708
rect 252204 239142 252324 239170
rect 252204 234161 252232 239142
rect 252284 237448 252336 237454
rect 252284 237390 252336 237396
rect 252296 236978 252324 237390
rect 252284 236972 252336 236978
rect 252284 236914 252336 236920
rect 252284 235612 252336 235618
rect 252284 235554 252336 235560
rect 252190 234152 252246 234161
rect 252190 234087 252246 234096
rect 252296 232898 252324 235554
rect 252284 232892 252336 232898
rect 252284 232834 252336 232840
rect 252296 231282 252324 232834
rect 252388 231470 252416 239702
rect 252376 231464 252428 231470
rect 252376 231406 252428 231412
rect 252296 231254 252416 231282
rect 252284 230920 252336 230926
rect 252284 230862 252336 230868
rect 252020 224926 252140 224954
rect 252020 224738 252048 224926
rect 252008 224732 252060 224738
rect 252008 224674 252060 224680
rect 251456 223576 251508 223582
rect 251456 223518 251508 223524
rect 251364 223508 251416 223514
rect 251364 223450 251416 223456
rect 251916 223508 251968 223514
rect 251916 223450 251968 223456
rect 251928 223174 251956 223450
rect 251916 223168 251968 223174
rect 251916 223110 251968 223116
rect 251272 222148 251324 222154
rect 251272 222090 251324 222096
rect 251822 221096 251878 221105
rect 251822 221031 251878 221040
rect 251088 146124 251140 146130
rect 251088 146066 251140 146072
rect 250996 146056 251048 146062
rect 250996 145998 251048 146004
rect 251008 145654 251036 145998
rect 251100 145722 251128 146066
rect 251088 145716 251140 145722
rect 251088 145658 251140 145664
rect 250996 145648 251048 145654
rect 250996 145590 251048 145596
rect 251836 145450 251864 221031
rect 251928 147218 251956 223110
rect 252020 148646 252048 224674
rect 252192 223576 252244 223582
rect 252192 223518 252244 223524
rect 252204 223106 252232 223518
rect 252192 223100 252244 223106
rect 252192 223042 252244 223048
rect 252100 222148 252152 222154
rect 252100 222090 252152 222096
rect 252112 221882 252140 222090
rect 252100 221876 252152 221882
rect 252100 221818 252152 221824
rect 252112 150006 252140 221818
rect 252204 153610 252232 223042
rect 252296 220425 252324 230862
rect 252388 224954 252416 231254
rect 252480 229634 252508 239822
rect 252618 239816 252646 240108
rect 252710 239902 252738 240108
rect 252698 239896 252750 239902
rect 252698 239838 252750 239844
rect 252572 239788 252646 239816
rect 252572 236366 252600 239788
rect 252802 239748 252830 240108
rect 252894 239850 252922 240108
rect 252986 239970 253014 240108
rect 252974 239964 253026 239970
rect 252974 239906 253026 239912
rect 253078 239907 253106 240108
rect 253064 239898 253120 239907
rect 253170 239902 253198 240108
rect 252894 239822 252968 239850
rect 253064 239833 253120 239842
rect 253158 239896 253210 239902
rect 253262 239873 253290 240108
rect 253158 239838 253210 239844
rect 253248 239864 253304 239873
rect 252756 239720 252830 239748
rect 252652 239692 252704 239698
rect 252652 239634 252704 239640
rect 252664 237454 252692 239634
rect 252652 237448 252704 237454
rect 252652 237390 252704 237396
rect 252652 237176 252704 237182
rect 252652 237118 252704 237124
rect 252560 236360 252612 236366
rect 252560 236302 252612 236308
rect 252558 233064 252614 233073
rect 252558 232999 252560 233008
rect 252612 232999 252614 233008
rect 252560 232970 252612 232976
rect 252468 229628 252520 229634
rect 252468 229570 252520 229576
rect 252388 224926 252508 224954
rect 252282 220416 252338 220425
rect 252282 220351 252338 220360
rect 252192 153604 252244 153610
rect 252192 153546 252244 153552
rect 252100 150000 252152 150006
rect 252100 149942 252152 149948
rect 252008 148640 252060 148646
rect 252008 148582 252060 148588
rect 251916 147212 251968 147218
rect 251916 147154 251968 147160
rect 251824 145444 251876 145450
rect 251824 145386 251876 145392
rect 252480 133890 252508 224926
rect 252664 222086 252692 237118
rect 252756 233234 252784 239720
rect 252834 239592 252890 239601
rect 252834 239527 252836 239536
rect 252888 239527 252890 239536
rect 252836 239498 252888 239504
rect 252940 235618 252968 239822
rect 253248 239799 253304 239808
rect 253354 239816 253382 240108
rect 253446 239970 253474 240108
rect 253538 239970 253566 240108
rect 253630 239970 253658 240108
rect 253434 239964 253486 239970
rect 253434 239906 253486 239912
rect 253526 239964 253578 239970
rect 253526 239906 253578 239912
rect 253618 239964 253670 239970
rect 253618 239906 253670 239912
rect 253722 239873 253750 240108
rect 253570 239864 253626 239873
rect 253492 239822 253570 239850
rect 253354 239788 253428 239816
rect 253020 239692 253072 239698
rect 253020 239634 253072 239640
rect 253204 239692 253256 239698
rect 253204 239634 253256 239640
rect 253296 239692 253348 239698
rect 253296 239634 253348 239640
rect 253032 236842 253060 239634
rect 253020 236836 253072 236842
rect 253020 236778 253072 236784
rect 252928 235612 252980 235618
rect 252928 235554 252980 235560
rect 252756 233206 252876 233234
rect 252744 229288 252796 229294
rect 252744 229230 252796 229236
rect 252756 222154 252784 229230
rect 252848 224058 252876 233206
rect 253216 233034 253244 239634
rect 253308 237425 253336 239634
rect 253294 237416 253350 237425
rect 253294 237351 253350 237360
rect 253294 237280 253350 237289
rect 253294 237215 253296 237224
rect 253348 237215 253350 237224
rect 253296 237186 253348 237192
rect 253296 237108 253348 237114
rect 253296 237050 253348 237056
rect 253308 236978 253336 237050
rect 253296 236972 253348 236978
rect 253296 236914 253348 236920
rect 253400 233234 253428 239788
rect 253492 236473 253520 239822
rect 253570 239799 253626 239808
rect 253708 239864 253764 239873
rect 253708 239799 253764 239808
rect 253814 239816 253842 240108
rect 253906 239970 253934 240108
rect 253998 239970 254026 240108
rect 253894 239964 253946 239970
rect 253894 239906 253946 239912
rect 253986 239964 254038 239970
rect 253986 239906 254038 239912
rect 254090 239816 254118 240108
rect 253814 239788 253888 239816
rect 253664 239692 253716 239698
rect 253664 239634 253716 239640
rect 253756 239692 253808 239698
rect 253756 239634 253808 239640
rect 253572 239624 253624 239630
rect 253572 239566 253624 239572
rect 253478 236464 253534 236473
rect 253478 236399 253534 236408
rect 253400 233206 253520 233234
rect 253204 233028 253256 233034
rect 253204 232970 253256 232976
rect 252836 224052 252888 224058
rect 252836 223994 252888 224000
rect 252744 222148 252796 222154
rect 252744 222090 252796 222096
rect 252652 222080 252704 222086
rect 252652 222022 252704 222028
rect 253216 160750 253244 232970
rect 253386 231976 253442 231985
rect 253386 231911 253442 231920
rect 253400 224777 253428 231911
rect 253492 224954 253520 233206
rect 253584 232558 253612 239566
rect 253676 237182 253704 239634
rect 253664 237176 253716 237182
rect 253664 237118 253716 237124
rect 253768 236722 253796 239634
rect 253676 236694 253796 236722
rect 253572 232552 253624 232558
rect 253572 232494 253624 232500
rect 253676 231985 253704 236694
rect 253860 233234 253888 239788
rect 254044 239788 254118 239816
rect 253940 239624 253992 239630
rect 253940 239566 253992 239572
rect 253952 237794 253980 239566
rect 253940 237788 253992 237794
rect 253940 237730 253992 237736
rect 253940 236496 253992 236502
rect 253940 236438 253992 236444
rect 253768 233206 253888 233234
rect 253662 231976 253718 231985
rect 253662 231911 253718 231920
rect 253768 229294 253796 233206
rect 253846 230480 253902 230489
rect 253846 230415 253902 230424
rect 253756 229288 253808 229294
rect 253756 229230 253808 229236
rect 253492 224926 253796 224954
rect 253386 224768 253442 224777
rect 253386 224703 253442 224712
rect 253296 224052 253348 224058
rect 253296 223994 253348 224000
rect 253204 160744 253256 160750
rect 253204 160686 253256 160692
rect 253204 153876 253256 153882
rect 253204 153818 253256 153824
rect 252468 133884 252520 133890
rect 252468 133826 252520 133832
rect 252480 133278 252508 133826
rect 252468 133272 252520 133278
rect 252468 133214 252520 133220
rect 251270 98832 251326 98841
rect 251270 98767 251326 98776
rect 251284 16574 251312 98767
rect 253216 16574 253244 153818
rect 253308 137737 253336 223994
rect 253478 222184 253534 222193
rect 253388 222148 253440 222154
rect 253478 222119 253534 222128
rect 253388 222090 253440 222096
rect 253400 221746 253428 222090
rect 253388 221740 253440 221746
rect 253388 221682 253440 221688
rect 253400 145994 253428 221682
rect 253492 152697 253520 222119
rect 253572 222080 253624 222086
rect 253572 222022 253624 222028
rect 253584 158030 253612 222022
rect 253768 219094 253796 224926
rect 253756 219088 253808 219094
rect 253756 219030 253808 219036
rect 253768 165646 253796 219030
rect 253756 165640 253808 165646
rect 253756 165582 253808 165588
rect 253768 161474 253796 165582
rect 253676 161446 253796 161474
rect 253676 158982 253704 161446
rect 253664 158976 253716 158982
rect 253664 158918 253716 158924
rect 253572 158024 253624 158030
rect 253572 157966 253624 157972
rect 253478 152688 253534 152697
rect 253478 152623 253534 152632
rect 253388 145988 253440 145994
rect 253388 145930 253440 145936
rect 253294 137728 253350 137737
rect 253294 137663 253350 137672
rect 253860 129674 253888 230415
rect 253952 218958 253980 236438
rect 254044 235210 254072 239788
rect 254182 239748 254210 240108
rect 254274 239970 254302 240108
rect 254262 239964 254314 239970
rect 254262 239906 254314 239912
rect 254366 239907 254394 240108
rect 254458 239970 254486 240108
rect 254446 239964 254498 239970
rect 254352 239898 254408 239907
rect 254446 239906 254498 239912
rect 254352 239833 254408 239842
rect 254136 239720 254210 239748
rect 254308 239760 254360 239766
rect 254032 235204 254084 235210
rect 254032 235146 254084 235152
rect 254032 221808 254084 221814
rect 254032 221750 254084 221756
rect 254044 221474 254072 221750
rect 254032 221468 254084 221474
rect 254032 221410 254084 221416
rect 254136 220017 254164 239720
rect 254550 239748 254578 240108
rect 254642 239902 254670 240108
rect 254734 239907 254762 240108
rect 254826 239970 254854 240108
rect 254814 239964 254866 239970
rect 254630 239896 254682 239902
rect 254630 239838 254682 239844
rect 254720 239898 254776 239907
rect 254814 239906 254866 239912
rect 254918 239907 254946 240108
rect 255010 239970 255038 240108
rect 255102 239970 255130 240108
rect 254998 239964 255050 239970
rect 254720 239833 254776 239842
rect 254904 239898 254960 239907
rect 254998 239906 255050 239912
rect 255090 239964 255142 239970
rect 255090 239906 255142 239912
rect 255194 239850 255222 240108
rect 255286 239970 255314 240108
rect 255274 239964 255326 239970
rect 255274 239906 255326 239912
rect 254904 239833 254960 239842
rect 255056 239822 255222 239850
rect 254952 239760 255004 239766
rect 254308 239702 254360 239708
rect 254398 239728 254454 239737
rect 254216 239624 254268 239630
rect 254216 239566 254268 239572
rect 254228 221814 254256 239566
rect 254320 237862 254348 239702
rect 254550 239720 254624 239748
rect 254398 239663 254454 239672
rect 254308 237856 254360 237862
rect 254308 237798 254360 237804
rect 254412 237368 254440 239663
rect 254492 239556 254544 239562
rect 254492 239498 254544 239504
rect 254504 237697 254532 239498
rect 254490 237688 254546 237697
rect 254490 237623 254546 237632
rect 254320 237340 254440 237368
rect 254320 222018 254348 237340
rect 254398 237280 254454 237289
rect 254398 237215 254400 237224
rect 254452 237215 254454 237224
rect 254400 237186 254452 237192
rect 254400 237040 254452 237046
rect 254400 236982 254452 236988
rect 254412 222154 254440 236982
rect 254596 236570 254624 239720
rect 254858 239728 254914 239737
rect 254768 239692 254820 239698
rect 254952 239702 255004 239708
rect 254858 239663 254914 239672
rect 254768 239634 254820 239640
rect 254584 236564 254636 236570
rect 254584 236506 254636 236512
rect 254676 235204 254728 235210
rect 254676 235146 254728 235152
rect 254490 231704 254546 231713
rect 254490 231639 254546 231648
rect 254504 230586 254532 231639
rect 254492 230580 254544 230586
rect 254492 230522 254544 230528
rect 254400 222148 254452 222154
rect 254400 222090 254452 222096
rect 254308 222012 254360 222018
rect 254308 221954 254360 221960
rect 254688 221814 254716 235146
rect 254780 231878 254808 239634
rect 254872 237046 254900 239663
rect 254860 237040 254912 237046
rect 254860 236982 254912 236988
rect 254768 231872 254820 231878
rect 254768 231814 254820 231820
rect 254964 229094 254992 239702
rect 255056 236502 255084 239822
rect 255378 239816 255406 240108
rect 255470 239970 255498 240108
rect 255458 239964 255510 239970
rect 255458 239906 255510 239912
rect 255562 239873 255590 240108
rect 255548 239864 255604 239873
rect 255378 239788 255452 239816
rect 255548 239799 255604 239808
rect 255136 239760 255188 239766
rect 255134 239728 255136 239737
rect 255188 239728 255190 239737
rect 255134 239663 255190 239672
rect 255228 239624 255280 239630
rect 255228 239566 255280 239572
rect 255136 239556 255188 239562
rect 255136 239498 255188 239504
rect 255148 236609 255176 239498
rect 255134 236600 255190 236609
rect 255134 236535 255190 236544
rect 255044 236496 255096 236502
rect 255044 236438 255096 236444
rect 255240 233234 255268 239566
rect 255424 239562 255452 239788
rect 255504 239760 255556 239766
rect 255654 239748 255682 240108
rect 255746 239902 255774 240108
rect 255838 239902 255866 240108
rect 255734 239896 255786 239902
rect 255734 239838 255786 239844
rect 255826 239896 255878 239902
rect 255826 239838 255878 239844
rect 255930 239816 255958 240108
rect 256022 239970 256050 240108
rect 256114 239970 256142 240108
rect 256010 239964 256062 239970
rect 256010 239906 256062 239912
rect 256102 239964 256154 239970
rect 256102 239906 256154 239912
rect 256206 239816 256234 240108
rect 256298 239902 256326 240108
rect 256390 239970 256418 240108
rect 256378 239964 256430 239970
rect 256378 239906 256430 239912
rect 256286 239896 256338 239902
rect 256286 239838 256338 239844
rect 256482 239816 256510 240108
rect 256574 239970 256602 240108
rect 256666 239970 256694 240108
rect 256562 239964 256614 239970
rect 256562 239906 256614 239912
rect 256654 239964 256706 239970
rect 256654 239906 256706 239912
rect 256758 239850 256786 240108
rect 255930 239788 256004 239816
rect 255654 239720 255728 239748
rect 255976 239737 256004 239788
rect 256160 239788 256234 239816
rect 256436 239788 256510 239816
rect 256620 239822 256786 239850
rect 255504 239702 255556 239708
rect 255412 239556 255464 239562
rect 255412 239498 255464 239504
rect 255410 239456 255466 239465
rect 255410 239391 255466 239400
rect 255318 239048 255374 239057
rect 255318 238983 255374 238992
rect 255148 233206 255268 233234
rect 255148 229945 255176 233206
rect 255134 229936 255190 229945
rect 255134 229871 255190 229880
rect 254964 229066 255176 229094
rect 254768 222148 254820 222154
rect 254768 222090 254820 222096
rect 254216 221808 254268 221814
rect 254216 221750 254268 221756
rect 254676 221808 254728 221814
rect 254676 221750 254728 221756
rect 254122 220008 254178 220017
rect 254122 219943 254178 219952
rect 254136 219434 254164 219943
rect 254136 219406 254624 219434
rect 253940 218952 253992 218958
rect 253940 218894 253992 218900
rect 254596 137873 254624 219406
rect 254688 145246 254716 221750
rect 254780 145314 254808 222090
rect 254860 222012 254912 222018
rect 254860 221954 254912 221960
rect 254952 222012 255004 222018
rect 254952 221954 255004 221960
rect 254872 145926 254900 221954
rect 254964 221882 254992 221954
rect 254952 221876 255004 221882
rect 254952 221818 255004 221824
rect 255044 221876 255096 221882
rect 255044 221818 255096 221824
rect 255056 221474 255084 221818
rect 255044 221468 255096 221474
rect 255044 221410 255096 221416
rect 255148 219162 255176 229066
rect 255136 219156 255188 219162
rect 255136 219098 255188 219104
rect 254952 218952 255004 218958
rect 254952 218894 255004 218900
rect 254964 218754 254992 218894
rect 254952 218748 255004 218754
rect 254952 218690 255004 218696
rect 254860 145920 254912 145926
rect 254860 145862 254912 145868
rect 254964 145858 254992 218690
rect 255148 214849 255176 219098
rect 255134 214840 255190 214849
rect 255134 214775 255190 214784
rect 255332 214713 255360 238983
rect 255318 214704 255374 214713
rect 255318 214639 255374 214648
rect 255424 147082 255452 239391
rect 255516 234841 255544 239702
rect 255596 239556 255648 239562
rect 255596 239498 255648 239504
rect 255502 234832 255558 234841
rect 255502 234767 255558 234776
rect 255608 225826 255636 239498
rect 255700 237318 255728 239720
rect 255962 239728 256018 239737
rect 255872 239692 255924 239698
rect 256160 239714 256188 239788
rect 255962 239663 256018 239672
rect 256068 239686 256188 239714
rect 256240 239692 256292 239698
rect 255872 239634 255924 239640
rect 255780 239624 255832 239630
rect 255780 239566 255832 239572
rect 255688 237312 255740 237318
rect 255688 237254 255740 237260
rect 255792 236881 255820 239566
rect 255884 239057 255912 239634
rect 255964 239624 256016 239630
rect 255964 239566 256016 239572
rect 255976 239465 256004 239566
rect 255962 239456 256018 239465
rect 255962 239391 256018 239400
rect 255870 239048 255926 239057
rect 255870 238983 255926 238992
rect 255778 236872 255834 236881
rect 255778 236807 255834 236816
rect 255872 236836 255924 236842
rect 255872 236778 255924 236784
rect 255780 236564 255832 236570
rect 255780 236506 255832 236512
rect 255792 226982 255820 236506
rect 255884 234569 255912 236778
rect 256068 236026 256096 239686
rect 256240 239634 256292 239640
rect 256332 239692 256384 239698
rect 256332 239634 256384 239640
rect 256148 239624 256200 239630
rect 256148 239566 256200 239572
rect 256056 236020 256108 236026
rect 256056 235962 256108 235968
rect 256054 234832 256110 234841
rect 256054 234767 256110 234776
rect 255870 234560 255926 234569
rect 255870 234495 255926 234504
rect 256068 232694 256096 234767
rect 256056 232688 256108 232694
rect 256056 232630 256108 232636
rect 256160 231854 256188 239566
rect 255976 231826 256188 231854
rect 255976 229094 256004 231826
rect 256252 229094 256280 239634
rect 256344 237017 256372 239634
rect 256330 237008 256386 237017
rect 256330 236943 256386 236952
rect 256436 236570 256464 239788
rect 256516 239556 256568 239562
rect 256516 239498 256568 239504
rect 256424 236564 256476 236570
rect 256424 236506 256476 236512
rect 256528 236450 256556 239498
rect 256436 236422 256556 236450
rect 256436 235482 256464 236422
rect 256514 236328 256570 236337
rect 256514 236263 256570 236272
rect 256424 235476 256476 235482
rect 256424 235418 256476 235424
rect 256436 234433 256464 235418
rect 256422 234424 256478 234433
rect 256422 234359 256478 234368
rect 255976 229066 256188 229094
rect 256252 229066 256464 229094
rect 255780 226976 255832 226982
rect 255780 226918 255832 226924
rect 255596 225820 255648 225826
rect 255596 225762 255648 225768
rect 255964 225820 256016 225826
rect 255964 225762 256016 225768
rect 255412 147076 255464 147082
rect 255412 147018 255464 147024
rect 254952 145852 255004 145858
rect 254952 145794 255004 145800
rect 255976 145790 256004 225762
rect 256056 223372 256108 223378
rect 256056 223314 256108 223320
rect 256068 148442 256096 223314
rect 256160 219434 256188 229066
rect 256436 223378 256464 229066
rect 256424 223372 256476 223378
rect 256424 223314 256476 223320
rect 256528 220289 256556 236263
rect 256620 227186 256648 239822
rect 256850 239748 256878 240108
rect 256942 239970 256970 240108
rect 256930 239964 256982 239970
rect 256930 239906 256982 239912
rect 257034 239816 257062 240108
rect 257126 239970 257154 240108
rect 257114 239964 257166 239970
rect 257114 239906 257166 239912
rect 257218 239902 257246 240108
rect 257310 239970 257338 240108
rect 257298 239964 257350 239970
rect 257298 239906 257350 239912
rect 257206 239896 257258 239902
rect 256804 239720 256878 239748
rect 256988 239788 257062 239816
rect 257204 239864 257206 239873
rect 257258 239864 257260 239873
rect 257402 239850 257430 240108
rect 257494 239970 257522 240108
rect 257586 239970 257614 240108
rect 257482 239964 257534 239970
rect 257482 239906 257534 239912
rect 257574 239964 257626 239970
rect 257574 239906 257626 239912
rect 257204 239799 257260 239808
rect 257356 239822 257430 239850
rect 256700 233640 256752 233646
rect 256700 233582 256752 233588
rect 256608 227180 256660 227186
rect 256608 227122 256660 227128
rect 256514 220280 256570 220289
rect 256514 220215 256570 220224
rect 256160 219406 256464 219434
rect 256436 219366 256464 219406
rect 256424 219360 256476 219366
rect 256424 219302 256476 219308
rect 256436 180794 256464 219302
rect 256160 180766 256464 180794
rect 256160 173942 256188 180766
rect 256528 174010 256556 220215
rect 256240 174004 256292 174010
rect 256240 173946 256292 173952
rect 256516 174004 256568 174010
rect 256516 173946 256568 173952
rect 256148 173936 256200 173942
rect 256148 173878 256200 173884
rect 256160 150249 256188 173878
rect 256252 163577 256280 173946
rect 256238 163568 256294 163577
rect 256238 163503 256294 163512
rect 256146 150240 256202 150249
rect 256146 150175 256202 150184
rect 256056 148436 256108 148442
rect 256056 148378 256108 148384
rect 255964 145784 256016 145790
rect 255964 145726 256016 145732
rect 254768 145308 254820 145314
rect 254768 145250 254820 145256
rect 254676 145240 254728 145246
rect 254676 145182 254728 145188
rect 254582 137864 254638 137873
rect 254582 137799 254638 137808
rect 255872 136536 255924 136542
rect 255872 136478 255924 136484
rect 255884 135930 255912 136478
rect 256620 135930 256648 227122
rect 256712 223446 256740 233582
rect 256804 231674 256832 239720
rect 256884 239624 256936 239630
rect 256884 239566 256936 239572
rect 256896 239465 256924 239566
rect 256882 239456 256938 239465
rect 256882 239391 256938 239400
rect 256896 238649 256924 239391
rect 256882 238640 256938 238649
rect 256882 238575 256938 238584
rect 256988 236094 257016 239788
rect 257160 239760 257212 239766
rect 257066 239728 257122 239737
rect 257160 239702 257212 239708
rect 257250 239728 257306 239737
rect 257066 239663 257122 239672
rect 257080 239562 257108 239663
rect 257068 239556 257120 239562
rect 257068 239498 257120 239504
rect 257172 238746 257200 239702
rect 257250 239663 257306 239672
rect 257160 238740 257212 238746
rect 257160 238682 257212 238688
rect 256976 236088 257028 236094
rect 256976 236030 257028 236036
rect 257264 235074 257292 239663
rect 256884 235068 256936 235074
rect 256884 235010 256936 235016
rect 257252 235068 257304 235074
rect 257252 235010 257304 235016
rect 256792 231668 256844 231674
rect 256792 231610 256844 231616
rect 256804 230926 256832 231610
rect 256792 230920 256844 230926
rect 256792 230862 256844 230868
rect 256896 223514 256924 235010
rect 257356 234614 257384 239822
rect 257678 239816 257706 240108
rect 257770 239970 257798 240108
rect 257862 239970 257890 240108
rect 257758 239964 257810 239970
rect 257758 239906 257810 239912
rect 257850 239964 257902 239970
rect 257850 239906 257902 239912
rect 257954 239850 257982 240108
rect 257494 239788 257706 239816
rect 257816 239822 257982 239850
rect 257494 239748 257522 239788
rect 256988 234586 257384 234614
rect 257448 239720 257522 239748
rect 257816 239737 257844 239822
rect 258046 239748 258074 240108
rect 258138 239907 258166 240108
rect 258124 239898 258180 239907
rect 258230 239902 258258 240108
rect 258124 239833 258180 239842
rect 258218 239896 258270 239902
rect 258322 239873 258350 240108
rect 258414 239970 258442 240108
rect 258506 239970 258534 240108
rect 258402 239964 258454 239970
rect 258402 239906 258454 239912
rect 258494 239964 258546 239970
rect 258494 239906 258546 239912
rect 258598 239873 258626 240108
rect 258690 239970 258718 240108
rect 258678 239964 258730 239970
rect 258678 239906 258730 239912
rect 258782 239873 258810 240108
rect 258874 239970 258902 240108
rect 258862 239964 258914 239970
rect 258862 239906 258914 239912
rect 258218 239838 258270 239844
rect 258308 239864 258364 239873
rect 258584 239864 258640 239873
rect 258308 239799 258364 239808
rect 258448 239828 258500 239834
rect 258768 239864 258824 239873
rect 258640 239808 258672 239816
rect 258584 239799 258672 239808
rect 258966 239816 258994 240108
rect 258768 239799 258824 239808
rect 258598 239788 258672 239799
rect 258448 239770 258500 239776
rect 258356 239760 258408 239766
rect 257802 239728 257858 239737
rect 256988 224233 257016 234586
rect 257448 233646 257476 239720
rect 257620 239692 257672 239698
rect 257620 239634 257672 239640
rect 257712 239692 257764 239698
rect 258046 239720 258212 239748
rect 257802 239663 257858 239672
rect 257712 239634 257764 239640
rect 257528 239624 257580 239630
rect 257528 239566 257580 239572
rect 257436 233640 257488 233646
rect 257436 233582 257488 233588
rect 257068 230920 257120 230926
rect 257068 230862 257120 230868
rect 257080 227254 257108 230862
rect 257540 229094 257568 239566
rect 257632 235210 257660 239634
rect 257620 235204 257672 235210
rect 257620 235146 257672 235152
rect 257724 233481 257752 239634
rect 257804 239556 257856 239562
rect 257804 239498 257856 239504
rect 257988 239556 258040 239562
rect 257988 239498 258040 239504
rect 257710 233472 257766 233481
rect 257710 233407 257766 233416
rect 257540 229066 257660 229094
rect 257068 227248 257120 227254
rect 257068 227190 257120 227196
rect 256974 224224 257030 224233
rect 256974 224159 257030 224168
rect 256884 223508 256936 223514
rect 256884 223450 256936 223456
rect 257344 223508 257396 223514
rect 257344 223450 257396 223456
rect 256700 223440 256752 223446
rect 256700 223382 256752 223388
rect 257356 145586 257384 223450
rect 257436 223440 257488 223446
rect 257436 223382 257488 223388
rect 257448 150074 257476 223382
rect 257526 221776 257582 221785
rect 257526 221711 257582 221720
rect 257540 210497 257568 221711
rect 257632 220182 257660 229066
rect 257620 220176 257672 220182
rect 257620 220118 257672 220124
rect 257526 210488 257582 210497
rect 257526 210423 257582 210432
rect 257816 186386 257844 239498
rect 257896 238740 257948 238746
rect 257896 238682 257948 238688
rect 257908 229094 257936 238682
rect 258000 237726 258028 239498
rect 258078 238776 258134 238785
rect 258078 238711 258134 238720
rect 257988 237720 258040 237726
rect 257988 237662 258040 237668
rect 257908 229066 258028 229094
rect 257528 186380 257580 186386
rect 257528 186322 257580 186328
rect 257804 186380 257856 186386
rect 257804 186322 257856 186328
rect 257436 150068 257488 150074
rect 257436 150010 257488 150016
rect 257344 145580 257396 145586
rect 257344 145522 257396 145528
rect 257540 144498 257568 186322
rect 258000 167074 258028 229066
rect 258092 215529 258120 238711
rect 258184 231713 258212 239720
rect 258356 239702 258408 239708
rect 258264 239624 258316 239630
rect 258264 239566 258316 239572
rect 258276 233889 258304 239566
rect 258368 235278 258396 239702
rect 258356 235272 258408 235278
rect 258356 235214 258408 235220
rect 258356 234728 258408 234734
rect 258356 234670 258408 234676
rect 258262 233880 258318 233889
rect 258262 233815 258318 233824
rect 258264 233300 258316 233306
rect 258264 233242 258316 233248
rect 258170 231704 258226 231713
rect 258170 231639 258226 231648
rect 258276 230722 258304 233242
rect 258264 230716 258316 230722
rect 258264 230658 258316 230664
rect 258276 226302 258304 230658
rect 258368 227254 258396 234670
rect 258460 229090 258488 239770
rect 258540 239692 258592 239698
rect 258540 239634 258592 239640
rect 258552 239465 258580 239634
rect 258538 239456 258594 239465
rect 258538 239391 258594 239400
rect 258644 239306 258672 239788
rect 258920 239788 258994 239816
rect 259058 239816 259086 240108
rect 259150 239970 259178 240108
rect 259138 239964 259190 239970
rect 259138 239906 259190 239912
rect 259242 239850 259270 240108
rect 259334 239970 259362 240108
rect 259322 239964 259374 239970
rect 259322 239906 259374 239912
rect 259242 239822 259316 239850
rect 259058 239788 259132 239816
rect 258816 239760 258868 239766
rect 258816 239702 258868 239708
rect 258722 239456 258778 239465
rect 258722 239391 258778 239400
rect 258552 239278 258672 239306
rect 258552 231130 258580 239278
rect 258630 238640 258686 238649
rect 258630 238575 258686 238584
rect 258644 238377 258672 238575
rect 258630 238368 258686 238377
rect 258630 238303 258686 238312
rect 258630 238232 258686 238241
rect 258630 238167 258686 238176
rect 258644 237697 258672 238167
rect 258630 237688 258686 237697
rect 258630 237623 258686 237632
rect 258630 237416 258686 237425
rect 258630 237351 258686 237360
rect 258540 231124 258592 231130
rect 258540 231066 258592 231072
rect 258448 229084 258500 229090
rect 258448 229026 258500 229032
rect 258460 228818 258488 229026
rect 258448 228812 258500 228818
rect 258448 228754 258500 228760
rect 258356 227248 258408 227254
rect 258356 227190 258408 227196
rect 258264 226296 258316 226302
rect 258264 226238 258316 226244
rect 258078 215520 258134 215529
rect 258078 215455 258134 215464
rect 257620 167068 257672 167074
rect 257620 167010 257672 167016
rect 257988 167068 258040 167074
rect 257988 167010 258040 167016
rect 257632 151473 257660 167010
rect 258644 152998 258672 237351
rect 258736 229094 258764 239391
rect 258828 238785 258856 239702
rect 258814 238776 258870 238785
rect 258814 238711 258870 238720
rect 258816 238672 258868 238678
rect 258816 238614 258868 238620
rect 258828 231130 258856 238614
rect 258920 238241 258948 239788
rect 259104 239714 259132 239788
rect 259012 239686 259132 239714
rect 259184 239760 259236 239766
rect 259184 239702 259236 239708
rect 258906 238232 258962 238241
rect 258906 238167 258962 238176
rect 258908 237924 258960 237930
rect 258908 237866 258960 237872
rect 258920 236978 258948 237866
rect 258908 236972 258960 236978
rect 258908 236914 258960 236920
rect 258816 231124 258868 231130
rect 258816 231066 258868 231072
rect 258736 229066 258948 229094
rect 258722 225992 258778 226001
rect 258722 225927 258778 225936
rect 258736 220794 258764 225927
rect 258920 223242 258948 229066
rect 259012 223582 259040 239686
rect 259092 239624 259144 239630
rect 259092 239566 259144 239572
rect 259104 231334 259132 239566
rect 259196 236570 259224 239702
rect 259184 236564 259236 236570
rect 259184 236506 259236 236512
rect 259288 234734 259316 239822
rect 259426 239816 259454 240108
rect 259518 239907 259546 240108
rect 259504 239898 259560 239907
rect 259504 239833 259560 239842
rect 259380 239788 259454 239816
rect 259610 239816 259638 240108
rect 259702 239970 259730 240108
rect 259690 239964 259742 239970
rect 259690 239906 259742 239912
rect 259794 239816 259822 240108
rect 259610 239788 259684 239816
rect 259276 234728 259328 234734
rect 259276 234670 259328 234676
rect 259380 233306 259408 239788
rect 259656 239737 259684 239788
rect 259748 239788 259822 239816
rect 259642 239728 259698 239737
rect 259460 239692 259512 239698
rect 259460 239634 259512 239640
rect 259564 239686 259642 239714
rect 259472 236337 259500 239634
rect 259564 237046 259592 239686
rect 259642 239663 259698 239672
rect 259644 239624 259696 239630
rect 259644 239566 259696 239572
rect 259552 237040 259604 237046
rect 259552 236982 259604 236988
rect 259458 236328 259514 236337
rect 259458 236263 259514 236272
rect 259550 235376 259606 235385
rect 259550 235311 259606 235320
rect 259460 235272 259512 235278
rect 259460 235214 259512 235220
rect 259472 235074 259500 235214
rect 259460 235068 259512 235074
rect 259460 235010 259512 235016
rect 259564 234977 259592 235311
rect 259550 234968 259606 234977
rect 259550 234903 259606 234912
rect 259368 233300 259420 233306
rect 259368 233242 259420 233248
rect 259092 231328 259144 231334
rect 259092 231270 259144 231276
rect 259656 231198 259684 239566
rect 259748 237930 259776 239788
rect 259886 239748 259914 240108
rect 259978 239850 260006 240108
rect 260070 239970 260098 240108
rect 260058 239964 260110 239970
rect 260058 239906 260110 239912
rect 260162 239850 260190 240108
rect 259978 239822 260052 239850
rect 259840 239720 259914 239748
rect 259840 238202 259868 239720
rect 259920 239624 259972 239630
rect 259920 239566 259972 239572
rect 259932 239465 259960 239566
rect 259918 239456 259974 239465
rect 259918 239391 259974 239400
rect 259828 238196 259880 238202
rect 259828 238138 259880 238144
rect 259736 237924 259788 237930
rect 259736 237866 259788 237872
rect 259734 237824 259790 237833
rect 259734 237759 259790 237768
rect 259748 235385 259776 237759
rect 259920 237720 259972 237726
rect 259920 237662 259972 237668
rect 259734 235376 259790 235385
rect 259734 235311 259790 235320
rect 259644 231192 259696 231198
rect 259644 231134 259696 231140
rect 259932 228750 259960 237662
rect 260024 233646 260052 239822
rect 260116 239822 260190 239850
rect 260012 233640 260064 233646
rect 260012 233582 260064 233588
rect 260116 229022 260144 239822
rect 260254 239748 260282 240108
rect 260346 239850 260374 240108
rect 260438 239970 260466 240108
rect 260530 239970 260558 240108
rect 260622 239970 260650 240108
rect 260714 239970 260742 240108
rect 260426 239964 260478 239970
rect 260426 239906 260478 239912
rect 260518 239964 260570 239970
rect 260518 239906 260570 239912
rect 260610 239964 260662 239970
rect 260610 239906 260662 239912
rect 260702 239964 260754 239970
rect 260702 239906 260754 239912
rect 260806 239873 260834 240108
rect 260792 239864 260848 239873
rect 260346 239822 260420 239850
rect 260254 239720 260328 239748
rect 260196 239624 260248 239630
rect 260196 239566 260248 239572
rect 260208 235618 260236 239566
rect 260300 237833 260328 239720
rect 260286 237824 260342 237833
rect 260286 237759 260342 237768
rect 260392 237425 260420 239822
rect 260472 239828 260524 239834
rect 260472 239770 260524 239776
rect 260564 239828 260616 239834
rect 260792 239799 260848 239808
rect 260898 239816 260926 240108
rect 260990 239970 261018 240108
rect 260978 239964 261030 239970
rect 260978 239906 261030 239912
rect 261082 239816 261110 240108
rect 261174 239907 261202 240108
rect 261160 239898 261216 239907
rect 261266 239902 261294 240108
rect 261358 239902 261386 240108
rect 261450 239970 261478 240108
rect 261438 239964 261490 239970
rect 261438 239906 261490 239912
rect 261160 239833 261216 239842
rect 261254 239896 261306 239902
rect 261254 239838 261306 239844
rect 261346 239896 261398 239902
rect 261542 239873 261570 240108
rect 261634 239902 261662 240108
rect 261726 239902 261754 240108
rect 261622 239896 261674 239902
rect 261346 239838 261398 239844
rect 261528 239864 261584 239873
rect 260898 239788 260972 239816
rect 260564 239770 260616 239776
rect 260484 238746 260512 239770
rect 260472 238740 260524 238746
rect 260472 238682 260524 238688
rect 260472 237856 260524 237862
rect 260472 237798 260524 237804
rect 260378 237416 260434 237425
rect 260378 237351 260434 237360
rect 260484 237046 260512 237798
rect 260288 237040 260340 237046
rect 260288 236982 260340 236988
rect 260472 237040 260524 237046
rect 260472 236982 260524 236988
rect 260196 235612 260248 235618
rect 260196 235554 260248 235560
rect 260196 232416 260248 232422
rect 260196 232358 260248 232364
rect 260104 229016 260156 229022
rect 260104 228958 260156 228964
rect 259920 228744 259972 228750
rect 259920 228686 259972 228692
rect 260116 228410 260144 228958
rect 260104 228404 260156 228410
rect 260104 228346 260156 228352
rect 259090 226400 259146 226409
rect 259090 226335 259146 226344
rect 260104 226364 260156 226370
rect 259000 223576 259052 223582
rect 259000 223518 259052 223524
rect 258908 223236 258960 223242
rect 258908 223178 258960 223184
rect 258724 220788 258776 220794
rect 258724 220730 258776 220736
rect 258632 152992 258684 152998
rect 258632 152934 258684 152940
rect 257618 151464 257674 151473
rect 257618 151399 257674 151408
rect 257528 144492 257580 144498
rect 257528 144434 257580 144440
rect 258736 139233 258764 220730
rect 258814 215384 258870 215393
rect 258814 215319 258870 215328
rect 258828 140622 258856 215319
rect 258920 160993 258948 223178
rect 259012 162217 259040 223518
rect 259104 202162 259132 226335
rect 260104 226306 260156 226312
rect 259366 216608 259422 216617
rect 259366 216543 259422 216552
rect 259380 215529 259408 216543
rect 259366 215520 259422 215529
rect 259366 215455 259422 215464
rect 259092 202156 259144 202162
rect 259092 202098 259144 202104
rect 259380 175302 259408 215455
rect 259460 186992 259512 186998
rect 259460 186934 259512 186940
rect 259368 175296 259420 175302
rect 259368 175238 259420 175244
rect 258998 162208 259054 162217
rect 258998 162143 259054 162152
rect 259380 161474 259408 175238
rect 259104 161446 259408 161474
rect 259104 161129 259132 161446
rect 259090 161120 259146 161129
rect 259090 161055 259146 161064
rect 258906 160984 258962 160993
rect 258906 160919 258962 160928
rect 259472 150210 259500 186934
rect 260116 159361 260144 226306
rect 260102 159352 260158 159361
rect 260102 159287 260158 159296
rect 259460 150204 259512 150210
rect 259460 150146 259512 150152
rect 259472 149122 259500 150146
rect 259460 149116 259512 149122
rect 259460 149058 259512 149064
rect 260104 149116 260156 149122
rect 260104 149058 260156 149064
rect 258816 140616 258868 140622
rect 258816 140558 258868 140564
rect 258722 139224 258778 139233
rect 258722 139159 258778 139168
rect 255872 135924 255924 135930
rect 255872 135866 255924 135872
rect 256608 135924 256660 135930
rect 256608 135866 256660 135872
rect 253848 129668 253900 129674
rect 253848 129610 253900 129616
rect 253860 129130 253888 129610
rect 253848 129124 253900 129130
rect 253848 129066 253900 129072
rect 255318 127664 255374 127673
rect 255318 127599 255374 127608
rect 255332 16574 255360 127599
rect 258722 124808 258778 124817
rect 258722 124743 258778 124752
rect 251284 16546 252416 16574
rect 253216 16546 253612 16574
rect 255332 16546 255912 16574
rect 251180 4072 251232 4078
rect 251180 4014 251232 4020
rect 249984 4004 250036 4010
rect 249984 3946 250036 3952
rect 250444 4004 250496 4010
rect 250444 3946 250496 3952
rect 249064 3528 249116 3534
rect 249064 3470 249116 3476
rect 247684 3120 247736 3126
rect 247684 3062 247736 3068
rect 248788 3120 248840 3126
rect 248788 3062 248840 3068
rect 248800 480 248828 3062
rect 249996 480 250024 3946
rect 251192 480 251220 4014
rect 252388 480 252416 16546
rect 253584 3602 253612 16546
rect 254676 4140 254728 4146
rect 254676 4082 254728 4088
rect 253480 3596 253532 3602
rect 253480 3538 253532 3544
rect 253572 3596 253624 3602
rect 253572 3538 253624 3544
rect 253492 480 253520 3538
rect 254688 480 254716 4082
rect 255884 480 255912 16546
rect 257068 3936 257120 3942
rect 257068 3878 257120 3884
rect 257080 480 257108 3878
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 258276 480 258304 3810
rect 258736 3398 258764 124743
rect 260116 3602 260144 149058
rect 260208 147422 260236 232358
rect 260300 157826 260328 236982
rect 260576 235414 260604 239770
rect 260656 239760 260708 239766
rect 260656 239702 260708 239708
rect 260838 239728 260894 239737
rect 260564 235408 260616 235414
rect 260564 235350 260616 235356
rect 260472 233640 260524 233646
rect 260472 233582 260524 233588
rect 260378 223544 260434 223553
rect 260378 223479 260434 223488
rect 260392 207641 260420 223479
rect 260484 223310 260512 233582
rect 260668 231854 260696 239702
rect 260838 239663 260840 239672
rect 260892 239663 260894 239672
rect 260840 239634 260892 239640
rect 260840 239556 260892 239562
rect 260840 239498 260892 239504
rect 260748 239488 260800 239494
rect 260748 239430 260800 239436
rect 260760 237425 260788 239430
rect 260746 237416 260802 237425
rect 260746 237351 260802 237360
rect 260852 235124 260880 239498
rect 260944 235278 260972 239788
rect 261036 239788 261110 239816
rect 261622 239838 261674 239844
rect 261714 239896 261766 239902
rect 261714 239838 261766 239844
rect 261528 239799 261584 239808
rect 261818 239816 261846 240108
rect 261910 239970 261938 240108
rect 262002 239970 262030 240108
rect 262094 239970 262122 240108
rect 262186 239970 262214 240108
rect 261898 239964 261950 239970
rect 261898 239906 261950 239912
rect 261990 239964 262042 239970
rect 261990 239906 262042 239912
rect 262082 239964 262134 239970
rect 262082 239906 262134 239912
rect 262174 239964 262226 239970
rect 262174 239906 262226 239912
rect 262034 239864 262090 239873
rect 261944 239828 261996 239834
rect 261818 239788 261892 239816
rect 261036 236881 261064 239788
rect 261484 239760 261536 239766
rect 261484 239702 261536 239708
rect 261576 239760 261628 239766
rect 261576 239702 261628 239708
rect 261668 239760 261720 239766
rect 261864 239748 261892 239788
rect 262034 239799 262090 239808
rect 262128 239828 262180 239834
rect 261944 239770 261996 239776
rect 261668 239702 261720 239708
rect 261772 239720 261892 239748
rect 261300 239692 261352 239698
rect 261300 239634 261352 239640
rect 261312 238610 261340 239634
rect 261392 239556 261444 239562
rect 261392 239498 261444 239504
rect 261300 238604 261352 238610
rect 261300 238546 261352 238552
rect 261022 236872 261078 236881
rect 261022 236807 261078 236816
rect 261208 236360 261260 236366
rect 261208 236302 261260 236308
rect 260932 235272 260984 235278
rect 260932 235214 260984 235220
rect 260852 235096 260972 235124
rect 260840 234728 260892 234734
rect 260840 234670 260892 234676
rect 260576 231826 260696 231854
rect 260576 227730 260604 231826
rect 260564 227724 260616 227730
rect 260564 227666 260616 227672
rect 260472 223304 260524 223310
rect 260472 223246 260524 223252
rect 260484 219434 260512 223246
rect 260852 221474 260880 234670
rect 260944 227526 260972 235096
rect 261220 232694 261248 236302
rect 261208 232688 261260 232694
rect 261208 232630 261260 232636
rect 261404 229094 261432 239498
rect 261496 237318 261524 239702
rect 261484 237312 261536 237318
rect 261484 237254 261536 237260
rect 261484 236020 261536 236026
rect 261484 235962 261536 235968
rect 261496 229809 261524 235962
rect 261588 234734 261616 239702
rect 261680 235346 261708 239702
rect 261668 235340 261720 235346
rect 261668 235282 261720 235288
rect 261576 234728 261628 234734
rect 261576 234670 261628 234676
rect 261574 233608 261630 233617
rect 261574 233543 261630 233552
rect 261588 231810 261616 233543
rect 261576 231804 261628 231810
rect 261576 231746 261628 231752
rect 261482 229800 261538 229809
rect 261482 229735 261538 229744
rect 261404 229066 261524 229094
rect 260932 227520 260984 227526
rect 260932 227462 260984 227468
rect 260944 226370 260972 227462
rect 260932 226364 260984 226370
rect 260932 226306 260984 226312
rect 260840 221468 260892 221474
rect 260840 221410 260892 221416
rect 260484 219406 260788 219434
rect 260378 207632 260434 207641
rect 260378 207567 260434 207576
rect 260760 171134 260788 219406
rect 261496 176089 261524 229066
rect 261482 176080 261538 176089
rect 261482 176015 261538 176024
rect 260392 171106 260788 171134
rect 260392 169794 260420 171106
rect 260380 169788 260432 169794
rect 260380 169730 260432 169736
rect 260288 157820 260340 157826
rect 260288 157762 260340 157768
rect 260196 147416 260248 147422
rect 260196 147358 260248 147364
rect 260392 144634 260420 169730
rect 260380 144628 260432 144634
rect 260380 144570 260432 144576
rect 261484 142928 261536 142934
rect 261484 142870 261536 142876
rect 260838 142216 260894 142225
rect 260838 142151 260840 142160
rect 260892 142151 260894 142160
rect 260840 142122 260892 142128
rect 260656 4004 260708 4010
rect 260656 3946 260708 3952
rect 260012 3596 260064 3602
rect 260012 3538 260064 3544
rect 260104 3596 260156 3602
rect 260104 3538 260156 3544
rect 260024 3398 260052 3538
rect 258724 3392 258776 3398
rect 258724 3334 258776 3340
rect 259460 3392 259512 3398
rect 259460 3334 259512 3340
rect 260012 3392 260064 3398
rect 260012 3334 260064 3340
rect 259472 480 259500 3334
rect 260668 480 260696 3946
rect 261496 3874 261524 142870
rect 261588 140690 261616 231746
rect 261772 231577 261800 239720
rect 261956 236609 261984 239770
rect 262048 239766 262076 239799
rect 262278 239816 262306 240108
rect 262370 239970 262398 240108
rect 262462 239970 262490 240108
rect 262358 239964 262410 239970
rect 262358 239906 262410 239912
rect 262450 239964 262502 239970
rect 262450 239906 262502 239912
rect 262554 239850 262582 240108
rect 262646 239873 262674 240108
rect 262404 239828 262456 239834
rect 262278 239788 262352 239816
rect 262128 239770 262180 239776
rect 262036 239760 262088 239766
rect 262036 239702 262088 239708
rect 262140 239193 262168 239770
rect 262218 239728 262274 239737
rect 262218 239663 262220 239672
rect 262272 239663 262274 239672
rect 262220 239634 262272 239640
rect 262232 239465 262260 239634
rect 262218 239456 262274 239465
rect 262218 239391 262274 239400
rect 262126 239184 262182 239193
rect 262126 239119 262182 239128
rect 262036 237992 262088 237998
rect 262036 237934 262088 237940
rect 261942 236600 261998 236609
rect 261942 236535 261998 236544
rect 261758 231568 261814 231577
rect 261758 231503 261760 231512
rect 261812 231503 261814 231512
rect 261760 231474 261812 231480
rect 261772 231443 261800 231474
rect 262048 226846 262076 237934
rect 262324 234938 262352 239788
rect 262404 239770 262456 239776
rect 262508 239822 262582 239850
rect 262632 239864 262688 239873
rect 262312 234932 262364 234938
rect 262312 234874 262364 234880
rect 262416 231962 262444 239770
rect 262508 237017 262536 239822
rect 262738 239850 262766 240108
rect 262830 239970 262858 240108
rect 262922 239970 262950 240108
rect 263014 239970 263042 240108
rect 262818 239964 262870 239970
rect 262818 239906 262870 239912
rect 262910 239964 262962 239970
rect 262910 239906 262962 239912
rect 263002 239964 263054 239970
rect 263002 239906 263054 239912
rect 263106 239873 263134 240108
rect 263198 239902 263226 240108
rect 263290 239970 263318 240108
rect 263382 239970 263410 240108
rect 263278 239964 263330 239970
rect 263278 239906 263330 239912
rect 263370 239964 263422 239970
rect 263370 239906 263422 239912
rect 263186 239896 263238 239902
rect 263092 239864 263148 239873
rect 262738 239822 262812 239850
rect 262632 239799 262688 239808
rect 262678 239728 262734 239737
rect 262678 239663 262734 239672
rect 262692 239562 262720 239663
rect 262680 239556 262732 239562
rect 262680 239498 262732 239504
rect 262784 239465 262812 239822
rect 262956 239828 263008 239834
rect 263186 239838 263238 239844
rect 263322 239864 263378 239873
rect 263092 239799 263148 239808
rect 263474 239816 263502 240108
rect 263566 239907 263594 240108
rect 263552 239898 263608 239907
rect 263552 239833 263608 239842
rect 263322 239799 263378 239808
rect 262956 239770 263008 239776
rect 262864 239692 262916 239698
rect 262864 239634 262916 239640
rect 262770 239456 262826 239465
rect 262770 239391 262826 239400
rect 262772 238876 262824 238882
rect 262772 238818 262824 238824
rect 262494 237008 262550 237017
rect 262494 236943 262550 236952
rect 262784 234614 262812 238818
rect 262876 234682 262904 239634
rect 262968 238921 262996 239770
rect 263048 239760 263100 239766
rect 263048 239702 263100 239708
rect 262954 238912 263010 238921
rect 262954 238847 263010 238856
rect 262956 238808 263008 238814
rect 262954 238776 262956 238785
rect 263008 238776 263010 238785
rect 262954 238711 263010 238720
rect 263060 234802 263088 239702
rect 263232 239692 263284 239698
rect 263232 239634 263284 239640
rect 263140 239624 263192 239630
rect 263140 239566 263192 239572
rect 263048 234796 263100 234802
rect 263048 234738 263100 234744
rect 262876 234654 262996 234682
rect 262784 234586 262904 234614
rect 262232 231934 262444 231962
rect 262036 226840 262088 226846
rect 262036 226782 262088 226788
rect 262232 223553 262260 231934
rect 262404 231804 262456 231810
rect 262404 231746 262456 231752
rect 262496 231804 262548 231810
rect 262496 231746 262548 231752
rect 262416 231538 262444 231746
rect 262404 231532 262456 231538
rect 262404 231474 262456 231480
rect 262508 231334 262536 231746
rect 262496 231328 262548 231334
rect 262496 231270 262548 231276
rect 262312 231192 262364 231198
rect 262312 231134 262364 231140
rect 262218 223544 262274 223553
rect 262218 223479 262274 223488
rect 262324 173194 262352 231134
rect 262876 229566 262904 234586
rect 262864 229560 262916 229566
rect 262864 229502 262916 229508
rect 262864 227792 262916 227798
rect 262864 227734 262916 227740
rect 262312 173188 262364 173194
rect 262312 173130 262364 173136
rect 262876 152833 262904 227734
rect 262968 227662 262996 234654
rect 263152 233073 263180 239566
rect 263138 233064 263194 233073
rect 263138 232999 263194 233008
rect 263152 229094 263180 232999
rect 263244 231198 263272 239634
rect 263336 235754 263364 239799
rect 263428 239788 263502 239816
rect 263324 235748 263376 235754
rect 263324 235690 263376 235696
rect 263232 231192 263284 231198
rect 263232 231134 263284 231140
rect 263060 229066 263180 229094
rect 263428 229072 263456 239788
rect 263658 239748 263686 240108
rect 263750 239816 263778 240108
rect 263842 239970 263870 240108
rect 263830 239964 263882 239970
rect 263830 239906 263882 239912
rect 263934 239816 263962 240108
rect 264026 239970 264054 240108
rect 264014 239964 264066 239970
rect 264014 239906 264066 239912
rect 264118 239816 264146 240108
rect 264210 239850 264238 240108
rect 264302 239970 264330 240108
rect 264394 239970 264422 240108
rect 264290 239964 264342 239970
rect 264290 239906 264342 239912
rect 264382 239964 264434 239970
rect 264382 239906 264434 239912
rect 264486 239873 264514 240108
rect 264472 239864 264528 239873
rect 264210 239822 264284 239850
rect 263750 239788 263824 239816
rect 263934 239788 264008 239816
rect 263658 239720 263732 239748
rect 263508 239692 263560 239698
rect 263508 239634 263560 239640
rect 263520 236366 263548 239634
rect 263600 239488 263652 239494
rect 263600 239430 263652 239436
rect 263508 236360 263560 236366
rect 263508 236302 263560 236308
rect 263508 234728 263560 234734
rect 263508 234670 263560 234676
rect 262956 227656 263008 227662
rect 262956 227598 263008 227604
rect 262968 154193 262996 227598
rect 263060 159089 263088 229066
rect 263244 229044 263456 229072
rect 263244 227594 263272 229044
rect 263520 228954 263548 234670
rect 263508 228948 263560 228954
rect 263508 228890 263560 228896
rect 263520 227798 263548 228890
rect 263508 227792 263560 227798
rect 263508 227734 263560 227740
rect 263232 227588 263284 227594
rect 263232 227530 263284 227536
rect 263138 223272 263194 223281
rect 263138 223207 263194 223216
rect 263152 161945 263180 223207
rect 263244 207806 263272 227530
rect 263322 223544 263378 223553
rect 263322 223479 263378 223488
rect 263336 223145 263364 223479
rect 263322 223136 263378 223145
rect 263322 223071 263378 223080
rect 263232 207800 263284 207806
rect 263232 207742 263284 207748
rect 263336 206310 263364 223071
rect 263324 206304 263376 206310
rect 263324 206246 263376 206252
rect 263612 167657 263640 239430
rect 263704 237153 263732 239720
rect 263690 237144 263746 237153
rect 263690 237079 263746 237088
rect 263796 234734 263824 239788
rect 263876 239692 263928 239698
rect 263876 239634 263928 239640
rect 263888 238513 263916 239634
rect 263980 238728 264008 239788
rect 264072 239788 264146 239816
rect 264072 238796 264100 239788
rect 264256 239329 264284 239822
rect 264336 239828 264388 239834
rect 264578 239850 264606 240108
rect 264670 239970 264698 240108
rect 264658 239964 264710 239970
rect 264658 239906 264710 239912
rect 264578 239822 264652 239850
rect 264472 239799 264528 239808
rect 264336 239770 264388 239776
rect 264242 239320 264298 239329
rect 264242 239255 264298 239264
rect 264348 238864 264376 239770
rect 264520 239760 264572 239766
rect 264520 239702 264572 239708
rect 264428 239692 264480 239698
rect 264428 239634 264480 239640
rect 264440 239057 264468 239634
rect 264426 239048 264482 239057
rect 264426 238983 264482 238992
rect 264256 238836 264376 238864
rect 264072 238768 264192 238796
rect 263980 238700 264100 238728
rect 263966 238640 264022 238649
rect 263966 238575 264022 238584
rect 263874 238504 263930 238513
rect 263874 238439 263930 238448
rect 263876 238196 263928 238202
rect 263876 238138 263928 238144
rect 263888 237862 263916 238138
rect 263980 238105 264008 238575
rect 263966 238096 264022 238105
rect 263966 238031 264022 238040
rect 263876 237856 263928 237862
rect 263876 237798 263928 237804
rect 264072 237726 264100 238700
rect 264060 237720 264112 237726
rect 264060 237662 264112 237668
rect 263876 235136 263928 235142
rect 263876 235078 263928 235084
rect 263784 234728 263836 234734
rect 263784 234670 263836 234676
rect 263888 233753 263916 235078
rect 263874 233744 263930 233753
rect 263874 233679 263930 233688
rect 263692 233572 263744 233578
rect 263692 233514 263744 233520
rect 263704 170377 263732 233514
rect 264164 230217 264192 238768
rect 264256 230489 264284 238836
rect 264428 238740 264480 238746
rect 264428 238682 264480 238688
rect 264440 238610 264468 238682
rect 264532 238649 264560 239702
rect 264518 238640 264574 238649
rect 264428 238604 264480 238610
rect 264518 238575 264574 238584
rect 264428 238546 264480 238552
rect 264532 233578 264560 238575
rect 264520 233572 264572 233578
rect 264520 233514 264572 233520
rect 264520 231872 264572 231878
rect 264520 231814 264572 231820
rect 264532 231198 264560 231814
rect 264520 231192 264572 231198
rect 264520 231134 264572 231140
rect 264242 230480 264298 230489
rect 264242 230415 264298 230424
rect 264150 230208 264206 230217
rect 264150 230143 264206 230152
rect 264164 223922 264192 230143
rect 264256 229094 264284 230415
rect 264256 229066 264376 229094
rect 264348 224074 264376 229066
rect 264624 227225 264652 239822
rect 264762 239816 264790 240108
rect 264854 239902 264882 240108
rect 264842 239896 264894 239902
rect 264842 239838 264894 239844
rect 264946 239850 264974 240108
rect 265038 239970 265066 240108
rect 265026 239964 265078 239970
rect 265026 239906 265078 239912
rect 265130 239902 265158 240108
rect 265222 239902 265250 240108
rect 265314 239902 265342 240108
rect 265118 239896 265170 239902
rect 264946 239822 265020 239850
rect 265118 239838 265170 239844
rect 265210 239896 265262 239902
rect 265210 239838 265262 239844
rect 265302 239896 265354 239902
rect 265406 239873 265434 240108
rect 265302 239838 265354 239844
rect 265392 239864 265448 239873
rect 264716 239788 264790 239816
rect 264716 235482 264744 239788
rect 264796 239692 264848 239698
rect 264796 239634 264848 239640
rect 264704 235476 264756 235482
rect 264704 235418 264756 235424
rect 264808 229094 264836 239634
rect 264888 239624 264940 239630
rect 264888 239566 264940 239572
rect 264900 237833 264928 239566
rect 264992 239494 265020 239822
rect 265392 239799 265448 239808
rect 265498 239816 265526 240108
rect 265590 239970 265618 240108
rect 265578 239964 265630 239970
rect 265578 239906 265630 239912
rect 265498 239788 265572 239816
rect 265544 239748 265572 239788
rect 265682 239748 265710 240108
rect 265774 239970 265802 240108
rect 265762 239964 265814 239970
rect 265762 239906 265814 239912
rect 265760 239864 265816 239873
rect 265866 239850 265894 240108
rect 265958 239902 265986 240108
rect 266050 239907 266078 240108
rect 266142 239970 266170 240108
rect 266130 239964 266182 239970
rect 265816 239822 265894 239850
rect 265946 239896 265998 239902
rect 265946 239838 265998 239844
rect 266036 239898 266092 239907
rect 266130 239906 266182 239912
rect 266234 239850 266262 240108
rect 266326 239970 266354 240108
rect 266314 239964 266366 239970
rect 266314 239906 266366 239912
rect 266418 239902 266446 240108
rect 266510 239902 266538 240108
rect 266036 239833 266092 239842
rect 266188 239822 266262 239850
rect 266406 239896 266458 239902
rect 266406 239838 266458 239844
rect 266498 239896 266550 239902
rect 266602 239873 266630 240108
rect 266694 239970 266722 240108
rect 266682 239964 266734 239970
rect 266682 239906 266734 239912
rect 266498 239838 266550 239844
rect 266588 239864 266644 239873
rect 265760 239799 265816 239808
rect 265452 239720 265572 239748
rect 265636 239720 265710 239748
rect 265900 239760 265952 239766
rect 265072 239692 265124 239698
rect 265124 239652 265204 239680
rect 265072 239634 265124 239640
rect 264980 239488 265032 239494
rect 264980 239430 265032 239436
rect 264992 239057 265020 239430
rect 264978 239048 265034 239057
rect 264978 238983 265034 238992
rect 264980 238808 265032 238814
rect 264978 238776 264980 238785
rect 265032 238776 265034 238785
rect 264978 238711 265034 238720
rect 264886 237824 264942 237833
rect 264886 237759 264942 237768
rect 265176 234734 265204 239652
rect 265256 239488 265308 239494
rect 265256 239430 265308 239436
rect 265268 238649 265296 239430
rect 265452 239057 265480 239720
rect 265636 239680 265664 239720
rect 265900 239702 265952 239708
rect 265992 239760 266044 239766
rect 266188 239714 266216 239822
rect 266786 239850 266814 240108
rect 266588 239799 266644 239808
rect 266740 239822 266814 239850
rect 266878 239850 266906 240108
rect 266970 239970 266998 240108
rect 267062 239970 267090 240108
rect 266958 239964 267010 239970
rect 266958 239906 267010 239912
rect 267050 239964 267102 239970
rect 267050 239906 267102 239912
rect 267154 239902 267182 240108
rect 267142 239896 267194 239902
rect 266878 239822 266952 239850
rect 267246 239884 267274 240108
rect 267338 239952 267366 240108
rect 267338 239924 267596 239952
rect 267246 239856 267504 239884
rect 267142 239838 267194 239844
rect 265992 239702 266044 239708
rect 265544 239652 265664 239680
rect 265438 239048 265494 239057
rect 265438 238983 265494 238992
rect 265254 238640 265310 238649
rect 265254 238575 265310 238584
rect 265268 236026 265296 238575
rect 265256 236020 265308 236026
rect 265256 235962 265308 235968
rect 265164 234728 265216 234734
rect 265164 234670 265216 234676
rect 265452 230738 265480 238983
rect 265544 238785 265572 239652
rect 265808 239556 265860 239562
rect 265808 239498 265860 239504
rect 265714 239320 265770 239329
rect 265714 239255 265770 239264
rect 265530 238776 265586 238785
rect 265530 238711 265586 238720
rect 264716 229066 264836 229094
rect 265084 230710 265480 230738
rect 264716 228682 264744 229066
rect 264704 228676 264756 228682
rect 264704 228618 264756 228624
rect 264716 227497 264744 228618
rect 264702 227488 264758 227497
rect 264702 227423 264758 227432
rect 264610 227216 264666 227225
rect 264610 227151 264666 227160
rect 264256 224046 264376 224074
rect 264152 223916 264204 223922
rect 264152 223858 264204 223864
rect 263690 170368 263746 170377
rect 263690 170303 263746 170312
rect 263598 167648 263654 167657
rect 263598 167583 263654 167592
rect 263138 161936 263194 161945
rect 263138 161871 263194 161880
rect 264256 161265 264284 224046
rect 264624 223990 264652 227151
rect 264336 223984 264388 223990
rect 264336 223926 264388 223932
rect 264612 223984 264664 223990
rect 264612 223926 264664 223932
rect 264348 207738 264376 223926
rect 264428 223916 264480 223922
rect 264428 223858 264480 223864
rect 264336 207732 264388 207738
rect 264336 207674 264388 207680
rect 264440 164937 264468 223858
rect 265084 165073 265112 230710
rect 265440 230648 265492 230654
rect 265440 230590 265492 230596
rect 265070 165064 265126 165073
rect 265070 164999 265126 165008
rect 264426 164928 264482 164937
rect 264426 164863 264482 164872
rect 264242 161256 264298 161265
rect 264242 161191 264298 161200
rect 263046 159080 263102 159089
rect 263046 159015 263102 159024
rect 262954 154184 263010 154193
rect 262954 154119 263010 154128
rect 262862 152824 262918 152833
rect 262862 152759 262918 152768
rect 264244 147416 264296 147422
rect 264244 147358 264296 147364
rect 263598 142896 263654 142905
rect 263598 142831 263600 142840
rect 263652 142831 263654 142840
rect 263600 142802 263652 142808
rect 261576 140684 261628 140690
rect 261576 140626 261628 140632
rect 261588 126342 261616 140626
rect 261576 126336 261628 126342
rect 261576 126278 261628 126284
rect 262220 111104 262272 111110
rect 262220 111046 262272 111052
rect 262232 16574 262260 111046
rect 262232 16546 262536 16574
rect 261484 3868 261536 3874
rect 261484 3810 261536 3816
rect 261760 3596 261812 3602
rect 261760 3538 261812 3544
rect 261772 480 261800 3538
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264256 3942 264284 147358
rect 265452 144362 265480 230590
rect 265544 226914 265572 238711
rect 265728 237289 265756 239255
rect 265820 238785 265848 239498
rect 265806 238776 265862 238785
rect 265806 238711 265862 238720
rect 265912 238377 265940 239702
rect 266004 238610 266032 239702
rect 266096 239686 266216 239714
rect 266268 239760 266320 239766
rect 266268 239702 266320 239708
rect 266360 239760 266412 239766
rect 266360 239702 266412 239708
rect 266544 239760 266596 239766
rect 266636 239760 266688 239766
rect 266544 239702 266596 239708
rect 266634 239728 266636 239737
rect 266688 239728 266690 239737
rect 266096 239562 266124 239686
rect 266176 239624 266228 239630
rect 266176 239566 266228 239572
rect 266084 239556 266136 239562
rect 266084 239498 266136 239504
rect 266082 239320 266138 239329
rect 266082 239255 266138 239264
rect 265992 238604 266044 238610
rect 265992 238546 266044 238552
rect 265898 238368 265954 238377
rect 265898 238303 265954 238312
rect 265808 238128 265860 238134
rect 265808 238070 265860 238076
rect 265820 237969 265848 238070
rect 265806 237960 265862 237969
rect 265806 237895 265862 237904
rect 265714 237280 265770 237289
rect 265714 237215 265770 237224
rect 265808 234864 265860 234870
rect 265808 234806 265860 234812
rect 265716 234728 265768 234734
rect 265716 234670 265768 234676
rect 265728 228857 265756 234670
rect 265714 228848 265770 228857
rect 265624 228812 265676 228818
rect 265714 228783 265770 228792
rect 265624 228754 265676 228760
rect 265532 226908 265584 226914
rect 265532 226850 265584 226856
rect 265636 161401 265664 228754
rect 265728 226794 265756 228783
rect 265820 226914 265848 234806
rect 265912 230654 265940 238303
rect 265992 236020 266044 236026
rect 265992 235962 266044 235968
rect 265900 230648 265952 230654
rect 265900 230590 265952 230596
rect 265808 226908 265860 226914
rect 265808 226850 265860 226856
rect 265728 226766 265848 226794
rect 265716 226704 265768 226710
rect 265716 226646 265768 226652
rect 265728 180033 265756 226646
rect 265820 207670 265848 226766
rect 266004 219434 266032 235962
rect 265912 219406 266032 219434
rect 265808 207664 265860 207670
rect 265808 207606 265860 207612
rect 265714 180024 265770 180033
rect 265714 179959 265770 179968
rect 265912 163441 265940 219406
rect 266096 166297 266124 239255
rect 266188 236026 266216 239566
rect 266176 236020 266228 236026
rect 266176 235962 266228 235968
rect 266176 235680 266228 235686
rect 266176 235622 266228 235628
rect 266188 231266 266216 235622
rect 266176 231260 266228 231266
rect 266176 231202 266228 231208
rect 266280 226710 266308 239702
rect 266372 236638 266400 239702
rect 266360 236632 266412 236638
rect 266360 236574 266412 236580
rect 266372 235249 266400 236574
rect 266358 235240 266414 235249
rect 266358 235175 266414 235184
rect 266452 235204 266504 235210
rect 266452 235146 266504 235152
rect 266360 235136 266412 235142
rect 266360 235078 266412 235084
rect 266268 226704 266320 226710
rect 266268 226646 266320 226652
rect 266280 226234 266308 226646
rect 266268 226228 266320 226234
rect 266268 226170 266320 226176
rect 266372 177342 266400 235078
rect 266464 231266 266492 235146
rect 266452 231260 266504 231266
rect 266452 231202 266504 231208
rect 266556 228410 266584 239702
rect 266634 239663 266690 239672
rect 266636 239488 266688 239494
rect 266634 239456 266636 239465
rect 266688 239456 266690 239465
rect 266634 239391 266690 239400
rect 266636 237992 266688 237998
rect 266636 237934 266688 237940
rect 266544 228404 266596 228410
rect 266544 228346 266596 228352
rect 266648 223574 266676 237934
rect 266740 228993 266768 239822
rect 266820 239760 266872 239766
rect 266820 239702 266872 239708
rect 266832 237998 266860 239702
rect 266924 239698 266952 239822
rect 267004 239828 267056 239834
rect 267004 239770 267056 239776
rect 266912 239692 266964 239698
rect 266912 239634 266964 239640
rect 266924 238513 266952 239634
rect 266910 238504 266966 238513
rect 266910 238439 266966 238448
rect 266820 237992 266872 237998
rect 266820 237934 266872 237940
rect 267016 235142 267044 239770
rect 267372 239624 267424 239630
rect 267372 239566 267424 239572
rect 267278 239320 267334 239329
rect 267278 239255 267334 239264
rect 267292 238474 267320 239255
rect 267280 238468 267332 238474
rect 267280 238410 267332 238416
rect 267384 238270 267412 239566
rect 267372 238264 267424 238270
rect 267372 238206 267424 238212
rect 267188 236088 267240 236094
rect 267188 236030 267240 236036
rect 267004 235136 267056 235142
rect 267004 235078 267056 235084
rect 267200 231334 267228 236030
rect 267476 235929 267504 239856
rect 267568 237998 267596 239924
rect 267646 239864 267702 239873
rect 267646 239799 267702 239808
rect 267556 237992 267608 237998
rect 267556 237934 267608 237940
rect 267556 237380 267608 237386
rect 267556 237322 267608 237328
rect 267462 235920 267518 235929
rect 267462 235855 267518 235864
rect 267476 235686 267504 235855
rect 267464 235680 267516 235686
rect 267464 235622 267516 235628
rect 267188 231328 267240 231334
rect 267094 231296 267150 231305
rect 267188 231270 267240 231276
rect 267094 231231 267150 231240
rect 266726 228984 266782 228993
rect 266726 228919 266782 228928
rect 267002 228984 267058 228993
rect 267002 228919 267058 228928
rect 266648 223546 266768 223574
rect 266360 177336 266412 177342
rect 266360 177278 266412 177284
rect 266740 174593 266768 223546
rect 266726 174584 266782 174593
rect 266726 174519 266782 174528
rect 266082 166288 266138 166297
rect 266082 166223 266138 166232
rect 265898 163432 265954 163441
rect 265898 163367 265954 163376
rect 265622 161392 265678 161401
rect 265622 161327 265678 161336
rect 267016 159225 267044 228919
rect 267108 171737 267136 231231
rect 267188 228404 267240 228410
rect 267188 228346 267240 228352
rect 267200 227497 267228 228346
rect 267186 227488 267242 227497
rect 267186 227423 267242 227432
rect 267200 204921 267228 227423
rect 267568 223574 267596 237322
rect 267476 223546 267596 223574
rect 267186 204912 267242 204921
rect 267186 204847 267242 204856
rect 267476 182889 267504 223546
rect 267462 182880 267518 182889
rect 267462 182815 267518 182824
rect 267094 171728 267150 171737
rect 267094 171663 267150 171672
rect 267660 162081 267688 239799
rect 267752 239748 267780 240128
rect 267844 239902 267872 248386
rect 267924 240508 267976 240514
rect 267924 240450 267976 240456
rect 267936 240106 267964 240450
rect 267924 240100 267976 240106
rect 267924 240042 267976 240048
rect 268028 239970 268056 250543
rect 268292 242072 268344 242078
rect 268292 242014 268344 242020
rect 268108 240916 268160 240922
rect 268108 240858 268160 240864
rect 268120 240417 268148 240858
rect 268106 240408 268162 240417
rect 268106 240343 268162 240352
rect 268108 240236 268160 240242
rect 268108 240178 268160 240184
rect 268016 239964 268068 239970
rect 268016 239906 268068 239912
rect 267832 239896 267884 239902
rect 267832 239838 267884 239844
rect 267752 239720 267872 239748
rect 267740 238264 267792 238270
rect 267740 238206 267792 238212
rect 267646 162072 267702 162081
rect 267646 162007 267702 162016
rect 267002 159216 267058 159225
rect 267002 159151 267058 159160
rect 267004 156664 267056 156670
rect 267004 156606 267056 156612
rect 265440 144356 265492 144362
rect 265440 144298 265492 144304
rect 265622 122224 265678 122233
rect 265622 122159 265678 122168
rect 264244 3936 264296 3942
rect 264244 3878 264296 3884
rect 265348 3800 265400 3806
rect 265348 3742 265400 3748
rect 264152 3392 264204 3398
rect 264152 3334 264204 3340
rect 264164 480 264192 3334
rect 265360 480 265388 3742
rect 265636 3602 265664 122159
rect 267016 3602 267044 156606
rect 267752 141914 267780 238206
rect 267844 237386 267872 239720
rect 268016 238060 268068 238066
rect 268016 238002 268068 238008
rect 267832 237380 267884 237386
rect 267832 237322 267884 237328
rect 267832 236904 267884 236910
rect 267832 236846 267884 236852
rect 267844 148918 267872 236846
rect 267924 235340 267976 235346
rect 267924 235282 267976 235288
rect 267936 235249 267964 235282
rect 267922 235240 267978 235249
rect 267922 235175 267978 235184
rect 267936 155174 267964 235175
rect 268028 234841 268056 238002
rect 268014 234832 268070 234841
rect 268014 234767 268070 234776
rect 268120 223574 268148 240178
rect 268200 239556 268252 239562
rect 268200 239498 268252 239504
rect 268212 228818 268240 239498
rect 268304 237561 268332 242014
rect 268396 238785 268424 287642
rect 268936 286340 268988 286346
rect 268936 286282 268988 286288
rect 268948 277394 268976 286282
rect 269028 284980 269080 284986
rect 269028 284922 269080 284928
rect 268488 277366 268976 277394
rect 268488 239970 268516 277366
rect 268936 254584 268988 254590
rect 268936 254526 268988 254532
rect 268948 253934 268976 254526
rect 268580 253906 268976 253934
rect 268476 239964 268528 239970
rect 268476 239906 268528 239912
rect 268382 238776 268438 238785
rect 268382 238711 268438 238720
rect 268396 238270 268424 238711
rect 268580 238542 268608 253906
rect 268936 251864 268988 251870
rect 268936 251806 268988 251812
rect 268948 249234 268976 251806
rect 268672 249206 268976 249234
rect 268672 243137 268700 249206
rect 268842 247888 268898 247897
rect 268842 247823 268898 247832
rect 268658 243128 268714 243137
rect 268658 243063 268714 243072
rect 268658 242992 268714 243001
rect 268658 242927 268714 242936
rect 268672 240145 268700 242927
rect 268658 240136 268714 240145
rect 268658 240071 268714 240080
rect 268568 238536 268620 238542
rect 268568 238478 268620 238484
rect 268856 238338 268884 247823
rect 268936 242412 268988 242418
rect 268936 242354 268988 242360
rect 268844 238332 268896 238338
rect 268844 238274 268896 238280
rect 268384 238264 268436 238270
rect 268384 238206 268436 238212
rect 268476 238196 268528 238202
rect 268476 238138 268528 238144
rect 268290 237552 268346 237561
rect 268290 237487 268346 237496
rect 268384 236972 268436 236978
rect 268384 236914 268436 236920
rect 268396 236502 268424 236914
rect 268384 236496 268436 236502
rect 268384 236438 268436 236444
rect 268488 234977 268516 238138
rect 268658 238096 268714 238105
rect 268658 238031 268714 238040
rect 268568 237992 268620 237998
rect 268568 237934 268620 237940
rect 268474 234968 268530 234977
rect 268474 234903 268530 234912
rect 268580 231305 268608 237934
rect 268672 232937 268700 238031
rect 268752 237992 268804 237998
rect 268752 237934 268804 237940
rect 268764 234297 268792 237934
rect 268948 237425 268976 242354
rect 268934 237416 268990 237425
rect 268934 237351 268990 237360
rect 269040 236026 269068 284922
rect 269118 247752 269174 247761
rect 269118 247687 269174 247696
rect 269132 239698 269160 247687
rect 269304 246356 269356 246362
rect 269304 246298 269356 246304
rect 269212 242208 269264 242214
rect 269212 242150 269264 242156
rect 269224 240689 269252 242150
rect 269210 240680 269266 240689
rect 269210 240615 269266 240624
rect 269210 240408 269266 240417
rect 269210 240343 269266 240352
rect 269224 240174 269252 240343
rect 269212 240168 269264 240174
rect 269212 240110 269264 240116
rect 269212 239964 269264 239970
rect 269212 239906 269264 239912
rect 269120 239692 269172 239698
rect 269120 239634 269172 239640
rect 269224 238746 269252 239906
rect 269316 239630 269344 246298
rect 269396 241664 269448 241670
rect 269396 241606 269448 241612
rect 269304 239624 269356 239630
rect 269304 239566 269356 239572
rect 269212 238740 269264 238746
rect 269212 238682 269264 238688
rect 269120 237924 269172 237930
rect 269120 237866 269172 237872
rect 269132 237386 269160 237866
rect 269120 237380 269172 237386
rect 269120 237322 269172 237328
rect 269028 236020 269080 236026
rect 269028 235962 269080 235968
rect 268936 235748 268988 235754
rect 268936 235690 268988 235696
rect 269028 235748 269080 235754
rect 269028 235690 269080 235696
rect 268948 235346 268976 235690
rect 268936 235340 268988 235346
rect 268936 235282 268988 235288
rect 269040 234938 269068 235690
rect 269120 235272 269172 235278
rect 269120 235214 269172 235220
rect 269028 234932 269080 234938
rect 269028 234874 269080 234880
rect 268750 234288 268806 234297
rect 268750 234223 268806 234232
rect 268658 232928 268714 232937
rect 268658 232863 268714 232872
rect 268566 231296 268622 231305
rect 268566 231231 268622 231240
rect 268200 228812 268252 228818
rect 268200 228754 268252 228760
rect 268028 223546 268148 223574
rect 268028 158953 268056 223546
rect 268014 158944 268070 158953
rect 268014 158879 268070 158888
rect 267924 155168 267976 155174
rect 267924 155110 267976 155116
rect 269040 153066 269068 234874
rect 269132 158914 269160 235214
rect 269224 160857 269252 238682
rect 269304 238468 269356 238474
rect 269304 238410 269356 238416
rect 269316 232422 269344 238410
rect 269408 237522 269436 241606
rect 269488 241596 269540 241602
rect 269488 241538 269540 241544
rect 269500 237590 269528 241538
rect 269592 239601 269620 315959
rect 269670 308680 269726 308689
rect 269670 308615 269726 308624
rect 269578 239592 269634 239601
rect 269578 239527 269634 239536
rect 269580 238876 269632 238882
rect 269580 238818 269632 238824
rect 269488 237584 269540 237590
rect 269488 237526 269540 237532
rect 269396 237516 269448 237522
rect 269396 237458 269448 237464
rect 269592 237425 269620 238818
rect 269394 237416 269450 237425
rect 269394 237351 269450 237360
rect 269578 237416 269634 237425
rect 269578 237351 269634 237360
rect 269304 232416 269356 232422
rect 269304 232358 269356 232364
rect 269408 227050 269436 237351
rect 269684 231810 269712 308615
rect 269672 231804 269724 231810
rect 269672 231746 269724 231752
rect 269396 227044 269448 227050
rect 269396 226986 269448 226992
rect 269776 226273 269804 319194
rect 269868 317393 269896 389846
rect 269948 385212 270000 385218
rect 269948 385154 270000 385160
rect 269854 317384 269910 317393
rect 269854 317319 269910 317328
rect 269854 315752 269910 315761
rect 269854 315687 269910 315696
rect 269868 229770 269896 315687
rect 269960 302190 269988 385154
rect 270052 320521 270080 396743
rect 270038 320512 270094 320521
rect 270038 320447 270094 320456
rect 270040 317756 270092 317762
rect 270040 317698 270092 317704
rect 269948 302184 270000 302190
rect 269948 302126 270000 302132
rect 269948 257372 270000 257378
rect 269948 257314 270000 257320
rect 269960 234569 269988 257314
rect 270052 240825 270080 317698
rect 270144 317354 270172 396879
rect 271512 396840 271564 396846
rect 271512 396782 271564 396788
rect 270222 396672 270278 396681
rect 270222 396607 270278 396616
rect 270132 317348 270184 317354
rect 270132 317290 270184 317296
rect 270144 316878 270172 317290
rect 270132 316872 270184 316878
rect 270132 316814 270184 316820
rect 270236 314294 270264 396607
rect 271234 395312 271290 395321
rect 271234 395247 271290 395256
rect 270406 394088 270462 394097
rect 270406 394023 270462 394032
rect 270316 391332 270368 391338
rect 270316 391274 270368 391280
rect 270224 314288 270276 314294
rect 270224 314230 270276 314236
rect 270236 313342 270264 314230
rect 270224 313336 270276 313342
rect 270224 313278 270276 313284
rect 270130 311672 270186 311681
rect 270130 311607 270186 311616
rect 270038 240816 270094 240825
rect 270038 240751 270094 240760
rect 270144 235074 270172 311607
rect 270328 310162 270356 391274
rect 270420 310321 270448 394023
rect 271248 325694 271276 395247
rect 271420 392624 271472 392630
rect 271420 392566 271472 392572
rect 271328 370456 271380 370462
rect 271328 370398 271380 370404
rect 271064 325666 271276 325694
rect 271064 320346 271092 325666
rect 271142 320376 271198 320385
rect 271052 320340 271104 320346
rect 271142 320311 271198 320320
rect 271052 320282 271104 320288
rect 271064 315897 271092 320282
rect 271050 315888 271106 315897
rect 271050 315823 271106 315832
rect 270684 313336 270736 313342
rect 270684 313278 270736 313284
rect 270406 310312 270462 310321
rect 270406 310247 270462 310256
rect 270328 310134 270448 310162
rect 270420 309058 270448 310134
rect 270408 309052 270460 309058
rect 270408 308994 270460 309000
rect 270420 308650 270448 308994
rect 270408 308644 270460 308650
rect 270408 308586 270460 308592
rect 270222 257544 270278 257553
rect 270222 257479 270278 257488
rect 270236 247034 270264 257479
rect 270236 247006 270356 247034
rect 270222 241632 270278 241641
rect 270222 241567 270278 241576
rect 270236 241534 270264 241567
rect 270224 241528 270276 241534
rect 270224 241470 270276 241476
rect 270328 238241 270356 247006
rect 270406 246392 270462 246401
rect 270406 246327 270462 246336
rect 270420 238377 270448 246327
rect 270592 243704 270644 243710
rect 270592 243646 270644 243652
rect 270498 240136 270554 240145
rect 270498 240071 270554 240080
rect 270512 240038 270540 240071
rect 270500 240032 270552 240038
rect 270500 239974 270552 239980
rect 270406 238368 270462 238377
rect 270406 238303 270462 238312
rect 270314 238232 270370 238241
rect 270314 238167 270370 238176
rect 270316 237924 270368 237930
rect 270316 237866 270368 237872
rect 270328 237726 270356 237866
rect 270316 237720 270368 237726
rect 270316 237662 270368 237668
rect 270224 235612 270276 235618
rect 270224 235554 270276 235560
rect 270132 235068 270184 235074
rect 270132 235010 270184 235016
rect 270132 234796 270184 234802
rect 270132 234738 270184 234744
rect 269946 234560 270002 234569
rect 269946 234495 270002 234504
rect 270144 234025 270172 234738
rect 270130 234016 270186 234025
rect 270130 233951 270186 233960
rect 269856 229764 269908 229770
rect 269856 229706 269908 229712
rect 269762 226264 269818 226273
rect 269762 226199 269818 226208
rect 270144 161474 270172 233951
rect 269776 161446 270172 161474
rect 269210 160848 269266 160857
rect 269210 160783 269266 160792
rect 269120 158908 269172 158914
rect 269120 158850 269172 158856
rect 269776 155990 269804 161446
rect 270236 159202 270264 235554
rect 270052 159174 270264 159202
rect 269764 155984 269816 155990
rect 269764 155926 269816 155932
rect 269120 154148 269172 154154
rect 269120 154090 269172 154096
rect 269028 153060 269080 153066
rect 269028 153002 269080 153008
rect 269040 152590 269068 153002
rect 269028 152584 269080 152590
rect 269028 152526 269080 152532
rect 267832 148912 267884 148918
rect 267832 148854 267884 148860
rect 268384 148912 268436 148918
rect 268384 148854 268436 148860
rect 267740 141908 267792 141914
rect 267740 141850 267792 141856
rect 267740 3936 267792 3942
rect 267740 3878 267792 3884
rect 265624 3596 265676 3602
rect 265624 3538 265676 3544
rect 266544 3596 266596 3602
rect 266544 3538 266596 3544
rect 267004 3596 267056 3602
rect 267004 3538 267056 3544
rect 266556 480 266584 3538
rect 267752 480 267780 3878
rect 268396 3806 268424 148854
rect 269132 148753 269160 154090
rect 269118 148744 269174 148753
rect 269118 148679 269174 148688
rect 269776 148617 269804 155926
rect 270052 154154 270080 159174
rect 270224 158908 270276 158914
rect 270224 158850 270276 158856
rect 270236 155310 270264 158850
rect 270224 155304 270276 155310
rect 270224 155246 270276 155252
rect 270040 154148 270092 154154
rect 270040 154090 270092 154096
rect 270052 153338 270080 154090
rect 270040 153332 270092 153338
rect 270040 153274 270092 153280
rect 269762 148608 269818 148617
rect 269762 148543 269818 148552
rect 270328 144702 270356 237662
rect 270408 237380 270460 237386
rect 270408 237322 270460 237328
rect 270316 144696 270368 144702
rect 270316 144638 270368 144644
rect 270328 144226 270356 144638
rect 270316 144220 270368 144226
rect 270316 144162 270368 144168
rect 269028 141908 269080 141914
rect 269028 141850 269080 141856
rect 269040 141438 269068 141850
rect 269028 141432 269080 141438
rect 269028 141374 269080 141380
rect 270420 129742 270448 237322
rect 270512 135250 270540 239974
rect 270604 237969 270632 243646
rect 270590 237960 270646 237969
rect 270590 237895 270646 237904
rect 270592 237856 270644 237862
rect 270592 237798 270644 237804
rect 270604 157049 270632 237798
rect 270696 231849 270724 313278
rect 270774 245440 270830 245449
rect 270774 245375 270830 245384
rect 270788 238406 270816 245375
rect 271052 241188 271104 241194
rect 271052 241130 271104 241136
rect 270866 240816 270922 240825
rect 271064 240786 271092 241130
rect 270866 240751 270922 240760
rect 271052 240780 271104 240786
rect 270880 239057 270908 240751
rect 271052 240722 271104 240728
rect 270960 239760 271012 239766
rect 270960 239702 271012 239708
rect 270866 239048 270922 239057
rect 270866 238983 270922 238992
rect 270972 238678 271000 239702
rect 270960 238672 271012 238678
rect 270960 238614 271012 238620
rect 271052 238672 271104 238678
rect 271052 238614 271104 238620
rect 270868 238604 270920 238610
rect 270868 238546 270920 238552
rect 270776 238400 270828 238406
rect 270776 238342 270828 238348
rect 270880 238241 270908 238546
rect 270866 238232 270922 238241
rect 270866 238167 270922 238176
rect 270774 236736 270830 236745
rect 270774 236671 270830 236680
rect 270788 236366 270816 236671
rect 270776 236360 270828 236366
rect 270776 236302 270828 236308
rect 270682 231840 270738 231849
rect 270682 231775 270738 231784
rect 270590 157040 270646 157049
rect 270590 156975 270646 156984
rect 270788 155145 270816 236302
rect 270880 158817 270908 238167
rect 271064 237454 271092 238614
rect 271052 237448 271104 237454
rect 271052 237390 271104 237396
rect 271156 232490 271184 320311
rect 271236 318096 271288 318102
rect 271236 318038 271288 318044
rect 271248 242418 271276 318038
rect 271340 292398 271368 370398
rect 271432 317257 271460 392566
rect 271524 319258 271552 396782
rect 271604 392488 271656 392494
rect 271604 392430 271656 392436
rect 271512 319252 271564 319258
rect 271512 319194 271564 319200
rect 271418 317248 271474 317257
rect 271418 317183 271474 317192
rect 271432 314022 271460 317183
rect 271616 314537 271644 392430
rect 271602 314528 271658 314537
rect 271602 314463 271658 314472
rect 271420 314016 271472 314022
rect 271420 313958 271472 313964
rect 271616 313857 271644 314463
rect 271602 313848 271658 313857
rect 271602 313783 271658 313792
rect 271708 311817 271736 400386
rect 274272 400240 274324 400246
rect 274272 400182 274324 400188
rect 274178 397080 274234 397089
rect 274178 397015 274234 397024
rect 272890 395584 272946 395593
rect 272890 395519 272946 395528
rect 271786 395448 271842 395457
rect 271786 395383 271842 395392
rect 271694 311808 271750 311817
rect 271694 311743 271750 311752
rect 271696 310548 271748 310554
rect 271696 310490 271748 310496
rect 271328 292392 271380 292398
rect 271328 292334 271380 292340
rect 271328 283620 271380 283626
rect 271328 283562 271380 283568
rect 271236 242412 271288 242418
rect 271236 242354 271288 242360
rect 271236 242276 271288 242282
rect 271236 242218 271288 242224
rect 271248 240378 271276 242218
rect 271340 241670 271368 283562
rect 271420 282192 271472 282198
rect 271420 282134 271472 282140
rect 271328 241664 271380 241670
rect 271328 241606 271380 241612
rect 271432 241482 271460 282134
rect 271512 280832 271564 280838
rect 271512 280774 271564 280780
rect 271524 241602 271552 280774
rect 271604 279472 271656 279478
rect 271604 279414 271656 279420
rect 271616 242078 271644 279414
rect 271604 242072 271656 242078
rect 271604 242014 271656 242020
rect 271708 241641 271736 310490
rect 271800 304842 271828 395383
rect 272616 394052 272668 394058
rect 272616 393994 272668 394000
rect 272524 382560 272576 382566
rect 272524 382502 272576 382508
rect 272432 320136 272484 320142
rect 272432 320078 272484 320084
rect 272444 319054 272472 320078
rect 272432 319048 272484 319054
rect 272432 318990 272484 318996
rect 272444 318238 272472 318990
rect 272432 318232 272484 318238
rect 272432 318174 272484 318180
rect 271788 304836 271840 304842
rect 271788 304778 271840 304784
rect 271800 304570 271828 304778
rect 271788 304564 271840 304570
rect 271788 304506 271840 304512
rect 271972 292188 272024 292194
rect 271972 292130 272024 292136
rect 271880 291712 271932 291718
rect 271880 291654 271932 291660
rect 271892 291242 271920 291654
rect 271880 291236 271932 291242
rect 271880 291178 271932 291184
rect 271788 250504 271840 250510
rect 271788 250446 271840 250452
rect 271694 241632 271750 241641
rect 271512 241596 271564 241602
rect 271694 241567 271750 241576
rect 271512 241538 271564 241544
rect 271432 241454 271644 241482
rect 271420 241392 271472 241398
rect 271420 241334 271472 241340
rect 271328 241324 271380 241330
rect 271328 241266 271380 241272
rect 271340 240854 271368 241266
rect 271432 240922 271460 241334
rect 271512 241120 271564 241126
rect 271512 241062 271564 241068
rect 271420 240916 271472 240922
rect 271420 240858 271472 240864
rect 271328 240848 271380 240854
rect 271328 240790 271380 240796
rect 271236 240372 271288 240378
rect 271236 240314 271288 240320
rect 271234 239320 271290 239329
rect 271234 239255 271290 239264
rect 271248 237794 271276 239255
rect 271524 238474 271552 241062
rect 271512 238468 271564 238474
rect 271512 238410 271564 238416
rect 271236 237788 271288 237794
rect 271236 237730 271288 237736
rect 271616 237658 271644 241454
rect 271696 240984 271748 240990
rect 271696 240926 271748 240932
rect 271604 237652 271656 237658
rect 271604 237594 271656 237600
rect 271708 237425 271736 240926
rect 271694 237416 271750 237425
rect 271694 237351 271750 237360
rect 271236 235340 271288 235346
rect 271236 235282 271288 235288
rect 271144 232484 271196 232490
rect 271144 232426 271196 232432
rect 271144 229152 271196 229158
rect 271144 229094 271196 229100
rect 270866 158808 270922 158817
rect 270866 158743 270922 158752
rect 270774 155136 270830 155145
rect 270774 155071 270830 155080
rect 271156 143274 271184 229094
rect 271248 155854 271276 235282
rect 271800 234433 271828 250446
rect 271786 234424 271842 234433
rect 271786 234359 271842 234368
rect 271788 233844 271840 233850
rect 271788 233786 271840 233792
rect 271800 233646 271828 233786
rect 271788 233640 271840 233646
rect 271788 233582 271840 233588
rect 271892 228614 271920 291178
rect 271880 228608 271932 228614
rect 271880 228550 271932 228556
rect 271984 228478 272012 292130
rect 272432 291848 272484 291854
rect 272432 291790 272484 291796
rect 272444 291310 272472 291790
rect 272536 291718 272564 382502
rect 272628 320142 272656 393994
rect 272800 374468 272852 374474
rect 272800 374410 272852 374416
rect 272708 374264 272760 374270
rect 272708 374206 272760 374212
rect 272616 320136 272668 320142
rect 272616 320078 272668 320084
rect 272616 318640 272668 318646
rect 272616 318582 272668 318588
rect 272628 318345 272656 318582
rect 272614 318336 272670 318345
rect 272614 318271 272670 318280
rect 272616 318232 272668 318238
rect 272616 318174 272668 318180
rect 272628 315518 272656 318174
rect 272616 315512 272668 315518
rect 272616 315454 272668 315460
rect 272616 313336 272668 313342
rect 272616 313278 272668 313284
rect 272524 291712 272576 291718
rect 272524 291654 272576 291660
rect 272432 291304 272484 291310
rect 272432 291246 272484 291252
rect 272248 291168 272300 291174
rect 272248 291110 272300 291116
rect 272154 243808 272210 243817
rect 272154 243743 272210 243752
rect 272064 241052 272116 241058
rect 272064 240994 272116 241000
rect 272076 237862 272104 240994
rect 272064 237856 272116 237862
rect 272064 237798 272116 237804
rect 272168 237374 272196 243743
rect 272076 237346 272196 237374
rect 271972 228472 272024 228478
rect 271972 228414 272024 228420
rect 271236 155848 271288 155854
rect 271236 155790 271288 155796
rect 271788 155848 271840 155854
rect 271788 155790 271840 155796
rect 271800 155242 271828 155790
rect 271788 155236 271840 155242
rect 271788 155178 271840 155184
rect 271880 148980 271932 148986
rect 271880 148922 271932 148928
rect 271892 148510 271920 148922
rect 271880 148504 271932 148510
rect 271880 148446 271932 148452
rect 271144 143268 271196 143274
rect 271144 143210 271196 143216
rect 270500 135244 270552 135250
rect 270500 135186 270552 135192
rect 270408 129736 270460 129742
rect 270408 129678 270460 129684
rect 270420 129062 270448 129678
rect 270408 129056 270460 129062
rect 270408 128998 270460 129004
rect 269120 94580 269172 94586
rect 269120 94522 269172 94528
rect 269132 16574 269160 94522
rect 269132 16546 270080 16574
rect 268384 3800 268436 3806
rect 268384 3742 268436 3748
rect 268844 3732 268896 3738
rect 268844 3674 268896 3680
rect 268856 480 268884 3674
rect 270052 480 270080 16546
rect 271156 3398 271184 143210
rect 271788 135244 271840 135250
rect 271788 135186 271840 135192
rect 271800 134570 271828 135186
rect 271788 134564 271840 134570
rect 271788 134506 271840 134512
rect 271892 16574 271920 148446
rect 272076 142361 272104 237346
rect 272154 236736 272210 236745
rect 272154 236671 272210 236680
rect 272168 236473 272196 236671
rect 272154 236464 272210 236473
rect 272154 236399 272210 236408
rect 272168 155922 272196 236399
rect 272260 211818 272288 291110
rect 272338 242584 272394 242593
rect 272338 242519 272394 242528
rect 272352 236337 272380 242519
rect 272338 236328 272394 236337
rect 272338 236263 272394 236272
rect 272248 211812 272300 211818
rect 272248 211754 272300 211760
rect 272352 158846 272380 236263
rect 272444 228138 272472 291246
rect 272524 233844 272576 233850
rect 272524 233786 272576 233792
rect 272536 233714 272564 233786
rect 272524 233708 272576 233714
rect 272524 233650 272576 233656
rect 272432 228132 272484 228138
rect 272432 228074 272484 228080
rect 272432 221536 272484 221542
rect 272432 221478 272484 221484
rect 272340 158840 272392 158846
rect 272340 158782 272392 158788
rect 272156 155916 272208 155922
rect 272156 155858 272208 155864
rect 272340 155916 272392 155922
rect 272340 155858 272392 155864
rect 272352 155378 272380 155858
rect 272340 155372 272392 155378
rect 272340 155314 272392 155320
rect 272444 148510 272472 221478
rect 272536 150278 272564 233650
rect 272628 224058 272656 313278
rect 272720 288697 272748 374206
rect 272812 290494 272840 374410
rect 272904 319297 272932 395519
rect 272984 394324 273036 394330
rect 272984 394266 273036 394272
rect 272890 319288 272946 319297
rect 272890 319223 272946 319232
rect 272996 318646 273024 394266
rect 273996 393984 274048 393990
rect 273718 393952 273774 393961
rect 273996 393926 274048 393932
rect 273718 393887 273774 393896
rect 273168 374604 273220 374610
rect 273168 374546 273220 374552
rect 273076 372700 273128 372706
rect 273076 372642 273128 372648
rect 272984 318640 273036 318646
rect 272984 318582 273036 318588
rect 272892 316600 272944 316606
rect 272892 316542 272944 316548
rect 272800 290488 272852 290494
rect 272800 290430 272852 290436
rect 272706 288688 272762 288697
rect 272706 288623 272762 288632
rect 272708 236020 272760 236026
rect 272708 235962 272760 235968
rect 272616 224052 272668 224058
rect 272616 223994 272668 224000
rect 272524 150272 272576 150278
rect 272524 150214 272576 150220
rect 272536 149802 272564 150214
rect 272524 149796 272576 149802
rect 272524 149738 272576 149744
rect 272432 148504 272484 148510
rect 272432 148446 272484 148452
rect 272062 142352 272118 142361
rect 272062 142287 272118 142296
rect 272720 137902 272748 235962
rect 272904 233850 272932 316542
rect 272984 316192 273036 316198
rect 272984 316134 273036 316140
rect 272996 236745 273024 316134
rect 273088 295322 273116 372642
rect 273180 296070 273208 374546
rect 273536 320408 273588 320414
rect 273536 320350 273588 320356
rect 273168 296064 273220 296070
rect 273168 296006 273220 296012
rect 273076 295316 273128 295322
rect 273076 295258 273128 295264
rect 273076 249076 273128 249082
rect 273076 249018 273128 249024
rect 273088 240242 273116 249018
rect 273352 243636 273404 243642
rect 273352 243578 273404 243584
rect 273364 241534 273392 243578
rect 273352 241528 273404 241534
rect 273352 241470 273404 241476
rect 273260 241324 273312 241330
rect 273260 241266 273312 241272
rect 273076 240236 273128 240242
rect 273076 240178 273128 240184
rect 273272 239494 273300 241266
rect 273260 239488 273312 239494
rect 273260 239430 273312 239436
rect 272982 236736 273038 236745
rect 272982 236671 273038 236680
rect 272892 233844 272944 233850
rect 272892 233786 272944 233792
rect 273272 143342 273300 239430
rect 273364 152969 273392 241470
rect 273548 233918 273576 320350
rect 273626 315888 273682 315897
rect 273626 315823 273682 315832
rect 273536 233912 273588 233918
rect 273536 233854 273588 233860
rect 273640 228206 273668 315823
rect 273732 313954 273760 393887
rect 273902 387288 273958 387297
rect 273902 387223 273958 387232
rect 273812 371544 273864 371550
rect 273812 371486 273864 371492
rect 273824 321162 273852 371486
rect 273916 321638 273944 387223
rect 273904 321632 273956 321638
rect 273904 321574 273956 321580
rect 273812 321156 273864 321162
rect 273812 321098 273864 321104
rect 273916 320657 273944 321574
rect 273902 320648 273958 320657
rect 273902 320583 273958 320592
rect 274008 319938 274036 393926
rect 274088 392692 274140 392698
rect 274088 392634 274140 392640
rect 273996 319932 274048 319938
rect 273996 319874 274048 319880
rect 273904 316872 273956 316878
rect 273904 316814 273956 316820
rect 273720 313948 273772 313954
rect 273720 313890 273772 313896
rect 273916 241330 273944 316814
rect 273904 241324 273956 241330
rect 273904 241266 273956 241272
rect 273904 235408 273956 235414
rect 273904 235350 273956 235356
rect 273628 228200 273680 228206
rect 273628 228142 273680 228148
rect 273812 153196 273864 153202
rect 273812 153138 273864 153144
rect 273350 152960 273406 152969
rect 273350 152895 273406 152904
rect 273824 152522 273852 153138
rect 273812 152516 273864 152522
rect 273812 152458 273864 152464
rect 273260 143336 273312 143342
rect 273260 143278 273312 143284
rect 273272 142934 273300 143278
rect 273260 142928 273312 142934
rect 273260 142870 273312 142876
rect 272708 137896 272760 137902
rect 272708 137838 272760 137844
rect 272720 137290 272748 137838
rect 272708 137284 272760 137290
rect 272708 137226 272760 137232
rect 272246 136640 272302 136649
rect 272246 136575 272248 136584
rect 272300 136575 272302 136584
rect 272248 136546 272300 136552
rect 272260 135318 272288 136546
rect 272248 135312 272300 135318
rect 272248 135254 272300 135260
rect 273916 126954 273944 235350
rect 274008 229702 274036 319874
rect 274100 314401 274128 392634
rect 274192 319530 274220 397015
rect 274284 345014 274312 400182
rect 274456 397724 274508 397730
rect 274456 397666 274508 397672
rect 274284 344986 274404 345014
rect 274376 320686 274404 344986
rect 274364 320680 274416 320686
rect 274364 320622 274416 320628
rect 274180 319524 274232 319530
rect 274180 319466 274232 319472
rect 274272 318912 274324 318918
rect 274272 318854 274324 318860
rect 274086 314392 274142 314401
rect 274086 314327 274142 314336
rect 274284 232830 274312 318854
rect 274376 233782 274404 320622
rect 274468 317121 274496 397666
rect 274560 374338 274588 465054
rect 280066 454064 280122 454073
rect 280066 453999 280122 454008
rect 278596 452192 278648 452198
rect 278596 452134 278648 452140
rect 278318 448624 278374 448633
rect 277768 448588 277820 448594
rect 278318 448559 278374 448568
rect 277768 448530 277820 448536
rect 277124 400376 277176 400382
rect 277124 400318 277176 400324
rect 275928 399356 275980 399362
rect 275928 399298 275980 399304
rect 275560 395480 275612 395486
rect 275560 395422 275612 395428
rect 275468 387252 275520 387258
rect 275468 387194 275520 387200
rect 275376 387116 275428 387122
rect 275376 387058 275428 387064
rect 274548 374332 274600 374338
rect 274548 374274 274600 374280
rect 274560 363662 274588 374274
rect 275192 372972 275244 372978
rect 275192 372914 275244 372920
rect 274548 363656 274600 363662
rect 274548 363598 274600 363604
rect 275098 320784 275154 320793
rect 275098 320719 275154 320728
rect 274454 317112 274510 317121
rect 274454 317047 274510 317056
rect 274364 233776 274416 233782
rect 274364 233718 274416 233724
rect 274272 232824 274324 232830
rect 274468 232801 274496 317047
rect 274548 314628 274600 314634
rect 274548 314570 274600 314576
rect 274560 313954 274588 314570
rect 274548 313948 274600 313954
rect 274548 313890 274600 313896
rect 274548 309188 274600 309194
rect 274548 309130 274600 309136
rect 274560 242049 274588 309130
rect 275112 248414 275140 320719
rect 275204 294710 275232 372914
rect 275284 371884 275336 371890
rect 275284 371826 275336 371832
rect 275296 324970 275324 371826
rect 275284 324964 275336 324970
rect 275284 324906 275336 324912
rect 275284 321428 275336 321434
rect 275284 321370 275336 321376
rect 275192 294704 275244 294710
rect 275192 294646 275244 294652
rect 274836 248386 275140 248414
rect 274546 242040 274602 242049
rect 274546 241975 274602 241984
rect 274548 241936 274600 241942
rect 274546 241904 274548 241913
rect 274600 241904 274602 241913
rect 274546 241839 274602 241848
rect 274272 232766 274324 232772
rect 274454 232792 274510 232801
rect 274454 232727 274510 232736
rect 273996 229696 274048 229702
rect 273996 229638 274048 229644
rect 274560 152522 274588 241839
rect 274640 241596 274692 241602
rect 274640 241538 274692 241544
rect 274652 237318 274680 241538
rect 274640 237312 274692 237318
rect 274640 237254 274692 237260
rect 274548 152516 274600 152522
rect 274548 152458 274600 152464
rect 274652 148889 274680 237254
rect 274836 233646 274864 248386
rect 274916 243568 274968 243574
rect 274916 243510 274968 243516
rect 274928 239193 274956 243510
rect 274914 239184 274970 239193
rect 274914 239119 274970 239128
rect 274824 233640 274876 233646
rect 274824 233582 274876 233588
rect 274732 229764 274784 229770
rect 274732 229706 274784 229712
rect 274744 229634 274772 229706
rect 274732 229628 274784 229634
rect 274732 229570 274784 229576
rect 274638 148880 274694 148889
rect 274638 148815 274694 148824
rect 274744 146962 274772 229570
rect 274836 149598 274864 233582
rect 274928 157185 274956 239119
rect 275296 232762 275324 321370
rect 275388 320793 275416 387058
rect 275374 320784 275430 320793
rect 275374 320719 275430 320728
rect 275480 319054 275508 387194
rect 275468 319048 275520 319054
rect 275468 318990 275520 318996
rect 275572 317762 275600 395422
rect 275744 395344 275796 395350
rect 275744 395286 275796 395292
rect 275652 374740 275704 374746
rect 275652 374682 275704 374688
rect 275560 317756 275612 317762
rect 275560 317698 275612 317704
rect 275376 316940 275428 316946
rect 275376 316882 275428 316888
rect 275284 232756 275336 232762
rect 275284 232698 275336 232704
rect 275388 229770 275416 316882
rect 275560 315512 275612 315518
rect 275560 315454 275612 315460
rect 275572 240009 275600 315454
rect 275664 292534 275692 374682
rect 275756 316674 275784 395286
rect 275836 373040 275888 373046
rect 275836 372982 275888 372988
rect 275744 316668 275796 316674
rect 275744 316610 275796 316616
rect 275744 313404 275796 313410
rect 275744 313346 275796 313352
rect 275652 292528 275704 292534
rect 275652 292470 275704 292476
rect 275652 253224 275704 253230
rect 275652 253166 275704 253172
rect 275664 241602 275692 253166
rect 275652 241596 275704 241602
rect 275652 241538 275704 241544
rect 275558 240000 275614 240009
rect 275558 239935 275614 239944
rect 275756 237930 275784 313346
rect 275848 293418 275876 372982
rect 275940 314673 275968 399298
rect 277032 397656 277084 397662
rect 277032 397598 277084 397604
rect 276940 396976 276992 396982
rect 276940 396918 276992 396924
rect 276756 394256 276808 394262
rect 276756 394198 276808 394204
rect 276296 392828 276348 392834
rect 276296 392770 276348 392776
rect 276018 368656 276074 368665
rect 276018 368591 276074 368600
rect 276032 368558 276060 368591
rect 276020 368552 276072 368558
rect 276020 368494 276072 368500
rect 276020 354000 276072 354006
rect 276020 353942 276072 353948
rect 276032 353326 276060 353942
rect 276020 353320 276072 353326
rect 276020 353262 276072 353268
rect 276308 316606 276336 392770
rect 276664 388612 276716 388618
rect 276664 388554 276716 388560
rect 276572 371476 276624 371482
rect 276572 371418 276624 371424
rect 276478 368656 276534 368665
rect 276478 368591 276534 368600
rect 276388 316668 276440 316674
rect 276388 316610 276440 316616
rect 276296 316600 276348 316606
rect 276296 316542 276348 316548
rect 275926 314664 275982 314673
rect 275926 314599 275982 314608
rect 275940 314566 275968 314599
rect 275928 314560 275980 314566
rect 275928 314502 275980 314508
rect 275928 309256 275980 309262
rect 275928 309198 275980 309204
rect 275836 293412 275888 293418
rect 275836 293354 275888 293360
rect 275940 241942 275968 309198
rect 276112 242208 276164 242214
rect 276112 242150 276164 242156
rect 275928 241936 275980 241942
rect 275928 241878 275980 241884
rect 276020 240168 276072 240174
rect 276020 240110 276072 240116
rect 275744 237924 275796 237930
rect 275744 237866 275796 237872
rect 276032 236842 276060 240110
rect 276020 236836 276072 236842
rect 276020 236778 276072 236784
rect 275376 229764 275428 229770
rect 275376 229706 275428 229712
rect 275928 229764 275980 229770
rect 275928 229706 275980 229712
rect 274914 157176 274970 157185
rect 274914 157111 274970 157120
rect 275940 156534 275968 229706
rect 275928 156528 275980 156534
rect 275928 156470 275980 156476
rect 276124 154465 276152 242150
rect 276296 237312 276348 237318
rect 276296 237254 276348 237260
rect 276308 236570 276336 237254
rect 276296 236564 276348 236570
rect 276296 236506 276348 236512
rect 276204 233232 276256 233238
rect 276204 233174 276256 233180
rect 276216 231062 276244 233174
rect 276204 231056 276256 231062
rect 276204 230998 276256 231004
rect 276110 154456 276166 154465
rect 276110 154391 276166 154400
rect 274824 149592 274876 149598
rect 274824 149534 274876 149540
rect 274836 149122 274864 149534
rect 274824 149116 274876 149122
rect 274824 149058 274876 149064
rect 275284 149116 275336 149122
rect 275284 149058 275336 149064
rect 274652 146934 274772 146962
rect 274652 144770 274680 146934
rect 274640 144764 274692 144770
rect 274640 144706 274692 144712
rect 274652 144362 274680 144706
rect 274640 144356 274692 144362
rect 274640 144298 274692 144304
rect 273904 126948 273956 126954
rect 273904 126890 273956 126896
rect 274088 126948 274140 126954
rect 274088 126890 274140 126896
rect 274100 126274 274128 126890
rect 274088 126268 274140 126274
rect 274088 126210 274140 126216
rect 271892 16546 272472 16574
rect 271236 3868 271288 3874
rect 271236 3810 271288 3816
rect 271144 3392 271196 3398
rect 271144 3334 271196 3340
rect 271248 480 271276 3810
rect 272444 480 272472 16546
rect 275296 4146 275324 149058
rect 276216 146742 276244 230998
rect 276308 153105 276336 236506
rect 276400 221610 276428 316610
rect 276388 221604 276440 221610
rect 276388 221546 276440 221552
rect 276492 153202 276520 368591
rect 276584 326398 276612 371418
rect 276572 326392 276624 326398
rect 276572 326334 276624 326340
rect 276676 322153 276704 388554
rect 276662 322144 276718 322153
rect 276662 322079 276718 322088
rect 276768 321065 276796 394198
rect 276754 321056 276810 321065
rect 276754 320991 276810 321000
rect 276664 318844 276716 318850
rect 276664 318786 276716 318792
rect 276676 229906 276704 318786
rect 276768 315353 276796 320991
rect 276952 319870 276980 396918
rect 276940 319864 276992 319870
rect 276940 319806 276992 319812
rect 276952 319462 276980 319806
rect 276940 319456 276992 319462
rect 276940 319398 276992 319404
rect 277044 318034 277072 397598
rect 277136 319598 277164 400318
rect 277216 399424 277268 399430
rect 277216 399366 277268 399372
rect 277124 319592 277176 319598
rect 277124 319534 277176 319540
rect 277228 318510 277256 399366
rect 277308 374060 277360 374066
rect 277308 374002 277360 374008
rect 277320 353326 277348 374002
rect 277780 371793 277808 448530
rect 278042 390280 278098 390289
rect 278042 390215 278098 390224
rect 277860 386028 277912 386034
rect 277860 385970 277912 385976
rect 277766 371784 277822 371793
rect 277766 371719 277822 371728
rect 277308 353320 277360 353326
rect 277308 353262 277360 353268
rect 277872 321026 277900 385970
rect 277952 373516 278004 373522
rect 277952 373458 278004 373464
rect 277860 321020 277912 321026
rect 277860 320962 277912 320968
rect 277858 320920 277914 320929
rect 277858 320855 277914 320864
rect 277872 320249 277900 320855
rect 277858 320240 277914 320249
rect 277858 320175 277914 320184
rect 277306 318880 277362 318889
rect 277306 318815 277362 318824
rect 277216 318504 277268 318510
rect 277216 318446 277268 318452
rect 277032 318028 277084 318034
rect 277032 317970 277084 317976
rect 276848 317484 276900 317490
rect 276848 317426 276900 317432
rect 276754 315344 276810 315353
rect 276754 315279 276810 315288
rect 276860 234054 276888 317426
rect 277044 317234 277072 317970
rect 277228 317490 277256 318446
rect 277216 317484 277268 317490
rect 277216 317426 277268 317432
rect 276952 317206 277072 317234
rect 276952 235890 276980 317206
rect 277032 317076 277084 317082
rect 277032 317018 277084 317024
rect 277044 237114 277072 317018
rect 277122 245168 277178 245177
rect 277122 245103 277178 245112
rect 277136 237318 277164 245103
rect 277124 237312 277176 237318
rect 277124 237254 277176 237260
rect 277032 237108 277084 237114
rect 277032 237050 277084 237056
rect 276940 235884 276992 235890
rect 276940 235826 276992 235832
rect 276848 234048 276900 234054
rect 276848 233990 276900 233996
rect 276664 229900 276716 229906
rect 276664 229842 276716 229848
rect 277044 229770 277072 237050
rect 277320 231441 277348 318815
rect 277768 317008 277820 317014
rect 277768 316950 277820 316956
rect 277492 242276 277544 242282
rect 277492 242218 277544 242224
rect 277400 237312 277452 237318
rect 277400 237254 277452 237260
rect 277412 236502 277440 237254
rect 277400 236496 277452 236502
rect 277400 236438 277452 236444
rect 277306 231432 277362 231441
rect 277306 231367 277362 231376
rect 277032 229764 277084 229770
rect 277032 229706 277084 229712
rect 277412 229158 277440 236438
rect 277400 229152 277452 229158
rect 277400 229094 277452 229100
rect 277504 160721 277532 242218
rect 277780 234122 277808 316950
rect 277860 312384 277912 312390
rect 277860 312326 277912 312332
rect 277872 235754 277900 312326
rect 277964 294642 277992 373458
rect 278056 361729 278084 390215
rect 278228 385688 278280 385694
rect 278228 385630 278280 385636
rect 278136 373108 278188 373114
rect 278136 373050 278188 373056
rect 278042 361720 278098 361729
rect 278042 361655 278098 361664
rect 278044 353320 278096 353326
rect 278044 353262 278096 353268
rect 277952 294636 278004 294642
rect 277952 294578 278004 294584
rect 277860 235748 277912 235754
rect 277860 235690 277912 235696
rect 277768 234116 277820 234122
rect 277768 234058 277820 234064
rect 278056 233306 278084 353262
rect 278148 293282 278176 373050
rect 278240 321554 278268 385630
rect 278332 373425 278360 448559
rect 278412 395548 278464 395554
rect 278412 395490 278464 395496
rect 278318 373416 278374 373425
rect 278318 373351 278320 373360
rect 278372 373351 278374 373360
rect 278320 373322 278372 373328
rect 278332 373291 278360 373322
rect 278318 371784 278374 371793
rect 278318 371719 278374 371728
rect 278332 370530 278360 371719
rect 278320 370524 278372 370530
rect 278320 370466 278372 370472
rect 278240 321526 278360 321554
rect 278226 320648 278282 320657
rect 278226 320583 278282 320592
rect 278240 320249 278268 320583
rect 278226 320240 278282 320249
rect 278226 320175 278282 320184
rect 278332 319569 278360 321526
rect 278318 319560 278374 319569
rect 278318 319495 278374 319504
rect 278332 318889 278360 319495
rect 278424 319025 278452 395490
rect 278504 374060 278556 374066
rect 278504 374002 278556 374008
rect 278516 319326 278544 374002
rect 278608 373318 278636 452134
rect 279884 450220 279936 450226
rect 279884 450162 279936 450168
rect 278688 399016 278740 399022
rect 278688 398958 278740 398964
rect 278596 373312 278648 373318
rect 278596 373254 278648 373260
rect 278596 373176 278648 373182
rect 278596 373118 278648 373124
rect 278504 319320 278556 319326
rect 278504 319262 278556 319268
rect 278410 319016 278466 319025
rect 278410 318951 278466 318960
rect 278318 318880 278374 318889
rect 278318 318815 278374 318824
rect 278318 317520 278374 317529
rect 278318 317455 278374 317464
rect 278228 315716 278280 315722
rect 278228 315658 278280 315664
rect 278136 293276 278188 293282
rect 278136 293218 278188 293224
rect 278136 240576 278188 240582
rect 278136 240518 278188 240524
rect 278148 239698 278176 240518
rect 278136 239692 278188 239698
rect 278136 239634 278188 239640
rect 278136 239488 278188 239494
rect 278136 239430 278188 239436
rect 278148 238814 278176 239430
rect 278136 238808 278188 238814
rect 278136 238750 278188 238756
rect 278044 233300 278096 233306
rect 278044 233242 278096 233248
rect 277860 232824 277912 232830
rect 277860 232766 277912 232772
rect 277872 231402 277900 232766
rect 277584 231396 277636 231402
rect 277584 231338 277636 231344
rect 277860 231396 277912 231402
rect 277860 231338 277912 231344
rect 277490 160712 277546 160721
rect 277490 160647 277546 160656
rect 276480 153196 276532 153202
rect 276480 153138 276532 153144
rect 276294 153096 276350 153105
rect 276294 153031 276350 153040
rect 276204 146736 276256 146742
rect 276204 146678 276256 146684
rect 277596 143478 277624 231338
rect 278044 148368 278096 148374
rect 278044 148310 278096 148316
rect 277584 143472 277636 143478
rect 277584 143414 277636 143420
rect 275284 4140 275336 4146
rect 275284 4082 275336 4088
rect 276020 3664 276072 3670
rect 276020 3606 276072 3612
rect 273626 3496 273682 3505
rect 273626 3431 273682 3440
rect 273640 480 273668 3431
rect 274824 3392 274876 3398
rect 274824 3334 274876 3340
rect 274836 480 274864 3334
rect 276032 480 276060 3606
rect 278056 3398 278084 148310
rect 278148 144838 278176 238750
rect 278240 227322 278268 315658
rect 278332 233238 278360 317455
rect 278424 312594 278452 318951
rect 278516 318850 278544 319262
rect 278504 318844 278556 318850
rect 278504 318786 278556 318792
rect 278504 316396 278556 316402
rect 278504 316338 278556 316344
rect 278412 312588 278464 312594
rect 278412 312530 278464 312536
rect 278412 239760 278464 239766
rect 278412 239702 278464 239708
rect 278424 239630 278452 239702
rect 278412 239624 278464 239630
rect 278412 239566 278464 239572
rect 278516 237318 278544 316338
rect 278608 293350 278636 373118
rect 278700 317286 278728 398958
rect 279700 394188 279752 394194
rect 279700 394130 279752 394136
rect 279148 386436 279200 386442
rect 279148 386378 279200 386384
rect 278780 373448 278832 373454
rect 278780 373390 278832 373396
rect 278792 373182 278820 373390
rect 278780 373176 278832 373182
rect 278780 373118 278832 373124
rect 279160 369238 279188 386378
rect 279516 385892 279568 385898
rect 279516 385834 279568 385840
rect 279424 381200 279476 381206
rect 279424 381142 279476 381148
rect 279240 372428 279292 372434
rect 279240 372370 279292 372376
rect 279148 369232 279200 369238
rect 279148 369174 279200 369180
rect 279252 349858 279280 372370
rect 279332 369980 279384 369986
rect 279332 369922 279384 369928
rect 279240 349852 279292 349858
rect 279240 349794 279292 349800
rect 279238 321872 279294 321881
rect 279238 321807 279294 321816
rect 279252 321609 279280 321807
rect 279238 321600 279294 321609
rect 279238 321535 279294 321544
rect 278688 317280 278740 317286
rect 278688 317222 278740 317228
rect 278700 317014 278728 317222
rect 278688 317008 278740 317014
rect 278688 316950 278740 316956
rect 279240 317008 279292 317014
rect 279240 316950 279292 316956
rect 278688 312588 278740 312594
rect 278688 312530 278740 312536
rect 278596 293344 278648 293350
rect 278596 293286 278648 293292
rect 278504 237312 278556 237318
rect 278504 237254 278556 237260
rect 278700 234025 278728 312530
rect 278778 243808 278834 243817
rect 278778 243743 278834 243752
rect 278792 243001 278820 243743
rect 278778 242992 278834 243001
rect 278834 242950 278912 242978
rect 278778 242927 278834 242936
rect 278780 236768 278832 236774
rect 278780 236710 278832 236716
rect 278792 235890 278820 236710
rect 278780 235884 278832 235890
rect 278780 235826 278832 235832
rect 278686 234016 278742 234025
rect 278686 233951 278742 233960
rect 278320 233232 278372 233238
rect 278320 233174 278372 233180
rect 278412 232620 278464 232626
rect 278412 232562 278464 232568
rect 278228 227316 278280 227322
rect 278228 227258 278280 227264
rect 278424 148170 278452 232562
rect 278412 148164 278464 148170
rect 278412 148106 278464 148112
rect 278136 144832 278188 144838
rect 278136 144774 278188 144780
rect 278688 143472 278740 143478
rect 278688 143414 278740 143420
rect 278700 143002 278728 143414
rect 278688 142996 278740 143002
rect 278688 142938 278740 142944
rect 278792 16574 278820 235826
rect 278884 144809 278912 242950
rect 279252 232626 279280 316950
rect 279344 291922 279372 369922
rect 279436 358086 279464 381142
rect 279424 358080 279476 358086
rect 279424 358022 279476 358028
rect 279528 321434 279556 385834
rect 279608 385756 279660 385762
rect 279608 385698 279660 385704
rect 279516 321428 279568 321434
rect 279516 321370 279568 321376
rect 279514 321328 279570 321337
rect 279514 321263 279570 321272
rect 279424 313472 279476 313478
rect 279424 313414 279476 313420
rect 279332 291916 279384 291922
rect 279332 291858 279384 291864
rect 279240 232620 279292 232626
rect 279240 232562 279292 232568
rect 278964 231192 279016 231198
rect 278964 231134 279016 231140
rect 278976 147490 279004 231134
rect 279436 220658 279464 313414
rect 279528 231198 279556 321263
rect 279620 318617 279648 385698
rect 279712 318889 279740 394130
rect 279792 392896 279844 392902
rect 279792 392838 279844 392844
rect 279698 318880 279754 318889
rect 279698 318815 279754 318824
rect 279606 318608 279662 318617
rect 279606 318543 279662 318552
rect 279620 317529 279648 318543
rect 279606 317520 279662 317529
rect 279606 317455 279662 317464
rect 279608 317212 279660 317218
rect 279608 317154 279660 317160
rect 279516 231192 279568 231198
rect 279516 231134 279568 231140
rect 279620 229838 279648 317154
rect 279712 233986 279740 318815
rect 279804 313614 279832 392838
rect 279896 371006 279924 450162
rect 279976 400512 280028 400518
rect 279976 400454 280028 400460
rect 279884 371000 279936 371006
rect 279884 370942 279936 370948
rect 279896 369986 279924 370942
rect 279884 369980 279936 369986
rect 279884 369922 279936 369928
rect 279882 361856 279938 361865
rect 279882 361791 279938 361800
rect 279896 361622 279924 361791
rect 279884 361616 279936 361622
rect 279884 361558 279936 361564
rect 279988 319666 280016 400454
rect 280080 371929 280108 453999
rect 280618 452024 280674 452033
rect 280618 451959 280674 451968
rect 280632 372065 280660 451959
rect 280712 385960 280764 385966
rect 280712 385902 280764 385908
rect 280618 372056 280674 372065
rect 280618 371991 280674 372000
rect 280632 371958 280660 371991
rect 280620 371952 280672 371958
rect 280066 371920 280122 371929
rect 280620 371894 280672 371900
rect 280066 371855 280122 371864
rect 280080 370666 280108 371855
rect 280620 371748 280672 371754
rect 280620 371690 280672 371696
rect 280528 371680 280580 371686
rect 280528 371622 280580 371628
rect 280068 370660 280120 370666
rect 280068 370602 280120 370608
rect 280540 362234 280568 371622
rect 280528 362228 280580 362234
rect 280528 362170 280580 362176
rect 280068 361616 280120 361622
rect 280068 361558 280120 361564
rect 279976 319660 280028 319666
rect 279976 319602 280028 319608
rect 279884 317552 279936 317558
rect 279884 317494 279936 317500
rect 279792 313608 279844 313614
rect 279792 313550 279844 313556
rect 279896 234394 279924 317494
rect 279884 234388 279936 234394
rect 279884 234330 279936 234336
rect 279700 233980 279752 233986
rect 279700 233922 279752 233928
rect 279608 229832 279660 229838
rect 279608 229774 279660 229780
rect 279424 220652 279476 220658
rect 279424 220594 279476 220600
rect 278964 147484 279016 147490
rect 278964 147426 279016 147432
rect 279976 147484 280028 147490
rect 279976 147426 280028 147432
rect 279988 146946 280016 147426
rect 279976 146940 280028 146946
rect 279976 146882 280028 146888
rect 278870 144800 278926 144809
rect 278870 144735 278926 144744
rect 280080 33114 280108 361558
rect 280632 359514 280660 371690
rect 280620 359508 280672 359514
rect 280620 359450 280672 359456
rect 280158 320784 280214 320793
rect 280158 320719 280214 320728
rect 280172 316810 280200 320719
rect 280620 320680 280672 320686
rect 280620 320622 280672 320628
rect 280528 319660 280580 319666
rect 280528 319602 280580 319608
rect 280540 318918 280568 319602
rect 280528 318912 280580 318918
rect 280528 318854 280580 318860
rect 280632 317490 280660 320622
rect 280724 320550 280752 385902
rect 280816 373969 280844 700266
rect 298744 670744 298796 670750
rect 298744 670686 298796 670692
rect 281448 464364 281500 464370
rect 281448 464306 281500 464312
rect 281460 463758 281488 464306
rect 281448 463752 281500 463758
rect 281448 463694 281500 463700
rect 281356 454980 281408 454986
rect 281356 454922 281408 454928
rect 280894 451616 280950 451625
rect 280894 451551 280950 451560
rect 280802 373960 280858 373969
rect 280802 373895 280858 373904
rect 280816 373017 280844 373895
rect 280908 373289 280936 451551
rect 281264 400580 281316 400586
rect 281264 400522 281316 400528
rect 281080 400308 281132 400314
rect 281080 400250 281132 400256
rect 280988 396908 281040 396914
rect 280988 396850 281040 396856
rect 280894 373280 280950 373289
rect 280894 373215 280950 373224
rect 280802 373008 280858 373017
rect 280802 372943 280858 372952
rect 280896 371612 280948 371618
rect 280896 371554 280948 371560
rect 280804 370048 280856 370054
rect 280804 369990 280856 369996
rect 280816 345710 280844 369990
rect 280908 351218 280936 371554
rect 280896 351212 280948 351218
rect 280896 351154 280948 351160
rect 280804 345704 280856 345710
rect 280804 345646 280856 345652
rect 281000 326602 281028 396850
rect 280988 326596 281040 326602
rect 280988 326538 281040 326544
rect 281092 326482 281120 400250
rect 281172 375352 281224 375358
rect 281172 375294 281224 375300
rect 281184 374814 281212 375294
rect 281172 374808 281224 374814
rect 281172 374750 281224 374756
rect 280816 326454 281120 326482
rect 280712 320544 280764 320550
rect 280712 320486 280764 320492
rect 280816 320226 280844 326454
rect 280988 326392 281040 326398
rect 281040 326340 281120 326346
rect 280988 326334 281120 326340
rect 281000 326318 281120 326334
rect 280988 322992 281040 322998
rect 280988 322934 281040 322940
rect 280896 320884 280948 320890
rect 280896 320826 280948 320832
rect 280724 320198 280844 320226
rect 280724 318850 280752 320198
rect 280908 319734 280936 320826
rect 280896 319728 280948 319734
rect 280896 319670 280948 319676
rect 280896 318912 280948 318918
rect 280896 318854 280948 318860
rect 280712 318844 280764 318850
rect 280712 318786 280764 318792
rect 280620 317484 280672 317490
rect 280620 317426 280672 317432
rect 280160 316804 280212 316810
rect 280160 316746 280212 316752
rect 280724 311894 280752 318786
rect 280804 318572 280856 318578
rect 280804 318514 280856 318520
rect 280632 311866 280752 311894
rect 280252 232484 280304 232490
rect 280252 232426 280304 232432
rect 280160 231124 280212 231130
rect 280160 231066 280212 231072
rect 280172 151774 280200 231066
rect 280264 229566 280292 232426
rect 280632 232354 280660 311866
rect 280712 307420 280764 307426
rect 280712 307362 280764 307368
rect 280724 239358 280752 307362
rect 280712 239352 280764 239358
rect 280712 239294 280764 239300
rect 280620 232348 280672 232354
rect 280620 232290 280672 232296
rect 280252 229560 280304 229566
rect 280252 229502 280304 229508
rect 280264 153134 280292 229502
rect 280816 223038 280844 318514
rect 280908 227118 280936 318854
rect 281000 318714 281028 322934
rect 280988 318708 281040 318714
rect 280988 318650 281040 318656
rect 281092 317422 281120 326318
rect 281080 317416 281132 317422
rect 281080 317358 281132 317364
rect 281078 316160 281134 316169
rect 281078 316095 281134 316104
rect 281092 232830 281120 316095
rect 281184 292466 281212 374750
rect 281276 317966 281304 400522
rect 281368 371210 281396 454922
rect 281460 375358 281488 463694
rect 298756 456822 298784 670686
rect 298744 456816 298796 456822
rect 298744 456758 298796 456764
rect 299388 456816 299440 456822
rect 299388 456758 299440 456764
rect 294696 454844 294748 454850
rect 294696 454786 294748 454792
rect 293868 454436 293920 454442
rect 293868 454378 293920 454384
rect 282826 451752 282882 451761
rect 282826 451687 282882 451696
rect 282182 448760 282238 448769
rect 282182 448695 282238 448704
rect 281632 395684 281684 395690
rect 281632 395626 281684 395632
rect 281540 395616 281592 395622
rect 281540 395558 281592 395564
rect 281448 375352 281500 375358
rect 281448 375294 281500 375300
rect 281448 373516 281500 373522
rect 281448 373458 281500 373464
rect 281460 373114 281488 373458
rect 281448 373108 281500 373114
rect 281448 373050 281500 373056
rect 281356 371204 281408 371210
rect 281356 371146 281408 371152
rect 281368 370734 281396 371146
rect 281356 370728 281408 370734
rect 281356 370670 281408 370676
rect 281448 370252 281500 370258
rect 281448 370194 281500 370200
rect 281356 320544 281408 320550
rect 281356 320486 281408 320492
rect 281368 318238 281396 320486
rect 281356 318232 281408 318238
rect 281356 318174 281408 318180
rect 281264 317960 281316 317966
rect 281264 317902 281316 317908
rect 281356 315648 281408 315654
rect 281356 315590 281408 315596
rect 281264 315580 281316 315586
rect 281264 315522 281316 315528
rect 281172 292460 281224 292466
rect 281172 292402 281224 292408
rect 281170 245304 281226 245313
rect 281170 245239 281226 245248
rect 281080 232824 281132 232830
rect 281080 232766 281132 232772
rect 280896 227112 280948 227118
rect 280896 227054 280948 227060
rect 280804 223032 280856 223038
rect 280804 222974 280856 222980
rect 281184 220590 281212 245239
rect 281276 235618 281304 315522
rect 281368 237386 281396 315590
rect 281460 291650 281488 370194
rect 281552 318306 281580 395558
rect 281644 319977 281672 395626
rect 281724 391400 281776 391406
rect 281724 391342 281776 391348
rect 281630 319968 281686 319977
rect 281630 319903 281686 319912
rect 281540 318300 281592 318306
rect 281540 318242 281592 318248
rect 281644 318170 281672 319903
rect 281736 319802 281764 391342
rect 281816 389972 281868 389978
rect 281816 389914 281868 389920
rect 281724 319796 281776 319802
rect 281724 319738 281776 319744
rect 281828 319705 281856 389914
rect 282000 374672 282052 374678
rect 282000 374614 282052 374620
rect 282012 372026 282040 374614
rect 282196 373250 282224 448695
rect 282368 392964 282420 392970
rect 282368 392906 282420 392912
rect 282276 373992 282328 373998
rect 282276 373934 282328 373940
rect 282184 373244 282236 373250
rect 282184 373186 282236 373192
rect 282000 372020 282052 372026
rect 282000 371962 282052 371968
rect 282012 363633 282040 371962
rect 282288 371822 282316 373934
rect 282276 371816 282328 371822
rect 282276 371758 282328 371764
rect 282276 370388 282328 370394
rect 282276 370330 282328 370336
rect 281998 363624 282054 363633
rect 281998 363559 282054 363568
rect 282182 361720 282238 361729
rect 282182 361655 282238 361664
rect 282090 322960 282146 322969
rect 282090 322895 282146 322904
rect 281906 322144 281962 322153
rect 281906 322079 281962 322088
rect 281920 320006 281948 322079
rect 281998 321736 282054 321745
rect 281998 321671 282054 321680
rect 282012 321434 282040 321671
rect 282000 321428 282052 321434
rect 282000 321370 282052 321376
rect 281998 321192 282054 321201
rect 281998 321127 282054 321136
rect 282012 320657 282040 321127
rect 282104 320754 282132 322895
rect 282092 320748 282144 320754
rect 282092 320690 282144 320696
rect 281998 320648 282054 320657
rect 282196 320634 282224 361655
rect 281998 320583 282054 320592
rect 282104 320606 282224 320634
rect 282000 320068 282052 320074
rect 282000 320010 282052 320016
rect 281908 320000 281960 320006
rect 281908 319942 281960 319948
rect 281814 319696 281870 319705
rect 281814 319631 281870 319640
rect 282012 319462 282040 320010
rect 282104 319954 282132 320606
rect 282184 320340 282236 320346
rect 282184 320282 282236 320288
rect 282196 320142 282224 320282
rect 282184 320136 282236 320142
rect 282184 320078 282236 320084
rect 282104 319926 282224 319954
rect 282000 319456 282052 319462
rect 282000 319398 282052 319404
rect 282196 318238 282224 319926
rect 282184 318232 282236 318238
rect 282184 318174 282236 318180
rect 281632 318164 281684 318170
rect 281632 318106 281684 318112
rect 281908 307488 281960 307494
rect 281908 307430 281960 307436
rect 281448 291644 281500 291650
rect 281448 291586 281500 291592
rect 281538 240272 281594 240281
rect 281538 240207 281594 240216
rect 281552 237454 281580 240207
rect 281540 237448 281592 237454
rect 281540 237390 281592 237396
rect 281356 237380 281408 237386
rect 281356 237322 281408 237328
rect 281264 235612 281316 235618
rect 281264 235554 281316 235560
rect 281920 234190 281948 307430
rect 282092 297220 282144 297226
rect 282092 297162 282144 297168
rect 282000 247716 282052 247722
rect 282000 247658 282052 247664
rect 281908 234184 281960 234190
rect 281908 234126 281960 234132
rect 282012 226846 282040 247658
rect 282104 239290 282132 297162
rect 282092 239284 282144 239290
rect 282092 239226 282144 239232
rect 282000 226840 282052 226846
rect 282000 226782 282052 226788
rect 282012 226370 282040 226782
rect 281540 226364 281592 226370
rect 281540 226306 281592 226312
rect 282000 226364 282052 226370
rect 282000 226306 282052 226312
rect 281172 220584 281224 220590
rect 281172 220526 281224 220532
rect 281184 219434 281212 220526
rect 280816 219406 281212 219434
rect 280816 160138 280844 219406
rect 280804 160132 280856 160138
rect 280804 160074 280856 160080
rect 280816 158778 280844 160074
rect 280804 158772 280856 158778
rect 280804 158714 280856 158720
rect 280252 153128 280304 153134
rect 280252 153070 280304 153076
rect 281448 153128 281500 153134
rect 281448 153070 281500 153076
rect 281460 152658 281488 153070
rect 281448 152652 281500 152658
rect 281448 152594 281500 152600
rect 280160 151768 280212 151774
rect 280160 151710 280212 151716
rect 280172 150482 280200 151710
rect 280160 150476 280212 150482
rect 280160 150418 280212 150424
rect 280804 150476 280856 150482
rect 280804 150418 280856 150424
rect 280816 140078 280844 150418
rect 281552 140758 281580 226306
rect 282196 216306 282224 318174
rect 282288 291990 282316 370330
rect 282380 321609 282408 392906
rect 282460 371816 282512 371822
rect 282460 371758 282512 371764
rect 282472 352617 282500 371758
rect 282840 371385 282868 451687
rect 285954 448896 286010 448905
rect 285954 448831 286010 448840
rect 282920 393304 282972 393310
rect 282920 393246 282972 393252
rect 282932 392057 282960 393246
rect 282918 392048 282974 392057
rect 282918 391983 282974 391992
rect 283564 384328 283616 384334
rect 283564 384270 283616 384276
rect 283576 374066 283604 384270
rect 283564 374060 283616 374066
rect 283564 374002 283616 374008
rect 282826 371376 282882 371385
rect 282826 371311 282882 371320
rect 283576 369866 283604 374002
rect 284114 373960 284170 373969
rect 284114 373895 284170 373904
rect 284128 371657 284156 373895
rect 284206 373280 284262 373289
rect 284206 373215 284262 373224
rect 284114 371648 284170 371657
rect 284114 371583 284170 371592
rect 284220 369866 284248 373215
rect 285220 371952 285272 371958
rect 285220 371894 285272 371900
rect 285080 369880 285136 369889
rect 283576 369838 284004 369866
rect 284220 369838 284372 369866
rect 285232 369866 285260 371894
rect 285968 370025 285996 448831
rect 290462 447944 290518 447953
rect 290462 447879 290518 447888
rect 286322 447808 286378 447817
rect 286322 447743 286378 447752
rect 286336 379514 286364 447743
rect 287704 435396 287756 435402
rect 287704 435338 287756 435344
rect 286416 409148 286468 409154
rect 286416 409090 286468 409096
rect 286060 379486 286364 379514
rect 286060 372745 286088 379486
rect 286046 372736 286102 372745
rect 286046 372671 286102 372680
rect 285954 370016 286010 370025
rect 285954 369951 286010 369960
rect 286060 369866 286088 372671
rect 286428 370161 286456 409090
rect 286784 378888 286836 378894
rect 286784 378830 286836 378836
rect 286508 373244 286560 373250
rect 286508 373186 286560 373192
rect 286414 370152 286470 370161
rect 286520 370138 286548 373186
rect 286520 370110 286594 370138
rect 286414 370087 286470 370096
rect 285232 369838 285476 369866
rect 285844 369838 286088 369866
rect 286566 369852 286594 370110
rect 285080 369815 285136 369824
rect 286184 369744 286240 369753
rect 286184 369679 286240 369688
rect 286796 369481 286824 378830
rect 287716 374513 287744 435338
rect 289728 418804 289780 418810
rect 289728 418746 289780 418752
rect 289084 398404 289136 398410
rect 289084 398346 289136 398352
rect 289096 376825 289124 398346
rect 289082 376816 289138 376825
rect 289082 376751 289138 376760
rect 287150 374504 287206 374513
rect 287150 374439 287206 374448
rect 287702 374504 287758 374513
rect 287702 374439 287758 374448
rect 287164 374105 287192 374439
rect 287150 374096 287206 374105
rect 287150 374031 287206 374040
rect 287058 370016 287114 370025
rect 287058 369951 287114 369960
rect 287072 369753 287100 369951
rect 286920 369744 286976 369753
rect 286920 369679 286976 369688
rect 287058 369744 287114 369753
rect 287058 369679 287114 369688
rect 284482 369472 284538 369481
rect 286782 369472 286838 369481
rect 284538 369430 284740 369458
rect 284482 369407 284538 369416
rect 287164 369458 287192 374031
rect 287428 373380 287480 373386
rect 287428 373322 287480 373328
rect 287440 369866 287468 373322
rect 288532 373312 288584 373318
rect 288532 373254 288584 373260
rect 288256 372088 288308 372094
rect 288256 372030 288308 372036
rect 287794 371920 287850 371929
rect 287794 371855 287850 371864
rect 287808 371278 287836 371855
rect 288268 371521 288296 372030
rect 288254 371512 288310 371521
rect 288254 371447 288310 371456
rect 287796 371272 287848 371278
rect 287796 371214 287848 371220
rect 287440 369838 287684 369866
rect 288268 369854 288296 371447
rect 288544 369866 288572 373254
rect 289740 372201 289768 418746
rect 290476 383654 290504 447879
rect 291842 443592 291898 443601
rect 291842 443527 291898 443536
rect 290200 383626 290504 383654
rect 290200 374134 290228 383626
rect 291856 375834 291884 443527
rect 291936 406496 291988 406502
rect 291936 406438 291988 406444
rect 291844 375828 291896 375834
rect 291844 375770 291896 375776
rect 291948 375426 291976 406438
rect 293880 386442 293908 454378
rect 294604 452124 294656 452130
rect 294604 452066 294656 452072
rect 292580 386436 292632 386442
rect 292580 386378 292632 386384
rect 293868 386436 293920 386442
rect 293868 386378 293920 386384
rect 292592 383654 292620 386378
rect 292592 383626 293356 383654
rect 292304 375828 292356 375834
rect 292304 375770 292356 375776
rect 291752 375420 291804 375426
rect 291752 375362 291804 375368
rect 291936 375420 291988 375426
rect 291936 375362 291988 375368
rect 290188 374128 290240 374134
rect 290188 374070 290240 374076
rect 289726 372192 289782 372201
rect 289726 372127 289782 372136
rect 289740 371385 289768 372127
rect 290002 371784 290058 371793
rect 290002 371719 290058 371728
rect 289726 371376 289782 371385
rect 289726 371311 289782 371320
rect 289740 369866 289768 371311
rect 288268 369826 288434 369854
rect 288544 369838 288788 369866
rect 289524 369838 289768 369866
rect 290016 369594 290044 371719
rect 290200 370138 290228 374070
rect 291764 372366 291792 375362
rect 291752 372360 291804 372366
rect 291752 372302 291804 372308
rect 290464 371884 290516 371890
rect 290464 371826 290516 371832
rect 290476 370530 290504 371826
rect 290740 371272 290792 371278
rect 290740 371214 290792 371220
rect 290464 370524 290516 370530
rect 290464 370466 290516 370472
rect 290200 370110 290274 370138
rect 290246 369852 290274 370110
rect 289892 369566 290044 369594
rect 290476 369594 290504 370466
rect 290752 369866 290780 371214
rect 291764 370138 291792 372302
rect 291844 371272 291896 371278
rect 291844 371214 291896 371220
rect 291718 370110 291792 370138
rect 290752 369838 290996 369866
rect 291120 369838 291608 369866
rect 291718 369852 291746 370110
rect 291856 369866 291884 371214
rect 292316 369866 292344 375770
rect 293224 372632 293276 372638
rect 293224 372574 293276 372580
rect 293040 372224 293092 372230
rect 293040 372166 293092 372172
rect 293052 369986 293080 372166
rect 293236 370138 293264 372574
rect 293190 370110 293264 370138
rect 293040 369980 293092 369986
rect 293040 369922 293092 369928
rect 291856 369838 292100 369866
rect 292316 369838 292468 369866
rect 290476 369566 290628 369594
rect 287288 369472 287344 369481
rect 287164 369430 287288 369458
rect 286782 369407 286838 369416
rect 291120 369442 291148 369838
rect 291580 369782 291608 369838
rect 291568 369776 291620 369782
rect 291568 369718 291620 369724
rect 292316 369442 292344 369838
rect 293052 369730 293080 369922
rect 293190 369852 293218 370110
rect 293328 369866 293356 383626
rect 294420 375760 294472 375766
rect 294420 375702 294472 375708
rect 294328 373516 294380 373522
rect 294328 373458 294380 373464
rect 293868 372156 293920 372162
rect 293868 372098 293920 372104
rect 293880 371414 293908 372098
rect 293868 371408 293920 371414
rect 293868 371350 293920 371356
rect 293880 370138 293908 371350
rect 294340 370138 294368 373458
rect 293880 370110 293954 370138
rect 293328 369838 293572 369866
rect 293926 369852 293954 370110
rect 294294 370110 294368 370138
rect 294294 369852 294322 370110
rect 294432 369866 294460 375702
rect 294616 370530 294644 452066
rect 294708 375766 294736 454786
rect 294788 452940 294840 452946
rect 294788 452882 294840 452888
rect 294696 375760 294748 375766
rect 294696 375702 294748 375708
rect 294800 374542 294828 452882
rect 297456 450832 297508 450838
rect 297456 450774 297508 450780
rect 297364 450288 297416 450294
rect 297364 450230 297416 450236
rect 295340 398472 295392 398478
rect 295340 398414 295392 398420
rect 295352 397225 295380 398414
rect 295338 397216 295394 397225
rect 295338 397151 295394 397160
rect 297376 379514 297404 450230
rect 297100 379486 297404 379514
rect 294788 374536 294840 374542
rect 294788 374478 294840 374484
rect 294800 373522 294828 374478
rect 297100 374406 297128 379486
rect 297468 375698 297496 450774
rect 298744 449200 298796 449206
rect 298744 449142 298796 449148
rect 297546 401296 297602 401305
rect 297546 401231 297602 401240
rect 297456 375692 297508 375698
rect 297456 375634 297508 375640
rect 297468 375426 297496 375634
rect 297560 375494 297588 401231
rect 298756 379514 298784 449142
rect 299400 403646 299428 456758
rect 299492 453422 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364524 700392 364576 700398
rect 364524 700334 364576 700340
rect 304264 700324 304316 700330
rect 304264 700266 304316 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 364432 700324 364484 700330
rect 364432 700266 364484 700272
rect 302884 455524 302936 455530
rect 302884 455466 302936 455472
rect 299480 453416 299532 453422
rect 299480 453358 299532 453364
rect 300124 451920 300176 451926
rect 300124 451862 300176 451868
rect 299388 403640 299440 403646
rect 299388 403582 299440 403588
rect 298388 379486 298784 379514
rect 297548 375488 297600 375494
rect 297548 375430 297600 375436
rect 297456 375420 297508 375426
rect 297456 375362 297508 375368
rect 297560 374898 297588 375430
rect 297732 375420 297784 375426
rect 297732 375362 297784 375368
rect 297468 374870 297588 374898
rect 297088 374400 297140 374406
rect 297088 374342 297140 374348
rect 295524 374128 295576 374134
rect 295524 374070 295576 374076
rect 294788 373516 294840 373522
rect 294788 373458 294840 373464
rect 295536 373182 295564 374070
rect 295616 373380 295668 373386
rect 295616 373322 295668 373328
rect 295524 373176 295576 373182
rect 295524 373118 295576 373124
rect 295248 372292 295300 372298
rect 295248 372234 295300 372240
rect 295260 371890 295288 372234
rect 295248 371884 295300 371890
rect 295248 371826 295300 371832
rect 294604 370524 294656 370530
rect 294604 370466 294656 370472
rect 295260 369866 295288 371826
rect 294432 369838 294676 369866
rect 295044 369838 295288 369866
rect 292836 369702 293080 369730
rect 295536 369594 295564 373118
rect 295628 373046 295656 373322
rect 296628 373312 296680 373318
rect 296628 373254 296680 373260
rect 295616 373040 295668 373046
rect 295616 372982 295668 372988
rect 296352 370796 296404 370802
rect 296352 370738 296404 370744
rect 295984 370660 296036 370666
rect 295984 370602 296036 370608
rect 295996 369866 296024 370602
rect 296364 370190 296392 370738
rect 296352 370184 296404 370190
rect 296352 370126 296404 370132
rect 296364 369866 296392 370126
rect 295780 369838 296024 369866
rect 296148 369838 296392 369866
rect 296640 369730 296668 373254
rect 297100 369866 297128 374342
rect 297468 369866 297496 374870
rect 297548 373380 297600 373386
rect 297548 373322 297600 373328
rect 297560 370002 297588 373322
rect 297560 369974 297634 370002
rect 296884 369838 297128 369866
rect 297252 369838 297496 369866
rect 297606 369852 297634 369974
rect 297744 369866 297772 375362
rect 298388 375018 298416 379486
rect 298376 375012 298428 375018
rect 298376 374954 298428 374960
rect 298388 370138 298416 374954
rect 300136 374134 300164 451862
rect 300308 450764 300360 450770
rect 300308 450706 300360 450712
rect 300214 449168 300270 449177
rect 300214 449103 300270 449112
rect 300124 374128 300176 374134
rect 300124 374070 300176 374076
rect 298468 373448 298520 373454
rect 298468 373390 298520 373396
rect 298480 373114 298508 373390
rect 298468 373108 298520 373114
rect 298468 373050 298520 373056
rect 298342 370110 298416 370138
rect 297744 369838 297988 369866
rect 298342 369852 298370 370110
rect 298480 369866 298508 373050
rect 300228 372978 300256 449103
rect 300320 376106 300348 450706
rect 301504 450356 301556 450362
rect 301504 450298 301556 450304
rect 300398 401024 300454 401033
rect 300398 400959 300454 400968
rect 300308 376100 300360 376106
rect 300308 376042 300360 376048
rect 300216 372972 300268 372978
rect 300216 372914 300268 372920
rect 299204 372768 299256 372774
rect 299204 372710 299256 372716
rect 299216 371210 299244 372710
rect 299204 371204 299256 371210
rect 299204 371146 299256 371152
rect 298836 370728 298888 370734
rect 298836 370670 298888 370676
rect 298848 370326 298876 370670
rect 298836 370320 298888 370326
rect 298836 370262 298888 370268
rect 298848 369866 298876 370262
rect 299216 369866 299244 371146
rect 300228 370104 300256 372914
rect 300044 370076 300256 370104
rect 300044 369866 300072 370076
rect 300320 369866 300348 376042
rect 300412 375630 300440 400959
rect 301516 379514 301544 450298
rect 301594 399800 301650 399809
rect 301594 399735 301650 399744
rect 301332 379486 301544 379514
rect 300400 375624 300452 375630
rect 300400 375566 300452 375572
rect 298480 369838 298724 369866
rect 298848 369838 299092 369866
rect 299216 369838 299460 369866
rect 299828 369838 300072 369866
rect 300196 369838 300348 369866
rect 300412 369866 300440 375566
rect 300860 374740 300912 374746
rect 300860 374682 300912 374688
rect 300872 370138 300900 374682
rect 301332 372910 301360 379486
rect 301608 374746 301636 399735
rect 301964 377460 302016 377466
rect 301964 377402 302016 377408
rect 301596 374740 301648 374746
rect 301596 374682 301648 374688
rect 301976 374610 302004 377402
rect 302896 376922 302924 455466
rect 304276 439521 304304 700266
rect 363604 698692 363656 698698
rect 363604 698634 363656 698640
rect 360108 670744 360160 670750
rect 360108 670686 360160 670692
rect 359464 643136 359516 643142
rect 359464 643078 359516 643084
rect 311164 618316 311216 618322
rect 311164 618258 311216 618264
rect 311176 456958 311204 618258
rect 358084 576904 358136 576910
rect 358084 576846 358136 576852
rect 355324 484424 355376 484430
rect 355324 484366 355376 484372
rect 315304 462392 315356 462398
rect 315304 462334 315356 462340
rect 315316 457094 315344 462334
rect 334716 457292 334768 457298
rect 334716 457234 334768 457240
rect 323768 457224 323820 457230
rect 323768 457166 323820 457172
rect 320916 457156 320968 457162
rect 320916 457098 320968 457104
rect 315304 457088 315356 457094
rect 315304 457030 315356 457036
rect 311164 456952 311216 456958
rect 311164 456894 311216 456900
rect 311808 456952 311860 456958
rect 311808 456894 311860 456900
rect 308402 454200 308458 454209
rect 308402 454135 308458 454144
rect 305000 450696 305052 450702
rect 305000 450638 305052 450644
rect 305012 450090 305040 450638
rect 306380 450560 306432 450566
rect 306380 450502 306432 450508
rect 305000 450084 305052 450090
rect 305000 450026 305052 450032
rect 304356 449268 304408 449274
rect 304356 449210 304408 449216
rect 304262 439512 304318 439521
rect 304262 439447 304318 439456
rect 303526 401160 303582 401169
rect 303526 401095 303582 401104
rect 302608 376916 302660 376922
rect 302608 376858 302660 376864
rect 302884 376916 302936 376922
rect 302884 376858 302936 376864
rect 301964 374604 302016 374610
rect 301964 374546 302016 374552
rect 301320 372904 301372 372910
rect 301320 372846 301372 372852
rect 301332 370138 301360 372846
rect 301412 370932 301464 370938
rect 301412 370874 301464 370880
rect 301424 370462 301452 370874
rect 301412 370456 301464 370462
rect 301412 370398 301464 370404
rect 300872 370110 300946 370138
rect 300412 369838 300564 369866
rect 300918 369852 300946 370110
rect 301286 370110 301360 370138
rect 301286 369852 301314 370110
rect 301424 369866 301452 370398
rect 301976 370138 302004 374546
rect 301976 370110 302050 370138
rect 301424 369838 301668 369866
rect 302022 369852 302050 370110
rect 302378 370116 302430 370122
rect 302378 370058 302430 370064
rect 302390 369852 302418 370058
rect 302620 369866 302648 376858
rect 303436 372700 303488 372706
rect 303436 372642 303488 372648
rect 303448 372570 303476 372642
rect 303436 372564 303488 372570
rect 303436 372506 303488 372512
rect 302884 371748 302936 371754
rect 302884 371690 302936 371696
rect 302896 371482 302924 371690
rect 302884 371476 302936 371482
rect 302884 371418 302936 371424
rect 303448 370954 303476 372506
rect 303540 371414 303568 401095
rect 303620 398540 303672 398546
rect 303620 398482 303672 398488
rect 303632 395690 303660 398482
rect 304276 398206 304304 439447
rect 304264 398200 304316 398206
rect 304264 398142 304316 398148
rect 303620 395684 303672 395690
rect 303620 395626 303672 395632
rect 303618 384296 303674 384305
rect 303618 384231 303674 384240
rect 303632 379642 303660 384231
rect 303620 379636 303672 379642
rect 303620 379578 303672 379584
rect 303528 371408 303580 371414
rect 303528 371350 303580 371356
rect 303356 370926 303476 370954
rect 303356 369866 303384 370926
rect 303436 370864 303488 370870
rect 303436 370806 303488 370812
rect 303448 370122 303476 370806
rect 303436 370116 303488 370122
rect 303436 370058 303488 370064
rect 302620 369838 302772 369866
rect 303140 369838 303384 369866
rect 303632 369866 303660 379578
rect 304368 374474 304396 449210
rect 305012 374626 305040 450026
rect 305734 399664 305790 399673
rect 305734 399599 305790 399608
rect 305092 398608 305144 398614
rect 305092 398550 305144 398556
rect 305104 395622 305132 398550
rect 305644 398200 305696 398206
rect 305644 398142 305696 398148
rect 305092 395616 305144 395622
rect 305092 395558 305144 395564
rect 305656 387530 305684 398142
rect 305092 387524 305144 387530
rect 305092 387466 305144 387472
rect 305644 387524 305696 387530
rect 305644 387466 305696 387472
rect 305104 381002 305132 387466
rect 305092 380996 305144 381002
rect 305092 380938 305144 380944
rect 305104 379514 305132 380938
rect 305104 379486 305684 379514
rect 305012 374598 305132 374626
rect 304356 374468 304408 374474
rect 304356 374410 304408 374416
rect 303988 371408 304040 371414
rect 303988 371350 304040 371356
rect 303632 369838 303876 369866
rect 304000 369753 304028 371350
rect 304368 370138 304396 374410
rect 304816 373992 304868 373998
rect 304816 373934 304868 373940
rect 304828 372842 304856 373934
rect 304816 372836 304868 372842
rect 304816 372778 304868 372784
rect 304724 371952 304776 371958
rect 304724 371894 304776 371900
rect 304230 370110 304396 370138
rect 304230 369852 304258 370110
rect 304356 369912 304408 369918
rect 304356 369854 304408 369860
rect 296516 369702 296668 369730
rect 303480 369744 303536 369753
rect 303480 369679 303536 369688
rect 303986 369744 304042 369753
rect 304368 369730 304396 369854
rect 304736 369730 304764 371894
rect 304368 369702 304764 369730
rect 304828 369730 304856 372778
rect 304828 369702 304980 369730
rect 303986 369679 304042 369688
rect 295412 369566 295564 369594
rect 304000 369442 304028 369679
rect 305104 369510 305132 374598
rect 305552 374536 305604 374542
rect 305552 374478 305604 374484
rect 305564 374202 305592 374478
rect 305552 374196 305604 374202
rect 305552 374138 305604 374144
rect 305564 369866 305592 374138
rect 305656 370274 305684 379486
rect 305748 374542 305776 399599
rect 306288 397044 306340 397050
rect 306288 396986 306340 396992
rect 305736 374536 305788 374542
rect 305736 374478 305788 374484
rect 305656 370246 305868 370274
rect 305348 369838 305592 369866
rect 305840 369866 305868 370246
rect 305840 369838 306084 369866
rect 305092 369504 305144 369510
rect 305092 369446 305144 369452
rect 305460 369504 305512 369510
rect 306300 369481 306328 396986
rect 306392 379778 306420 450502
rect 307666 449984 307722 449993
rect 307666 449919 307722 449928
rect 307024 449336 307076 449342
rect 307024 449278 307076 449284
rect 306380 379772 306432 379778
rect 306380 379714 306432 379720
rect 306564 379772 306616 379778
rect 306564 379714 306616 379720
rect 306426 370116 306478 370122
rect 306426 370058 306478 370064
rect 306438 369852 306466 370058
rect 306576 369866 306604 379714
rect 307036 374270 307064 449278
rect 307680 404297 307708 449919
rect 307666 404288 307722 404297
rect 307666 404223 307722 404232
rect 308416 383654 308444 454135
rect 308496 451988 308548 451994
rect 308496 451930 308548 451936
rect 308324 383626 308444 383654
rect 307668 378820 307720 378826
rect 307668 378762 307720 378768
rect 307300 374808 307352 374814
rect 307300 374750 307352 374756
rect 307024 374264 307076 374270
rect 307024 374206 307076 374212
rect 306932 372700 306984 372706
rect 306932 372642 306984 372648
rect 306944 372026 306972 372642
rect 306932 372020 306984 372026
rect 306932 371962 306984 371968
rect 306576 369838 306820 369866
rect 306944 369594 306972 371962
rect 307036 370122 307064 374206
rect 307024 370116 307076 370122
rect 307024 370058 307076 370064
rect 307312 369866 307340 374750
rect 307312 369838 307556 369866
rect 306944 369566 307188 369594
rect 307680 369481 307708 378762
rect 308324 371822 308352 383626
rect 308404 374332 308456 374338
rect 308404 374274 308456 374280
rect 308312 371816 308364 371822
rect 308312 371758 308364 371764
rect 307760 371000 307812 371006
rect 307760 370942 307812 370948
rect 307772 369866 307800 370942
rect 308324 370138 308352 371758
rect 308278 370110 308352 370138
rect 307772 369838 307924 369866
rect 308278 369852 308306 370110
rect 308416 369866 308444 374274
rect 308508 372706 308536 451930
rect 309784 451580 309836 451586
rect 309784 451522 309836 451528
rect 309138 450528 309194 450537
rect 309138 450463 309194 450472
rect 309152 379914 309180 450463
rect 309140 379908 309192 379914
rect 309140 379850 309192 379856
rect 309324 379908 309376 379914
rect 309324 379850 309376 379856
rect 309336 379514 309364 379850
rect 309336 379486 309732 379514
rect 309598 375456 309654 375465
rect 309598 375391 309654 375400
rect 308496 372700 308548 372706
rect 308496 372642 308548 372648
rect 309508 372496 309560 372502
rect 309508 372438 309560 372444
rect 309520 371550 309548 372438
rect 309508 371544 309560 371550
rect 308770 371512 308826 371521
rect 309508 371486 309560 371492
rect 308770 371447 308826 371456
rect 308784 369866 308812 371447
rect 309520 369866 309548 371486
rect 308416 369838 308660 369866
rect 308784 369838 309028 369866
rect 309396 369838 309548 369866
rect 309612 369866 309640 375391
rect 309704 370138 309732 379486
rect 309796 373998 309824 451522
rect 309874 450120 309930 450129
rect 309874 450055 309930 450064
rect 309784 373992 309836 373998
rect 309784 373934 309836 373940
rect 309888 372314 309916 450055
rect 311164 422340 311216 422346
rect 311164 422282 311216 422288
rect 311176 415478 311204 422282
rect 311164 415472 311216 415478
rect 311164 415414 311216 415420
rect 311256 410576 311308 410582
rect 311256 410518 311308 410524
rect 309968 406428 310020 406434
rect 309968 406370 310020 406376
rect 309980 405618 310008 406370
rect 309968 405612 310020 405618
rect 309968 405554 310020 405560
rect 309980 372502 310008 405554
rect 310520 403640 310572 403646
rect 310520 403582 310572 403588
rect 310060 399628 310112 399634
rect 310060 399570 310112 399576
rect 310072 375465 310100 399570
rect 310058 375456 310114 375465
rect 310058 375391 310114 375400
rect 310532 372609 310560 403582
rect 311268 401577 311296 410518
rect 311820 402974 311848 456894
rect 314016 450424 314068 450430
rect 314016 450366 314068 450372
rect 312542 449032 312598 449041
rect 312542 448967 312598 448976
rect 311900 411936 311952 411942
rect 311900 411878 311952 411884
rect 311912 411262 311940 411878
rect 311900 411256 311952 411262
rect 311900 411198 311952 411204
rect 311820 402946 312124 402974
rect 311254 401568 311310 401577
rect 311254 401503 311310 401512
rect 311164 399560 311216 399566
rect 311164 399502 311216 399508
rect 311176 383654 311204 399502
rect 310900 383626 311204 383654
rect 310900 376038 310928 383626
rect 311268 381138 311296 401503
rect 311808 391468 311860 391474
rect 311808 391410 311860 391416
rect 311256 381132 311308 381138
rect 311256 381074 311308 381080
rect 310888 376032 310940 376038
rect 310888 375974 310940 375980
rect 310518 372600 310574 372609
rect 310518 372535 310574 372544
rect 309968 372496 310020 372502
rect 309968 372438 310020 372444
rect 309888 372286 310284 372314
rect 310256 371793 310284 372286
rect 310242 371784 310298 371793
rect 310242 371719 310298 371728
rect 309704 370110 309916 370138
rect 309888 369866 309916 370110
rect 310256 369866 310284 371719
rect 310900 370138 310928 375974
rect 311268 370138 311296 381074
rect 311346 372600 311402 372609
rect 311346 372535 311402 372544
rect 310854 370110 310928 370138
rect 311222 370110 311296 370138
rect 309612 369838 309764 369866
rect 309888 369838 310132 369866
rect 310256 369838 310500 369866
rect 310854 369852 310882 370110
rect 311222 369852 311250 370110
rect 311360 369866 311388 372535
rect 311360 369838 311604 369866
rect 311820 369481 311848 391410
rect 312096 370394 312124 402946
rect 312556 383654 312584 448967
rect 313924 414724 313976 414730
rect 313924 414666 313976 414672
rect 313936 413982 313964 414666
rect 313924 413976 313976 413982
rect 313924 413918 313976 413924
rect 313280 413908 313332 413914
rect 313280 413850 313332 413856
rect 312636 411256 312688 411262
rect 312636 411198 312688 411204
rect 312188 383626 312584 383654
rect 312188 375970 312216 383626
rect 312648 379514 312676 411198
rect 313292 402974 313320 413850
rect 313292 402946 313504 402974
rect 313280 402280 313332 402286
rect 313280 402222 313332 402228
rect 313292 401606 313320 402222
rect 313280 401600 313332 401606
rect 313280 401542 313332 401548
rect 312728 399492 312780 399498
rect 312728 399434 312780 399440
rect 312464 379486 312676 379514
rect 312740 379514 312768 399434
rect 313188 390652 313240 390658
rect 313188 390594 313240 390600
rect 312740 379486 312860 379514
rect 312176 375964 312228 375970
rect 312176 375906 312228 375912
rect 312084 370388 312136 370394
rect 312084 370330 312136 370336
rect 312096 370122 312124 370330
rect 312084 370116 312136 370122
rect 312084 370058 312136 370064
rect 312188 369730 312216 375906
rect 311972 369702 312216 369730
rect 306286 369472 306342 369481
rect 305512 369452 305716 369458
rect 305460 369446 305716 369452
rect 287288 369407 287344 369416
rect 291108 369436 291160 369442
rect 291108 369378 291160 369384
rect 292304 369436 292356 369442
rect 292304 369378 292356 369384
rect 303988 369436 304040 369442
rect 305472 369430 305716 369446
rect 306286 369407 306342 369416
rect 307666 369472 307722 369481
rect 307666 369407 307722 369416
rect 311806 369472 311862 369481
rect 311806 369407 311862 369416
rect 312312 369472 312368 369481
rect 312464 369458 312492 379486
rect 312832 375902 312860 379486
rect 312820 375896 312872 375902
rect 312820 375838 312872 375844
rect 312682 370116 312734 370122
rect 312682 370058 312734 370064
rect 312694 369852 312722 370058
rect 312832 369866 312860 375838
rect 313200 370161 313228 390594
rect 313476 382430 313504 402946
rect 313936 383654 313964 413918
rect 314028 413914 314056 450366
rect 314752 416764 314804 416770
rect 314752 416706 314804 416712
rect 314016 413908 314068 413914
rect 314016 413850 314068 413856
rect 314016 401600 314068 401606
rect 314016 401542 314068 401548
rect 313924 383648 313976 383654
rect 313924 383590 313976 383596
rect 313464 382424 313516 382430
rect 313464 382366 313516 382372
rect 313186 370152 313242 370161
rect 313476 370138 313504 382366
rect 314028 371482 314056 401542
rect 314106 400888 314162 400897
rect 314106 400823 314162 400832
rect 314120 378282 314148 400823
rect 314384 390584 314436 390590
rect 314384 390526 314436 390532
rect 314200 383648 314252 383654
rect 314200 383590 314252 383596
rect 314108 378276 314160 378282
rect 314108 378218 314160 378224
rect 314016 371476 314068 371482
rect 314016 371418 314068 371424
rect 313186 370087 313242 370096
rect 313430 370110 313504 370138
rect 312832 369838 313076 369866
rect 313430 369852 313458 370110
rect 314028 369866 314056 371418
rect 314120 370002 314148 378218
rect 314212 370258 314240 383590
rect 314200 370252 314252 370258
rect 314200 370194 314252 370200
rect 314212 370122 314240 370194
rect 314200 370116 314252 370122
rect 314200 370058 314252 370064
rect 314120 369974 314194 370002
rect 313812 369838 314056 369866
rect 314166 369852 314194 369974
rect 314396 369481 314424 390526
rect 314764 379846 314792 416706
rect 314844 383104 314896 383110
rect 314844 383046 314896 383052
rect 314856 382294 314884 383046
rect 314844 382288 314896 382294
rect 314844 382230 314896 382236
rect 314752 379840 314804 379846
rect 314752 379782 314804 379788
rect 314764 374678 314792 379782
rect 314752 374672 314804 374678
rect 314752 374614 314804 374620
rect 314856 370138 314884 382230
rect 315316 379514 315344 457030
rect 320824 457020 320876 457026
rect 320824 456962 320876 456968
rect 319536 454912 319588 454918
rect 319536 454854 319588 454860
rect 318248 454368 318300 454374
rect 318248 454310 318300 454316
rect 316868 454300 316920 454306
rect 316868 454242 316920 454248
rect 315396 453212 315448 453218
rect 315396 453154 315448 453160
rect 315408 416770 315436 453154
rect 316684 453144 316736 453150
rect 316684 453086 316736 453092
rect 315488 417444 315540 417450
rect 315488 417386 315540 417392
rect 315396 416764 315448 416770
rect 315396 416706 315448 416712
rect 315500 404326 315528 417386
rect 316040 405680 316092 405686
rect 316040 405622 316092 405628
rect 315488 404320 315540 404326
rect 315488 404262 315540 404268
rect 315394 399936 315450 399945
rect 315394 399871 315450 399880
rect 315224 379486 315344 379514
rect 315224 372502 315252 379486
rect 315408 376786 315436 399871
rect 315500 383110 315528 404262
rect 315856 393032 315908 393038
rect 315856 392974 315908 392980
rect 315488 383104 315540 383110
rect 315488 383046 315540 383052
rect 315396 376780 315448 376786
rect 315396 376722 315448 376728
rect 315408 375442 315436 376722
rect 315316 375414 315436 375442
rect 315212 372496 315264 372502
rect 315212 372438 315264 372444
rect 315316 370138 315344 375414
rect 315396 374672 315448 374678
rect 315396 374614 315448 374620
rect 314522 370116 314574 370122
rect 314856 370110 314930 370138
rect 314522 370058 314574 370064
rect 314534 369852 314562 370058
rect 314902 369852 314930 370110
rect 315270 370110 315344 370138
rect 315270 369852 315298 370110
rect 315408 369866 315436 374614
rect 315764 372496 315816 372502
rect 315764 372438 315816 372444
rect 315776 371686 315804 372438
rect 315764 371680 315816 371686
rect 315764 371622 315816 371628
rect 315408 369838 315652 369866
rect 315776 369730 315804 371622
rect 315868 369889 315896 392974
rect 316052 372298 316080 405622
rect 316132 401668 316184 401674
rect 316132 401610 316184 401616
rect 316144 379710 316172 401610
rect 316696 385082 316724 453086
rect 316776 453008 316828 453014
rect 316776 452950 316828 452956
rect 316788 415478 316816 452950
rect 316776 415472 316828 415478
rect 316776 415414 316828 415420
rect 316788 401674 316816 415414
rect 316880 405686 316908 454242
rect 318064 453552 318116 453558
rect 318064 453494 318116 453500
rect 316868 405680 316920 405686
rect 316868 405622 316920 405628
rect 316776 401668 316828 401674
rect 316776 401610 316828 401616
rect 317694 385792 317750 385801
rect 317694 385727 317750 385736
rect 316224 385076 316276 385082
rect 316224 385018 316276 385024
rect 316684 385076 316736 385082
rect 316684 385018 316736 385024
rect 316236 383654 316264 385018
rect 316236 383626 316540 383654
rect 316132 379704 316184 379710
rect 316132 379646 316184 379652
rect 316040 372292 316092 372298
rect 316040 372234 316092 372240
rect 316052 371618 316080 372234
rect 316040 371612 316092 371618
rect 316040 371554 316092 371560
rect 315854 369880 315910 369889
rect 316144 369866 316172 379646
rect 316512 369866 316540 383626
rect 317512 381200 317564 381206
rect 317512 381142 317564 381148
rect 317524 378418 317552 381142
rect 317604 379024 317656 379030
rect 317604 378966 317656 378972
rect 317512 378412 317564 378418
rect 317512 378354 317564 378360
rect 317616 378350 317644 378966
rect 317604 378344 317656 378350
rect 317604 378286 317656 378292
rect 316868 372292 316920 372298
rect 316868 372234 316920 372240
rect 316880 369866 316908 372234
rect 317616 369866 317644 378286
rect 317708 370054 317736 385727
rect 317972 378412 318024 378418
rect 317972 378354 318024 378360
rect 317696 370048 317748 370054
rect 317696 369990 317748 369996
rect 316144 369838 316388 369866
rect 316512 369838 316756 369866
rect 316880 369838 317124 369866
rect 317492 369838 317644 369866
rect 317708 369866 317736 369990
rect 317984 369866 318012 378354
rect 318076 370598 318104 453494
rect 318156 453076 318208 453082
rect 318156 453018 318208 453024
rect 318168 379030 318196 453018
rect 318260 381206 318288 454310
rect 319444 450628 319496 450634
rect 319444 450570 319496 450576
rect 319168 390176 319220 390182
rect 319168 390118 319220 390124
rect 318708 389224 318760 389230
rect 318708 389166 318760 389172
rect 318248 381200 318300 381206
rect 318248 381142 318300 381148
rect 318720 379514 318748 389166
rect 319076 385008 319128 385014
rect 319076 384950 319128 384956
rect 319088 383722 319116 384950
rect 319076 383716 319128 383722
rect 319076 383658 319128 383664
rect 318892 383036 318944 383042
rect 318892 382978 318944 382984
rect 318904 382498 318932 382978
rect 318984 382628 319036 382634
rect 318984 382570 319036 382576
rect 318892 382492 318944 382498
rect 318892 382434 318944 382440
rect 318444 379486 318748 379514
rect 318156 379024 318208 379030
rect 318156 378966 318208 378972
rect 318064 370592 318116 370598
rect 318064 370534 318116 370540
rect 317708 369838 317860 369866
rect 317984 369838 318228 369866
rect 315854 369815 315910 369824
rect 315776 369702 316020 369730
rect 318444 369481 318472 379486
rect 318904 371142 318932 382434
rect 318996 382362 319024 382570
rect 318984 382356 319036 382362
rect 318984 382298 319036 382304
rect 318892 371136 318944 371142
rect 318892 371078 318944 371084
rect 318708 370592 318760 370598
rect 318708 370534 318760 370540
rect 318720 369730 318748 370534
rect 318996 370122 319024 382298
rect 318984 370116 319036 370122
rect 318984 370058 319036 370064
rect 319088 369866 319116 383658
rect 319180 383654 319208 390118
rect 319180 383626 319300 383654
rect 319272 374660 319300 383626
rect 319456 379514 319484 450570
rect 319548 382634 319576 454854
rect 319628 454572 319680 454578
rect 319628 454514 319680 454520
rect 319640 383042 319668 454514
rect 319720 454504 319772 454510
rect 319720 454446 319772 454452
rect 319732 385014 319760 454446
rect 319812 390108 319864 390114
rect 319812 390050 319864 390056
rect 319720 385008 319772 385014
rect 319720 384950 319772 384956
rect 319628 383036 319680 383042
rect 319628 382978 319680 382984
rect 319536 382628 319588 382634
rect 319536 382570 319588 382576
rect 319456 379486 319576 379514
rect 319548 374950 319576 379486
rect 319536 374944 319588 374950
rect 319536 374886 319588 374892
rect 319272 374632 319484 374660
rect 319168 371136 319220 371142
rect 319168 371078 319220 371084
rect 318964 369838 319116 369866
rect 319180 369866 319208 371078
rect 319456 369889 319484 374632
rect 319442 369880 319498 369889
rect 319180 369838 319332 369866
rect 319548 369866 319576 374886
rect 319548 369838 319700 369866
rect 319442 369815 319498 369824
rect 318596 369702 318748 369730
rect 319824 369617 319852 390050
rect 319904 390040 319956 390046
rect 319904 389982 319956 389988
rect 319810 369608 319866 369617
rect 319810 369543 319866 369552
rect 319916 369481 319944 389982
rect 320456 386368 320508 386374
rect 320456 386310 320508 386316
rect 320468 385218 320496 386310
rect 320456 385212 320508 385218
rect 320456 385154 320508 385160
rect 320468 383654 320496 385154
rect 320468 383626 320772 383654
rect 320364 379568 320416 379574
rect 320364 379514 320416 379516
rect 320364 379510 320588 379514
rect 320376 379486 320588 379510
rect 320272 371408 320324 371414
rect 320272 371350 320324 371356
rect 320042 370116 320094 370122
rect 320042 370058 320094 370064
rect 320054 369852 320082 370058
rect 320284 369594 320312 371350
rect 320560 369866 320588 379486
rect 320744 370138 320772 383626
rect 320836 372434 320864 456962
rect 320928 386374 320956 457098
rect 322296 455456 322348 455462
rect 322296 455398 322348 455404
rect 322204 452872 322256 452878
rect 322204 452814 322256 452820
rect 321008 450696 321060 450702
rect 321008 450638 321060 450644
rect 320916 386368 320968 386374
rect 320916 386310 320968 386316
rect 321020 379574 321048 450638
rect 321376 393372 321428 393378
rect 321376 393314 321428 393320
rect 321008 379568 321060 379574
rect 321008 379510 321060 379516
rect 320824 372428 320876 372434
rect 320824 372370 320876 372376
rect 320744 370110 320956 370138
rect 320928 369866 320956 370110
rect 320560 369838 320804 369866
rect 320928 369838 321172 369866
rect 320284 369566 320436 369594
rect 321388 369481 321416 393314
rect 321744 387796 321796 387802
rect 321744 387738 321796 387744
rect 321756 386510 321784 387738
rect 321744 386504 321796 386510
rect 321744 386446 321796 386452
rect 321756 383654 321784 386446
rect 321756 383626 322060 383654
rect 321652 382560 321704 382566
rect 321652 382502 321704 382508
rect 321664 374678 321692 382502
rect 321836 375556 321888 375562
rect 321836 375498 321888 375504
rect 321652 374672 321704 374678
rect 321652 374614 321704 374620
rect 321468 372428 321520 372434
rect 321468 372370 321520 372376
rect 321480 370138 321508 372370
rect 321848 370138 321876 375498
rect 321480 370110 321554 370138
rect 321848 370110 321922 370138
rect 321526 369852 321554 370110
rect 321894 369852 321922 370110
rect 322032 369866 322060 383626
rect 322216 375562 322244 452814
rect 322308 383858 322336 455398
rect 323584 453620 323636 453626
rect 323584 453562 323636 453568
rect 322388 438184 322440 438190
rect 322388 438126 322440 438132
rect 322296 383852 322348 383858
rect 322296 383794 322348 383800
rect 322204 375556 322256 375562
rect 322204 375498 322256 375504
rect 322308 370122 322336 383794
rect 322400 382566 322428 438126
rect 322478 399528 322534 399537
rect 322478 399463 322534 399472
rect 322492 387802 322520 399463
rect 322848 394392 322900 394398
rect 322848 394334 322900 394340
rect 322480 387796 322532 387802
rect 322480 387738 322532 387744
rect 322388 382560 322440 382566
rect 322388 382502 322440 382508
rect 322388 374672 322440 374678
rect 322388 374614 322440 374620
rect 322296 370116 322348 370122
rect 322296 370058 322348 370064
rect 322400 369866 322428 374614
rect 322032 369838 322276 369866
rect 322400 369838 322644 369866
rect 322860 369481 322888 394334
rect 322940 378208 322992 378214
rect 322940 378150 322992 378156
rect 322952 370138 322980 378150
rect 323596 376854 323624 453562
rect 323676 450492 323728 450498
rect 323676 450434 323728 450440
rect 323688 378214 323716 450434
rect 323780 385150 323808 457166
rect 334624 455932 334676 455938
rect 334624 455874 334676 455880
rect 332140 455864 332192 455870
rect 332140 455806 332192 455812
rect 332048 455796 332100 455802
rect 332048 455738 332100 455744
rect 324964 452804 325016 452810
rect 324964 452746 325016 452752
rect 323768 385144 323820 385150
rect 323768 385086 323820 385092
rect 323676 378208 323728 378214
rect 323676 378150 323728 378156
rect 323584 376848 323636 376854
rect 323584 376790 323636 376796
rect 323780 372502 323808 385086
rect 324976 382022 325004 452746
rect 331494 449576 331550 449585
rect 331494 449511 331550 449520
rect 330208 449268 330260 449274
rect 330208 449210 330260 449216
rect 330220 449138 330248 449210
rect 330208 449132 330260 449138
rect 330208 449074 330260 449080
rect 331508 448769 331536 449511
rect 331494 448760 331550 448769
rect 331494 448695 331550 448704
rect 325056 445052 325108 445058
rect 325056 444994 325108 445000
rect 324412 382016 324464 382022
rect 324412 381958 324464 381964
rect 324964 382016 325016 382022
rect 324964 381958 325016 381964
rect 324424 380934 324452 381958
rect 325068 380934 325096 444994
rect 326344 407788 326396 407794
rect 326344 407730 326396 407736
rect 326356 385014 326384 407730
rect 331864 399696 331916 399702
rect 331864 399638 331916 399644
rect 330760 398676 330812 398682
rect 330760 398618 330812 398624
rect 330668 397248 330720 397254
rect 330668 397190 330720 397196
rect 330576 395752 330628 395758
rect 330576 395694 330628 395700
rect 329288 395684 329340 395690
rect 329288 395626 329340 395632
rect 328000 395208 328052 395214
rect 328000 395150 328052 395156
rect 325700 385008 325752 385014
rect 325700 384950 325752 384956
rect 326344 385008 326396 385014
rect 326344 384950 326396 384956
rect 325712 383790 325740 384950
rect 325700 383784 325752 383790
rect 325700 383726 325752 383732
rect 324412 380928 324464 380934
rect 324412 380870 324464 380876
rect 324596 380928 324648 380934
rect 324596 380870 324648 380876
rect 325056 380928 325108 380934
rect 325056 380870 325108 380876
rect 323860 376848 323912 376854
rect 323860 376790 323912 376796
rect 323768 372496 323820 372502
rect 323768 372438 323820 372444
rect 323584 371272 323636 371278
rect 323584 371214 323636 371220
rect 322952 370110 323026 370138
rect 322998 369852 323026 370110
rect 323354 370116 323406 370122
rect 323354 370058 323406 370064
rect 323366 369852 323394 370058
rect 323596 369594 323624 371214
rect 323872 369866 323900 376790
rect 324424 374678 324452 380870
rect 324412 374672 324464 374678
rect 324412 374614 324464 374620
rect 324320 372496 324372 372502
rect 324320 372438 324372 372444
rect 324332 369866 324360 372438
rect 324608 369866 324636 380870
rect 324964 374672 325016 374678
rect 324964 374614 325016 374620
rect 324976 369866 325004 374614
rect 325424 371340 325476 371346
rect 325424 371282 325476 371288
rect 323872 369838 324116 369866
rect 324332 369838 324484 369866
rect 324608 369838 324852 369866
rect 324976 369838 325220 369866
rect 325436 369594 325464 371282
rect 325712 369866 325740 383726
rect 327724 372360 327776 372366
rect 327724 372302 327776 372308
rect 325712 369838 325956 369866
rect 323596 369566 323748 369594
rect 325436 369566 325588 369594
rect 312368 369430 312492 369458
rect 314382 369472 314438 369481
rect 312312 369407 312368 369416
rect 314382 369407 314438 369416
rect 318430 369472 318486 369481
rect 318430 369407 318486 369416
rect 319902 369472 319958 369481
rect 319902 369407 319958 369416
rect 321374 369472 321430 369481
rect 321374 369407 321430 369416
rect 322846 369472 322902 369481
rect 322846 369407 322902 369416
rect 303988 369378 304040 369384
rect 288024 369336 288080 369345
rect 288024 369271 288080 369280
rect 289128 369336 289184 369345
rect 289128 369271 289184 369280
rect 312312 369336 312368 369345
rect 312312 369271 312368 369280
rect 327736 360913 327764 372302
rect 327722 360904 327778 360913
rect 327722 360839 327778 360848
rect 327722 359408 327778 359417
rect 327722 359343 327778 359352
rect 327446 355328 327502 355337
rect 327446 355263 327502 355272
rect 282458 352608 282514 352617
rect 282458 352543 282514 352552
rect 327460 321910 327488 355263
rect 327538 330440 327594 330449
rect 327538 330375 327594 330384
rect 327448 321904 327500 321910
rect 327448 321846 327500 321852
rect 282366 321600 282422 321609
rect 282366 321535 282422 321544
rect 282458 321464 282514 321473
rect 282458 321399 282514 321408
rect 282472 321065 282500 321399
rect 282458 321056 282514 321065
rect 282458 320991 282514 321000
rect 282688 320784 282744 320793
rect 282688 320719 282744 320728
rect 283976 320784 284032 320793
rect 283976 320719 284032 320728
rect 284344 320784 284400 320793
rect 284344 320719 284400 320728
rect 285540 320784 285596 320793
rect 288392 320784 288448 320793
rect 285922 320754 285950 320756
rect 285540 320719 285596 320728
rect 285910 320748 285962 320754
rect 288392 320719 288448 320728
rect 289128 320784 289184 320793
rect 289128 320719 289184 320728
rect 289312 320784 289368 320793
rect 289312 320719 289368 320728
rect 289864 320784 289920 320793
rect 291428 320784 291484 320793
rect 290246 320754 290274 320756
rect 289864 320719 289920 320728
rect 290234 320748 290286 320754
rect 285910 320690 285962 320696
rect 291428 320719 291484 320728
rect 295384 320784 295440 320793
rect 295384 320719 295440 320728
rect 297040 320784 297096 320793
rect 297040 320719 297096 320728
rect 301272 320784 301328 320793
rect 301272 320719 301328 320728
rect 304032 320784 304088 320793
rect 304032 320719 304088 320728
rect 304768 320784 304824 320793
rect 304768 320719 304824 320728
rect 307528 320784 307584 320793
rect 307528 320719 307584 320728
rect 311116 320784 311172 320793
rect 311116 320719 311172 320728
rect 314796 320784 314852 320793
rect 314796 320719 314798 320728
rect 290234 320690 290286 320696
rect 314850 320719 314852 320728
rect 315808 320784 315864 320793
rect 315808 320719 315864 320728
rect 318476 320784 318532 320793
rect 318476 320719 318532 320728
rect 321696 320784 321752 320793
rect 321696 320719 321752 320728
rect 322432 320784 322488 320793
rect 322432 320719 322488 320728
rect 324088 320784 324144 320793
rect 324088 320719 324144 320728
rect 324640 320784 324696 320793
rect 324640 320719 324696 320728
rect 325192 320784 325248 320793
rect 325192 320719 325248 320728
rect 326480 320784 326536 320793
rect 326480 320719 326536 320728
rect 327400 320784 327456 320793
rect 327400 320719 327456 320728
rect 314798 320690 314850 320696
rect 284712 320648 284768 320657
rect 284712 320583 284768 320592
rect 285080 320648 285136 320657
rect 285080 320583 285136 320592
rect 288300 320648 288356 320657
rect 288300 320583 288356 320592
rect 292164 320648 292220 320657
rect 292164 320583 292220 320592
rect 293452 320648 293508 320657
rect 293452 320583 293508 320592
rect 294096 320648 294152 320657
rect 294096 320583 294152 320592
rect 298144 320648 298200 320657
rect 298144 320583 298200 320592
rect 298512 320648 298568 320657
rect 298512 320583 298568 320592
rect 299248 320648 299304 320657
rect 299248 320583 299304 320592
rect 304492 320648 304548 320657
rect 304492 320583 304548 320592
rect 305320 320648 305376 320657
rect 305320 320583 305376 320592
rect 307620 320648 307676 320657
rect 307620 320583 307622 320592
rect 307674 320583 307676 320592
rect 313784 320648 313840 320657
rect 313784 320583 313840 320592
rect 317832 320648 317888 320657
rect 317832 320583 317888 320592
rect 326756 320648 326812 320657
rect 326756 320583 326812 320592
rect 327308 320648 327364 320657
rect 327308 320583 327364 320592
rect 307622 320554 307674 320560
rect 299984 320512 300040 320521
rect 299984 320447 300040 320456
rect 300536 320512 300592 320521
rect 300536 320447 300592 320456
rect 302100 320512 302156 320521
rect 302100 320447 302156 320456
rect 305504 320512 305560 320521
rect 305504 320447 305560 320456
rect 312588 320512 312644 320521
rect 312588 320447 312644 320456
rect 313508 320512 313564 320521
rect 313508 320447 313564 320456
rect 319672 320512 319728 320521
rect 319672 320447 319728 320456
rect 322984 320512 323040 320521
rect 322984 320447 323040 320456
rect 324364 320512 324420 320521
rect 324364 320447 324420 320456
rect 325008 320512 325064 320521
rect 325008 320447 325064 320456
rect 308724 320376 308780 320385
rect 308724 320311 308780 320320
rect 309460 320376 309516 320385
rect 309460 320311 309516 320320
rect 310932 320376 310988 320385
rect 310932 320311 310988 320320
rect 311484 320376 311540 320385
rect 311484 320311 311540 320320
rect 323536 320376 323592 320385
rect 323536 320311 323592 320320
rect 325468 320376 325524 320385
rect 325468 320311 325524 320320
rect 326296 320376 326352 320385
rect 326296 320311 326352 320320
rect 284528 320240 284584 320249
rect 284528 320175 284584 320184
rect 284896 320240 284952 320249
rect 284896 320175 284952 320184
rect 285448 320240 285504 320249
rect 285448 320175 285504 320184
rect 286828 320240 286884 320249
rect 286828 320175 286884 320184
rect 287288 320240 287344 320249
rect 287288 320175 287344 320184
rect 288024 320240 288080 320249
rect 288024 320175 288080 320184
rect 290324 320240 290380 320249
rect 290324 320175 290380 320184
rect 291980 320240 292036 320249
rect 291980 320175 292036 320184
rect 292440 320240 292496 320249
rect 292440 320175 292496 320184
rect 293728 320240 293784 320249
rect 293728 320175 293784 320184
rect 294280 320240 294336 320249
rect 294280 320175 294336 320184
rect 294648 320240 294704 320249
rect 294648 320175 294704 320184
rect 295016 320240 295072 320249
rect 295016 320175 295072 320184
rect 296028 320240 296084 320249
rect 296028 320175 296084 320184
rect 296488 320240 296544 320249
rect 296488 320175 296544 320184
rect 296948 320240 297004 320249
rect 296948 320175 297004 320184
rect 298696 320240 298752 320249
rect 298696 320175 298752 320184
rect 299156 320240 299212 320249
rect 299156 320175 299212 320184
rect 300168 320240 300224 320249
rect 300168 320175 300224 320184
rect 302744 320240 302800 320249
rect 302744 320175 302800 320184
rect 305136 320240 305192 320249
rect 305136 320175 305192 320184
rect 306240 320240 306296 320249
rect 306240 320175 306296 320184
rect 307068 320240 307124 320249
rect 307068 320175 307124 320184
rect 308448 320240 308504 320249
rect 308448 320175 308504 320184
rect 308632 320240 308688 320249
rect 308632 320175 308688 320184
rect 309644 320240 309700 320249
rect 309644 320175 309700 320184
rect 312496 320240 312552 320249
rect 312496 320175 312552 320184
rect 314152 320240 314208 320249
rect 314152 320175 314208 320184
rect 314980 320240 315036 320249
rect 314980 320175 315036 320184
rect 316912 320240 316968 320249
rect 316912 320175 316968 320184
rect 319120 320240 319176 320249
rect 319120 320175 319176 320184
rect 319856 320240 319912 320249
rect 319856 320175 319912 320184
rect 320592 320240 320648 320249
rect 320592 320175 320648 320184
rect 282872 320104 282928 320113
rect 282518 319841 282546 320076
rect 282610 319870 282638 320076
rect 282794 319920 282822 320076
rect 283332 320104 283388 320113
rect 282872 320039 282928 320048
rect 282748 319892 282822 319920
rect 282598 319864 282650 319870
rect 282504 319832 282560 319841
rect 282598 319806 282650 319812
rect 282504 319767 282560 319776
rect 282748 318306 282776 319892
rect 282978 319852 283006 320076
rect 282932 319824 283006 319852
rect 282828 319796 282880 319802
rect 282828 319738 282880 319744
rect 282840 319530 282868 319738
rect 282828 319524 282880 319530
rect 282828 319466 282880 319472
rect 282932 319297 282960 319824
rect 283070 319784 283098 320076
rect 283162 319818 283190 320076
rect 283254 319920 283282 320076
rect 283608 320104 283664 320113
rect 283332 320039 283388 320048
rect 283254 319892 283328 319920
rect 283162 319790 283236 319818
rect 283024 319756 283098 319784
rect 282918 319288 282974 319297
rect 282918 319223 282974 319232
rect 282920 319184 282972 319190
rect 282920 319126 282972 319132
rect 282932 319054 282960 319126
rect 282920 319048 282972 319054
rect 282920 318990 282972 318996
rect 282736 318300 282788 318306
rect 282736 318242 282788 318248
rect 282642 317792 282698 317801
rect 282642 317727 282698 317736
rect 282366 316840 282422 316849
rect 282366 316775 282422 316784
rect 282276 291984 282328 291990
rect 282276 291926 282328 291932
rect 282276 241188 282328 241194
rect 282276 241130 282328 241136
rect 282184 216300 282236 216306
rect 282184 216242 282236 216248
rect 282184 146192 282236 146198
rect 282184 146134 282236 146140
rect 281540 140752 281592 140758
rect 281540 140694 281592 140700
rect 281552 140146 281580 140694
rect 281540 140140 281592 140146
rect 281540 140082 281592 140088
rect 280804 140072 280856 140078
rect 280804 140014 280856 140020
rect 280068 33108 280120 33114
rect 280068 33050 280120 33056
rect 278792 16546 279096 16574
rect 278320 4140 278372 4146
rect 278320 4082 278372 4088
rect 278044 3392 278096 3398
rect 277122 3360 277178 3369
rect 278044 3334 278096 3340
rect 277122 3295 277178 3304
rect 277136 480 277164 3295
rect 278332 480 278360 4082
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280710 6080 280766 6089
rect 280710 6015 280766 6024
rect 280724 480 280752 6015
rect 281908 3392 281960 3398
rect 281908 3334 281960 3340
rect 281920 480 281948 3334
rect 282196 3194 282224 146134
rect 282288 139398 282316 241130
rect 282380 227186 282408 316775
rect 282552 316056 282604 316062
rect 282552 315998 282604 316004
rect 282460 313948 282512 313954
rect 282460 313890 282512 313896
rect 282472 240281 282500 313890
rect 282458 240272 282514 240281
rect 282458 240207 282514 240216
rect 282460 235476 282512 235482
rect 282460 235418 282512 235424
rect 282368 227180 282420 227186
rect 282368 227122 282420 227128
rect 282472 149025 282500 235418
rect 282564 232490 282592 315998
rect 282656 304978 282684 317727
rect 282828 317620 282880 317626
rect 282828 317562 282880 317568
rect 282736 311228 282788 311234
rect 282736 311170 282788 311176
rect 282644 304972 282696 304978
rect 282644 304914 282696 304920
rect 282552 232484 282604 232490
rect 282552 232426 282604 232432
rect 282656 225418 282684 304914
rect 282748 234258 282776 311170
rect 282840 298110 282868 317562
rect 282828 298104 282880 298110
rect 282828 298046 282880 298052
rect 282840 297226 282868 298046
rect 282828 297220 282880 297226
rect 282828 297162 282880 297168
rect 282932 239222 282960 318990
rect 283024 317830 283052 319756
rect 283102 319696 283158 319705
rect 283102 319631 283158 319640
rect 283012 317824 283064 317830
rect 283012 317766 283064 317772
rect 283010 307728 283066 307737
rect 283010 307663 283066 307672
rect 282920 239216 282972 239222
rect 282920 239158 282972 239164
rect 282736 234252 282788 234258
rect 282736 234194 282788 234200
rect 283024 230353 283052 307663
rect 283116 304774 283144 319631
rect 283208 318306 283236 319790
rect 283300 319580 283328 319892
rect 283438 319784 283466 320076
rect 283392 319756 283466 319784
rect 283530 319784 283558 320076
rect 284068 320104 284124 320113
rect 283608 320039 283664 320048
rect 283530 319756 283604 319784
rect 283392 319648 283420 319756
rect 283392 319620 283512 319648
rect 283300 319552 283420 319580
rect 283288 319388 283340 319394
rect 283288 319330 283340 319336
rect 283196 318300 283248 318306
rect 283196 318242 283248 318248
rect 283196 318096 283248 318102
rect 283196 318038 283248 318044
rect 283208 307766 283236 318038
rect 283300 310418 283328 319330
rect 283392 318782 283420 319552
rect 283380 318776 283432 318782
rect 283380 318718 283432 318724
rect 283380 317416 283432 317422
rect 283380 317358 283432 317364
rect 283288 310412 283340 310418
rect 283288 310354 283340 310360
rect 283196 307760 283248 307766
rect 283196 307702 283248 307708
rect 283104 304768 283156 304774
rect 283104 304710 283156 304716
rect 283392 241369 283420 317358
rect 283484 315994 283512 319620
rect 283576 319530 283604 319756
rect 283714 319682 283742 320076
rect 283806 319943 283834 320076
rect 283792 319934 283848 319943
rect 283792 319869 283848 319878
rect 283898 319852 283926 320076
rect 285632 320104 285688 320113
rect 284068 320039 284124 320048
rect 283898 319824 283972 319852
rect 283714 319654 283788 319682
rect 283564 319524 283616 319530
rect 283564 319466 283616 319472
rect 283654 319424 283710 319433
rect 283564 319388 283616 319394
rect 283760 319394 283788 319654
rect 283654 319359 283710 319368
rect 283748 319388 283800 319394
rect 283564 319330 283616 319336
rect 283576 317529 283604 319330
rect 283668 318374 283696 319359
rect 283748 319330 283800 319336
rect 283748 319048 283800 319054
rect 283748 318990 283800 318996
rect 283838 319016 283894 319025
rect 283760 318850 283788 318990
rect 283838 318951 283894 318960
rect 283852 318850 283880 318951
rect 283748 318844 283800 318850
rect 283748 318786 283800 318792
rect 283840 318844 283892 318850
rect 283840 318786 283892 318792
rect 283656 318368 283708 318374
rect 283656 318310 283708 318316
rect 283562 317520 283618 317529
rect 283562 317455 283618 317464
rect 283472 315988 283524 315994
rect 283472 315930 283524 315936
rect 283852 315382 283880 318786
rect 283944 318102 283972 319824
rect 284174 319818 284202 320076
rect 284266 319943 284294 320076
rect 284252 319934 284308 319943
rect 284252 319869 284308 319878
rect 284450 319852 284478 320076
rect 284450 319824 284524 319852
rect 284174 319790 284248 319818
rect 284022 319696 284078 319705
rect 284022 319631 284078 319640
rect 284036 319433 284064 319631
rect 284022 319424 284078 319433
rect 284022 319359 284078 319368
rect 284036 318458 284064 319359
rect 284220 319190 284248 319790
rect 284298 319696 284354 319705
rect 284298 319631 284354 319640
rect 284208 319184 284260 319190
rect 284208 319126 284260 319132
rect 284312 318481 284340 319631
rect 284496 319444 284524 319824
rect 284634 319784 284662 320076
rect 284818 319954 284846 320076
rect 284818 319938 284892 319954
rect 284818 319932 284904 319938
rect 284818 319926 284852 319932
rect 284852 319874 284904 319880
rect 284852 319796 284904 319802
rect 284634 319756 284708 319784
rect 284404 319416 284524 319444
rect 284298 318472 284354 318481
rect 284036 318430 284156 318458
rect 284024 318300 284076 318306
rect 284024 318242 284076 318248
rect 283932 318096 283984 318102
rect 283932 318038 283984 318044
rect 283930 317928 283986 317937
rect 283930 317863 283986 317872
rect 283840 315376 283892 315382
rect 283840 315318 283892 315324
rect 283654 314664 283710 314673
rect 283654 314599 283710 314608
rect 283564 310412 283616 310418
rect 283564 310354 283616 310360
rect 283576 309534 283604 310354
rect 283564 309528 283616 309534
rect 283564 309470 283616 309476
rect 283576 296002 283604 309470
rect 283564 295996 283616 296002
rect 283564 295938 283616 295944
rect 283378 241360 283434 241369
rect 283378 241295 283434 241304
rect 283564 241256 283616 241262
rect 283564 241198 283616 241204
rect 283010 230344 283066 230353
rect 283010 230279 283066 230288
rect 282644 225412 282696 225418
rect 282644 225354 282696 225360
rect 282458 149016 282514 149025
rect 282458 148951 282514 148960
rect 282472 148345 282500 148951
rect 282458 148336 282514 148345
rect 282458 148271 282514 148280
rect 282920 143404 282972 143410
rect 282920 143346 282972 143352
rect 282932 142866 282960 143346
rect 282920 142860 282972 142866
rect 282920 142802 282972 142808
rect 282276 139392 282328 139398
rect 282276 139334 282328 139340
rect 282288 138786 282316 139334
rect 282276 138780 282328 138786
rect 282276 138722 282328 138728
rect 282920 137964 282972 137970
rect 282920 137906 282972 137912
rect 282932 137426 282960 137906
rect 283576 137426 283604 241198
rect 283668 216442 283696 314599
rect 283746 310584 283802 310593
rect 283746 310519 283802 310528
rect 283760 224194 283788 310519
rect 283840 307216 283892 307222
rect 283840 307158 283892 307164
rect 283748 224188 283800 224194
rect 283748 224130 283800 224136
rect 283852 221678 283880 307158
rect 283944 305833 283972 317863
rect 283930 305824 283986 305833
rect 283930 305759 283986 305768
rect 283930 299024 283986 299033
rect 283930 298959 283986 298968
rect 283840 221672 283892 221678
rect 283840 221614 283892 221620
rect 283748 220176 283800 220182
rect 283748 220118 283800 220124
rect 283656 216436 283708 216442
rect 283656 216378 283708 216384
rect 283760 142866 283788 220118
rect 283944 216374 283972 298959
rect 284036 295322 284064 318242
rect 284128 316713 284156 318430
rect 284298 318407 284354 318416
rect 284208 318368 284260 318374
rect 284208 318310 284260 318316
rect 284220 317422 284248 318310
rect 284208 317416 284260 317422
rect 284404 317393 284432 319416
rect 284482 319288 284538 319297
rect 284482 319223 284538 319232
rect 284208 317358 284260 317364
rect 284390 317384 284446 317393
rect 284390 317319 284446 317328
rect 284114 316704 284170 316713
rect 284114 316639 284170 316648
rect 284496 316146 284524 319223
rect 284680 317665 284708 319756
rect 285002 319784 285030 320076
rect 285186 319920 285214 320076
rect 284852 319738 284904 319744
rect 284956 319756 285030 319784
rect 285094 319892 285214 319920
rect 284760 319184 284812 319190
rect 284760 319126 284812 319132
rect 284772 319025 284800 319126
rect 284758 319016 284814 319025
rect 284758 318951 284814 318960
rect 284864 318782 284892 319738
rect 284852 318776 284904 318782
rect 284852 318718 284904 318724
rect 284852 317688 284904 317694
rect 284666 317656 284722 317665
rect 284852 317630 284904 317636
rect 284666 317591 284722 317600
rect 284496 316118 284616 316146
rect 284484 315988 284536 315994
rect 284484 315930 284536 315936
rect 284300 314492 284352 314498
rect 284300 314434 284352 314440
rect 284312 313614 284340 314434
rect 284300 313608 284352 313614
rect 284300 313550 284352 313556
rect 284116 304088 284168 304094
rect 284116 304030 284168 304036
rect 284024 295316 284076 295322
rect 284024 295258 284076 295264
rect 284036 295089 284064 295258
rect 284022 295080 284078 295089
rect 284022 295015 284078 295024
rect 284024 232552 284076 232558
rect 284024 232494 284076 232500
rect 283932 216368 283984 216374
rect 283932 216310 283984 216316
rect 284036 151745 284064 232494
rect 284128 225486 284156 304030
rect 284312 241097 284340 313550
rect 284496 310486 284524 315930
rect 284484 310480 284536 310486
rect 284484 310422 284536 310428
rect 284588 296750 284616 316118
rect 284864 316033 284892 317630
rect 284956 317529 284984 319756
rect 285094 319716 285122 319892
rect 285278 319818 285306 320076
rect 285370 319920 285398 320076
rect 286276 320104 286332 320113
rect 285632 320039 285688 320048
rect 285738 319920 285766 320076
rect 285370 319892 285444 319920
rect 285416 319818 285444 319892
rect 285692 319892 285766 319920
rect 285830 319920 285858 320076
rect 286014 319920 286042 320076
rect 286106 319938 286134 320076
rect 285830 319892 285904 319920
rect 285586 319832 285642 319841
rect 285278 319790 285352 319818
rect 285416 319790 285490 319818
rect 285094 319688 285168 319716
rect 285034 319016 285090 319025
rect 285034 318951 285090 318960
rect 285048 317694 285076 318951
rect 285140 317898 285168 319688
rect 285324 318866 285352 319790
rect 285462 319784 285490 319790
rect 285462 319756 285536 319784
rect 285586 319767 285642 319776
rect 285232 318838 285352 318866
rect 285128 317892 285180 317898
rect 285128 317834 285180 317840
rect 285036 317688 285088 317694
rect 285036 317630 285088 317636
rect 284942 317520 284998 317529
rect 285126 317520 285182 317529
rect 284942 317455 284998 317464
rect 285048 317478 285126 317506
rect 284850 316024 284906 316033
rect 284850 315959 284906 315968
rect 285048 311894 285076 317478
rect 285126 317455 285182 317464
rect 285128 315376 285180 315382
rect 285128 315318 285180 315324
rect 284956 311866 285076 311894
rect 284576 296744 284628 296750
rect 284576 296686 284628 296692
rect 284588 295186 284616 296686
rect 284576 295180 284628 295186
rect 284576 295122 284628 295128
rect 284852 242344 284904 242350
rect 284852 242286 284904 242292
rect 284298 241088 284354 241097
rect 284298 241023 284354 241032
rect 284484 237448 284536 237454
rect 284484 237390 284536 237396
rect 284300 234728 284352 234734
rect 284300 234670 284352 234676
rect 284116 225480 284168 225486
rect 284116 225422 284168 225428
rect 284022 151736 284078 151745
rect 284022 151671 284078 151680
rect 284036 151201 284064 151671
rect 284022 151192 284078 151201
rect 284022 151127 284078 151136
rect 283748 142860 283800 142866
rect 283748 142802 283800 142808
rect 282920 137420 282972 137426
rect 282920 137362 282972 137368
rect 283564 137420 283616 137426
rect 283564 137362 283616 137368
rect 284312 128314 284340 234670
rect 284392 231804 284444 231810
rect 284392 231746 284444 231752
rect 284404 231470 284432 231746
rect 284392 231464 284444 231470
rect 284392 231406 284444 231412
rect 284404 139330 284432 231406
rect 284496 151609 284524 237390
rect 284864 235822 284892 242286
rect 284852 235816 284904 235822
rect 284852 235758 284904 235764
rect 284864 234734 284892 235758
rect 284852 234728 284904 234734
rect 284852 234670 284904 234676
rect 284956 217841 284984 311866
rect 285036 311160 285088 311166
rect 285036 311102 285088 311108
rect 285048 225554 285076 311102
rect 285140 231810 285168 315318
rect 285232 314498 285260 318838
rect 285312 318164 285364 318170
rect 285312 318106 285364 318112
rect 285220 314492 285272 314498
rect 285220 314434 285272 314440
rect 285220 307352 285272 307358
rect 285220 307294 285272 307300
rect 285128 231804 285180 231810
rect 285128 231746 285180 231752
rect 285036 225548 285088 225554
rect 285036 225490 285088 225496
rect 285232 224466 285260 307294
rect 285324 239426 285352 318106
rect 285404 317484 285456 317490
rect 285404 317426 285456 317432
rect 285416 315858 285444 317426
rect 285404 315852 285456 315858
rect 285404 315794 285456 315800
rect 285508 307290 285536 319756
rect 285600 315994 285628 319767
rect 285692 316130 285720 319892
rect 285770 319832 285826 319841
rect 285770 319767 285826 319776
rect 285784 318714 285812 319767
rect 285772 318708 285824 318714
rect 285772 318650 285824 318656
rect 285876 318646 285904 319892
rect 285968 319892 286042 319920
rect 286094 319932 286146 319938
rect 285968 319274 285996 319892
rect 286094 319874 286146 319880
rect 286198 319841 286226 320076
rect 286920 320104 286976 320113
rect 286276 320039 286332 320048
rect 286184 319832 286240 319841
rect 286184 319767 286240 319776
rect 286290 319682 286318 320039
rect 286382 319784 286410 320076
rect 286474 319943 286502 320076
rect 286460 319934 286516 319943
rect 286460 319869 286516 319878
rect 286566 319784 286594 320076
rect 286382 319756 286456 319784
rect 286244 319654 286318 319682
rect 285968 319246 286088 319274
rect 285864 318640 285916 318646
rect 285864 318582 285916 318588
rect 285864 318300 285916 318306
rect 285864 318242 285916 318248
rect 285680 316124 285732 316130
rect 285680 316066 285732 316072
rect 285588 315988 285640 315994
rect 285588 315930 285640 315936
rect 285588 315852 285640 315858
rect 285588 315794 285640 315800
rect 285496 307284 285548 307290
rect 285496 307226 285548 307232
rect 285402 297120 285458 297129
rect 285402 297055 285458 297064
rect 285312 239420 285364 239426
rect 285312 239362 285364 239368
rect 285220 224460 285272 224466
rect 285220 224402 285272 224408
rect 285416 222737 285444 297055
rect 285508 242729 285536 307226
rect 285600 298994 285628 315794
rect 285678 309360 285734 309369
rect 285678 309295 285734 309304
rect 285692 309262 285720 309295
rect 285680 309256 285732 309262
rect 285680 309198 285732 309204
rect 285876 306066 285904 318242
rect 286060 317694 286088 319246
rect 286244 318345 286272 319654
rect 286230 318336 286286 318345
rect 286230 318271 286286 318280
rect 286048 317688 286100 317694
rect 286048 317630 286100 317636
rect 286230 317656 286286 317665
rect 285956 315988 286008 315994
rect 285956 315930 286008 315936
rect 285968 309126 285996 315930
rect 286060 313478 286088 317630
rect 286230 317591 286286 317600
rect 286140 316124 286192 316130
rect 286140 316066 286192 316072
rect 286048 313472 286100 313478
rect 286048 313414 286100 313420
rect 286152 310185 286180 316066
rect 286138 310176 286194 310185
rect 286138 310111 286194 310120
rect 285956 309120 286008 309126
rect 285956 309062 286008 309068
rect 285864 306060 285916 306066
rect 285864 306002 285916 306008
rect 285876 304366 285904 306002
rect 285864 304360 285916 304366
rect 285864 304302 285916 304308
rect 285588 298988 285640 298994
rect 285588 298930 285640 298936
rect 285494 242720 285550 242729
rect 285494 242655 285550 242664
rect 285600 241233 285628 298930
rect 285864 244928 285916 244934
rect 285864 244870 285916 244876
rect 285586 241224 285642 241233
rect 285586 241159 285642 241168
rect 285876 237046 285904 244870
rect 286244 242865 286272 317591
rect 286428 306338 286456 319756
rect 286520 319756 286594 319784
rect 286520 318753 286548 319756
rect 286658 319716 286686 320076
rect 286750 319784 286778 320076
rect 287196 320104 287252 320113
rect 286920 320039 286976 320048
rect 287026 319954 287054 320076
rect 286980 319926 287054 319954
rect 286750 319756 286916 319784
rect 286658 319688 286732 319716
rect 286600 319592 286652 319598
rect 286600 319534 286652 319540
rect 286506 318744 286562 318753
rect 286506 318679 286562 318688
rect 286520 317665 286548 318679
rect 286612 318578 286640 319534
rect 286600 318572 286652 318578
rect 286600 318514 286652 318520
rect 286704 318306 286732 319688
rect 286782 319696 286838 319705
rect 286782 319631 286838 319640
rect 286692 318300 286744 318306
rect 286692 318242 286744 318248
rect 286600 318096 286652 318102
rect 286600 318038 286652 318044
rect 286692 318096 286744 318102
rect 286692 318038 286744 318044
rect 286612 317898 286640 318038
rect 286600 317892 286652 317898
rect 286600 317834 286652 317840
rect 286506 317656 286562 317665
rect 286506 317591 286562 317600
rect 286704 311894 286732 318038
rect 286612 311866 286732 311894
rect 286508 310072 286560 310078
rect 286508 310014 286560 310020
rect 286416 306332 286468 306338
rect 286416 306274 286468 306280
rect 286324 305856 286376 305862
rect 286324 305798 286376 305804
rect 286230 242856 286286 242865
rect 286230 242791 286286 242800
rect 285864 237040 285916 237046
rect 285864 236982 285916 236988
rect 285680 235544 285732 235550
rect 285680 235486 285732 235492
rect 285692 234394 285720 235486
rect 285680 234388 285732 234394
rect 285680 234330 285732 234336
rect 285402 222728 285458 222737
rect 285402 222663 285458 222672
rect 284942 217832 284998 217841
rect 284942 217767 284998 217776
rect 284482 151600 284538 151609
rect 284482 151535 284538 151544
rect 284496 151065 284524 151535
rect 284482 151056 284538 151065
rect 284482 150991 284538 151000
rect 284944 144832 284996 144838
rect 284944 144774 284996 144780
rect 284392 139324 284444 139330
rect 284392 139266 284444 139272
rect 284404 138718 284432 139266
rect 284392 138712 284444 138718
rect 284392 138654 284444 138660
rect 284300 128308 284352 128314
rect 284300 128250 284352 128256
rect 284312 127702 284340 128250
rect 284300 127696 284352 127702
rect 284300 127638 284352 127644
rect 284298 6896 284354 6905
rect 284298 6831 284354 6840
rect 283104 3800 283156 3806
rect 283104 3742 283156 3748
rect 282184 3188 282236 3194
rect 282184 3130 282236 3136
rect 283116 480 283144 3742
rect 284312 480 284340 6831
rect 284956 3738 284984 144774
rect 285692 16574 285720 234330
rect 285772 226908 285824 226914
rect 285772 226850 285824 226856
rect 285784 226710 285812 226850
rect 285772 226704 285824 226710
rect 285772 226646 285824 226652
rect 285784 125594 285812 226646
rect 285876 142118 285904 236982
rect 286336 221542 286364 305798
rect 286414 298072 286470 298081
rect 286414 298007 286470 298016
rect 286428 296993 286456 298007
rect 286414 296984 286470 296993
rect 286414 296919 286470 296928
rect 286324 221536 286376 221542
rect 286324 221478 286376 221484
rect 286428 216510 286456 296919
rect 286520 228274 286548 310014
rect 286612 237182 286640 311866
rect 286692 304564 286744 304570
rect 286692 304506 286744 304512
rect 286600 237176 286652 237182
rect 286600 237118 286652 237124
rect 286508 228268 286560 228274
rect 286508 228210 286560 228216
rect 286704 224126 286732 304506
rect 286796 298081 286824 319631
rect 286888 317490 286916 319756
rect 286876 317484 286928 317490
rect 286876 317426 286928 317432
rect 286980 315994 287008 319926
rect 287118 319920 287146 320076
rect 287472 320104 287528 320113
rect 287196 320039 287252 320048
rect 287118 319892 287192 319920
rect 287058 319288 287114 319297
rect 287058 319223 287114 319232
rect 287072 318986 287100 319223
rect 287060 318980 287112 318986
rect 287060 318922 287112 318928
rect 287060 318776 287112 318782
rect 287060 318718 287112 318724
rect 286968 315988 287020 315994
rect 286968 315930 287020 315936
rect 287072 313274 287100 318718
rect 287164 317422 287192 319892
rect 287242 319832 287298 319841
rect 287394 319784 287422 320076
rect 287840 320104 287896 320113
rect 287472 320039 287528 320048
rect 287578 319852 287606 320076
rect 287242 319767 287298 319776
rect 287256 319161 287284 319767
rect 287348 319756 287422 319784
rect 287532 319824 287606 319852
rect 287242 319152 287298 319161
rect 287242 319087 287298 319096
rect 287242 319016 287298 319025
rect 287242 318951 287298 318960
rect 287256 318782 287284 318951
rect 287244 318776 287296 318782
rect 287244 318718 287296 318724
rect 287348 318073 287376 319756
rect 287426 319696 287482 319705
rect 287426 319631 287482 319640
rect 287334 318064 287390 318073
rect 287334 317999 287390 318008
rect 287336 317688 287388 317694
rect 287334 317656 287336 317665
rect 287388 317656 287390 317665
rect 287334 317591 287390 317600
rect 287152 317416 287204 317422
rect 287152 317358 287204 317364
rect 287152 315988 287204 315994
rect 287152 315930 287204 315936
rect 287060 313268 287112 313274
rect 287060 313210 287112 313216
rect 286876 310004 286928 310010
rect 286876 309946 286928 309952
rect 286782 298072 286838 298081
rect 286782 298007 286838 298016
rect 286782 297664 286838 297673
rect 286782 297599 286838 297608
rect 286692 224120 286744 224126
rect 286692 224062 286744 224068
rect 286796 221921 286824 297599
rect 286888 234462 286916 309946
rect 287164 298042 287192 315930
rect 287244 315852 287296 315858
rect 287244 315794 287296 315800
rect 287256 311846 287284 315794
rect 287336 314900 287388 314906
rect 287336 314842 287388 314848
rect 287244 311840 287296 311846
rect 287244 311782 287296 311788
rect 287348 302161 287376 314842
rect 287440 311778 287468 319631
rect 287428 311772 287480 311778
rect 287428 311714 287480 311720
rect 287334 302152 287390 302161
rect 287334 302087 287390 302096
rect 287532 301578 287560 319824
rect 287670 319818 287698 320076
rect 287762 319920 287790 320076
rect 288116 320104 288172 320113
rect 287840 320039 287896 320048
rect 287762 319892 287836 319920
rect 287670 319790 287744 319818
rect 287610 319696 287666 319705
rect 287610 319631 287666 319640
rect 287624 319598 287652 319631
rect 287612 319592 287664 319598
rect 287612 319534 287664 319540
rect 287612 319456 287664 319462
rect 287612 319398 287664 319404
rect 287624 318714 287652 319398
rect 287716 318782 287744 319790
rect 287704 318776 287756 318782
rect 287704 318718 287756 318724
rect 287612 318708 287664 318714
rect 287612 318650 287664 318656
rect 287704 318572 287756 318578
rect 287704 318514 287756 318520
rect 287610 318064 287666 318073
rect 287716 318034 287744 318514
rect 287610 317999 287666 318008
rect 287704 318028 287756 318034
rect 287520 301572 287572 301578
rect 287520 301514 287572 301520
rect 287152 298036 287204 298042
rect 287152 297978 287204 297984
rect 287624 296041 287652 317999
rect 287704 317970 287756 317976
rect 287808 315994 287836 319892
rect 287946 319841 287974 320076
rect 288484 320104 288540 320113
rect 288116 320039 288172 320048
rect 288222 319954 288250 320076
rect 288668 320104 288724 320113
rect 288484 320039 288540 320048
rect 288590 319954 288618 320076
rect 289220 320104 289276 320113
rect 288668 320039 288724 320048
rect 288222 319926 288296 319954
rect 287932 319832 287988 319841
rect 287932 319767 287988 319776
rect 288268 319784 288296 319926
rect 288452 319926 288618 319954
rect 288268 319756 288342 319784
rect 287978 319696 288034 319705
rect 287978 319631 288034 319640
rect 287888 318776 287940 318782
rect 287888 318718 287940 318724
rect 287796 315988 287848 315994
rect 287796 315930 287848 315936
rect 287702 313848 287758 313857
rect 287702 313783 287758 313792
rect 287716 313410 287744 313783
rect 287704 313404 287756 313410
rect 287704 313346 287756 313352
rect 287796 311500 287848 311506
rect 287796 311442 287848 311448
rect 287704 307692 287756 307698
rect 287704 307634 287756 307640
rect 287610 296032 287666 296041
rect 287610 295967 287666 295976
rect 287612 244996 287664 245002
rect 287612 244938 287664 244944
rect 286968 239556 287020 239562
rect 286968 239498 287020 239504
rect 286876 234456 286928 234462
rect 286876 234398 286928 234404
rect 286980 226710 287008 239498
rect 287518 233880 287574 233889
rect 287518 233815 287574 233824
rect 287152 232688 287204 232694
rect 287152 232630 287204 232636
rect 286968 226704 287020 226710
rect 286968 226646 287020 226652
rect 286782 221912 286838 221921
rect 286782 221847 286838 221856
rect 286416 216504 286468 216510
rect 286416 216446 286468 216452
rect 287060 168428 287112 168434
rect 287060 168370 287112 168376
rect 285864 142112 285916 142118
rect 285864 142054 285916 142060
rect 285876 140826 285904 142054
rect 285864 140820 285916 140826
rect 285864 140762 285916 140768
rect 286324 140820 286376 140826
rect 286324 140762 286376 140768
rect 286336 130422 286364 140762
rect 286324 130416 286376 130422
rect 286324 130358 286376 130364
rect 285772 125588 285824 125594
rect 285772 125530 285824 125536
rect 286232 125588 286284 125594
rect 286232 125530 286284 125536
rect 286244 124914 286272 125530
rect 286232 124908 286284 124914
rect 286232 124850 286284 124856
rect 287072 16574 287100 168370
rect 287164 132462 287192 232630
rect 287532 227322 287560 233815
rect 287624 232694 287652 244938
rect 287716 236910 287744 307634
rect 287704 236904 287756 236910
rect 287704 236846 287756 236852
rect 287612 232688 287664 232694
rect 287612 232630 287664 232636
rect 287808 229974 287836 311442
rect 287900 309641 287928 318718
rect 287992 317937 288020 319631
rect 288314 319580 288342 319756
rect 288176 319552 288342 319580
rect 288070 319288 288126 319297
rect 288070 319223 288126 319232
rect 287978 317928 288034 317937
rect 287978 317863 288034 317872
rect 287980 311364 288032 311370
rect 287980 311306 288032 311312
rect 287886 309632 287942 309641
rect 287886 309567 287942 309576
rect 287888 301572 287940 301578
rect 287888 301514 287940 301520
rect 287796 229968 287848 229974
rect 287702 229936 287758 229945
rect 287796 229910 287848 229916
rect 287702 229871 287758 229880
rect 287520 227316 287572 227322
rect 287520 227258 287572 227264
rect 287532 226370 287560 227258
rect 287520 226364 287572 226370
rect 287520 226306 287572 226312
rect 287244 154148 287296 154154
rect 287244 154090 287296 154096
rect 287256 147558 287284 154090
rect 287244 147552 287296 147558
rect 287244 147494 287296 147500
rect 287716 142154 287744 229871
rect 287796 226364 287848 226370
rect 287796 226306 287848 226312
rect 287532 142126 287744 142154
rect 287532 142050 287560 142126
rect 287520 142044 287572 142050
rect 287520 141986 287572 141992
rect 287532 141574 287560 141986
rect 287808 141982 287836 226306
rect 287900 217394 287928 301514
rect 287992 230042 288020 311306
rect 288084 309058 288112 319223
rect 288176 314906 288204 319552
rect 288256 319456 288308 319462
rect 288256 319398 288308 319404
rect 288268 315858 288296 319398
rect 288348 318980 288400 318986
rect 288348 318922 288400 318928
rect 288360 318753 288388 318922
rect 288346 318744 288402 318753
rect 288346 318679 288402 318688
rect 288452 318442 288480 319926
rect 288774 319920 288802 320076
rect 288728 319892 288802 319920
rect 288622 319832 288678 319841
rect 288622 319767 288678 319776
rect 288530 319696 288586 319705
rect 288530 319631 288586 319640
rect 288544 319462 288572 319631
rect 288532 319456 288584 319462
rect 288532 319398 288584 319404
rect 288532 318980 288584 318986
rect 288532 318922 288584 318928
rect 288440 318436 288492 318442
rect 288440 318378 288492 318384
rect 288440 318300 288492 318306
rect 288440 318242 288492 318248
rect 288348 317416 288400 317422
rect 288348 317358 288400 317364
rect 288256 315852 288308 315858
rect 288256 315794 288308 315800
rect 288164 314900 288216 314906
rect 288164 314842 288216 314848
rect 288254 309496 288310 309505
rect 288254 309431 288310 309440
rect 288268 309194 288296 309431
rect 288256 309188 288308 309194
rect 288256 309130 288308 309136
rect 288072 309052 288124 309058
rect 288072 308994 288124 309000
rect 288164 305040 288216 305046
rect 288164 304982 288216 304988
rect 288070 298208 288126 298217
rect 288070 298143 288126 298152
rect 287980 230036 288032 230042
rect 287980 229978 288032 229984
rect 288084 219094 288112 298143
rect 288176 228342 288204 304982
rect 288256 303068 288308 303074
rect 288256 303010 288308 303016
rect 288268 230110 288296 303010
rect 288360 296614 288388 317358
rect 288452 317121 288480 318242
rect 288438 317112 288494 317121
rect 288438 317047 288494 317056
rect 288544 316962 288572 318922
rect 288452 316934 288572 316962
rect 288348 296608 288400 296614
rect 288348 296550 288400 296556
rect 288360 296313 288388 296550
rect 288346 296304 288402 296313
rect 288346 296239 288402 296248
rect 288346 236600 288402 236609
rect 288346 236535 288402 236544
rect 288360 235958 288388 236535
rect 288348 235952 288400 235958
rect 288348 235894 288400 235900
rect 288256 230104 288308 230110
rect 288256 230046 288308 230052
rect 288164 228336 288216 228342
rect 288164 228278 288216 228284
rect 288072 219088 288124 219094
rect 288072 219030 288124 219036
rect 287888 217388 287940 217394
rect 287888 217330 287940 217336
rect 288360 154154 288388 235894
rect 288452 217977 288480 316934
rect 288532 315920 288584 315926
rect 288532 315862 288584 315868
rect 288544 306374 288572 315862
rect 288636 315858 288664 319767
rect 288624 315852 288676 315858
rect 288624 315794 288676 315800
rect 288544 306346 288664 306374
rect 288636 295254 288664 306346
rect 288728 296682 288756 319892
rect 288866 319852 288894 320076
rect 288958 319943 288986 320076
rect 288944 319934 289000 319943
rect 288944 319869 289000 319878
rect 288820 319824 288894 319852
rect 288820 317626 288848 319824
rect 289050 319818 289078 320076
rect 289772 320104 289828 320113
rect 289220 320039 289276 320048
rect 289268 319864 289320 319870
rect 289004 319790 289078 319818
rect 289174 319832 289230 319841
rect 289004 319784 289032 319790
rect 288958 319756 289032 319784
rect 289418 319852 289446 320076
rect 289268 319806 289320 319812
rect 289372 319824 289446 319852
rect 289174 319767 289230 319776
rect 288958 319682 288986 319756
rect 288958 319654 289032 319682
rect 288898 319288 288954 319297
rect 288898 319223 288954 319232
rect 288808 317620 288860 317626
rect 288808 317562 288860 317568
rect 288808 315988 288860 315994
rect 288808 315930 288860 315936
rect 288820 298897 288848 315930
rect 288912 315926 288940 319223
rect 289004 318730 289032 319654
rect 289084 319592 289136 319598
rect 289084 319534 289136 319540
rect 289096 319297 289124 319534
rect 289082 319288 289138 319297
rect 289082 319223 289138 319232
rect 289004 318702 289124 318730
rect 289096 318617 289124 318702
rect 289082 318608 289138 318617
rect 289082 318543 289138 318552
rect 288900 315920 288952 315926
rect 288900 315862 288952 315868
rect 288992 315920 289044 315926
rect 288992 315862 289044 315868
rect 288900 311296 288952 311302
rect 288900 311238 288952 311244
rect 288806 298888 288862 298897
rect 288806 298823 288862 298832
rect 288716 296676 288768 296682
rect 288716 296618 288768 296624
rect 288728 296177 288756 296618
rect 288714 296168 288770 296177
rect 288714 296103 288770 296112
rect 288624 295248 288676 295254
rect 288624 295190 288676 295196
rect 288636 294953 288664 295190
rect 288622 294944 288678 294953
rect 288622 294879 288678 294888
rect 288532 243772 288584 243778
rect 288532 243714 288584 243720
rect 288544 239057 288572 243714
rect 288912 243710 288940 311238
rect 289004 304910 289032 315862
rect 289096 311302 289124 318543
rect 289188 317937 289216 319767
rect 289280 319462 289308 319806
rect 289268 319456 289320 319462
rect 289268 319398 289320 319404
rect 289174 317928 289230 317937
rect 289174 317863 289230 317872
rect 289372 315994 289400 319824
rect 289510 319784 289538 320076
rect 289464 319756 289538 319784
rect 289464 318986 289492 319756
rect 289602 319546 289630 320076
rect 289694 319784 289722 320076
rect 290416 320104 290472 320113
rect 289772 320039 289828 320048
rect 289970 319938 289998 320076
rect 289958 319932 290010 319938
rect 289958 319874 290010 319880
rect 289818 319832 289874 319841
rect 289694 319756 289768 319784
rect 289818 319767 289874 319776
rect 290062 319784 290090 320076
rect 290154 319938 290182 320076
rect 290692 320104 290748 320113
rect 290416 320039 290472 320048
rect 290142 319932 290194 319938
rect 290142 319874 290194 319880
rect 290280 319932 290332 319938
rect 290280 319874 290332 319880
rect 290188 319796 290240 319802
rect 289556 319518 289630 319546
rect 289452 318980 289504 318986
rect 289452 318922 289504 318928
rect 289452 318844 289504 318850
rect 289452 318786 289504 318792
rect 289464 318034 289492 318786
rect 289556 318209 289584 319518
rect 289740 319444 289768 319756
rect 289648 319416 289768 319444
rect 289542 318200 289598 318209
rect 289542 318135 289598 318144
rect 289452 318028 289504 318034
rect 289452 317970 289504 317976
rect 289360 315988 289412 315994
rect 289360 315930 289412 315936
rect 289648 315926 289676 319416
rect 289726 319016 289782 319025
rect 289726 318951 289782 318960
rect 289636 315920 289688 315926
rect 289636 315862 289688 315868
rect 289360 315852 289412 315858
rect 289360 315794 289412 315800
rect 289176 311432 289228 311438
rect 289176 311374 289228 311380
rect 289084 311296 289136 311302
rect 289084 311238 289136 311244
rect 288992 304904 289044 304910
rect 288992 304846 289044 304852
rect 289084 300144 289136 300150
rect 289084 300086 289136 300092
rect 288900 243704 288952 243710
rect 288900 243646 288952 243652
rect 288530 239048 288586 239057
rect 288530 238983 288586 238992
rect 288438 217968 288494 217977
rect 288438 217903 288494 217912
rect 288348 154148 288400 154154
rect 288348 154090 288400 154096
rect 288360 153270 288388 154090
rect 288348 153264 288400 153270
rect 288348 153206 288400 153212
rect 288544 143546 288572 238983
rect 289096 235006 289124 300086
rect 289084 235000 289136 235006
rect 289084 234942 289136 234948
rect 288532 143540 288584 143546
rect 288532 143482 288584 143488
rect 287796 141976 287848 141982
rect 287796 141918 287848 141924
rect 287520 141568 287572 141574
rect 287520 141510 287572 141516
rect 287808 134638 287836 141918
rect 288544 137358 288572 143482
rect 288532 137352 288584 137358
rect 288532 137294 288584 137300
rect 287796 134632 287848 134638
rect 287796 134574 287848 134580
rect 287152 132456 287204 132462
rect 287152 132398 287204 132404
rect 288348 132456 288400 132462
rect 288348 132398 288400 132404
rect 287704 131844 287756 131850
rect 287704 131786 287756 131792
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 284944 3732 284996 3738
rect 284944 3674 284996 3680
rect 285404 3188 285456 3194
rect 285404 3130 285456 3136
rect 285416 480 285444 3130
rect 286612 480 286640 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 3670 287744 131786
rect 288360 131782 288388 132398
rect 288348 131776 288400 131782
rect 288348 131718 288400 131724
rect 287704 3664 287756 3670
rect 287704 3606 287756 3612
rect 289096 3534 289124 234942
rect 289188 227390 289216 311374
rect 289372 310457 289400 315794
rect 289358 310448 289414 310457
rect 289358 310383 289414 310392
rect 289360 302116 289412 302122
rect 289360 302058 289412 302064
rect 289176 227384 289228 227390
rect 289176 227326 289228 227332
rect 289268 226976 289320 226982
rect 289268 226918 289320 226924
rect 289176 156664 289228 156670
rect 289176 156606 289228 156612
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289084 3528 289136 3534
rect 289084 3470 289136 3476
rect 289004 480 289032 3470
rect 289188 3058 289216 156606
rect 289280 144906 289308 226918
rect 289372 223009 289400 302058
rect 289450 297256 289506 297265
rect 289450 297191 289506 297200
rect 289358 223000 289414 223009
rect 289358 222935 289414 222944
rect 289464 221785 289492 297191
rect 289740 294681 289768 318951
rect 289832 318794 289860 319767
rect 290062 319756 290136 319784
rect 290004 319524 290056 319530
rect 290004 319466 290056 319472
rect 289832 318766 289952 318794
rect 289818 318336 289874 318345
rect 289818 318271 289874 318280
rect 289832 317966 289860 318271
rect 289820 317960 289872 317966
rect 289820 317902 289872 317908
rect 289924 294817 289952 318766
rect 290016 299033 290044 319466
rect 290108 305590 290136 319756
rect 290188 319738 290240 319744
rect 290200 318850 290228 319738
rect 290188 318844 290240 318850
rect 290188 318786 290240 318792
rect 290200 311273 290228 318786
rect 290292 317830 290320 319874
rect 290522 319784 290550 320076
rect 290614 319841 290642 320076
rect 290968 320104 291024 320113
rect 290692 320039 290748 320048
rect 290706 319870 290734 320039
rect 290798 319870 290826 320076
rect 290890 319938 290918 320076
rect 291152 320104 291208 320113
rect 290968 320039 291024 320048
rect 290878 319932 290930 319938
rect 291074 319920 291102 320076
rect 291704 320104 291760 320113
rect 291152 320039 291208 320048
rect 291166 319938 291194 320039
rect 290878 319874 290930 319880
rect 291028 319892 291102 319920
rect 291154 319932 291206 319938
rect 290694 319864 290746 319870
rect 290476 319756 290550 319784
rect 290600 319832 290656 319841
rect 290694 319806 290746 319812
rect 290786 319864 290838 319870
rect 290786 319806 290838 319812
rect 290600 319767 290656 319776
rect 290370 319696 290426 319705
rect 290370 319631 290426 319640
rect 290384 318782 290412 319631
rect 290372 318776 290424 318782
rect 290372 318718 290424 318724
rect 290280 317824 290332 317830
rect 290280 317766 290332 317772
rect 290292 317490 290320 317766
rect 290280 317484 290332 317490
rect 290280 317426 290332 317432
rect 290186 311264 290242 311273
rect 290186 311199 290242 311208
rect 290096 305584 290148 305590
rect 290096 305526 290148 305532
rect 290002 299024 290058 299033
rect 290002 298959 290058 298968
rect 289910 294808 289966 294817
rect 289910 294743 289966 294752
rect 289726 294672 289782 294681
rect 289726 294607 289782 294616
rect 290384 254590 290412 318718
rect 290476 318374 290504 319756
rect 290738 319696 290794 319705
rect 290738 319631 290794 319640
rect 290556 319592 290608 319598
rect 290556 319534 290608 319540
rect 290464 318368 290516 318374
rect 290464 318310 290516 318316
rect 290568 318073 290596 319534
rect 290752 318560 290780 319631
rect 290752 318532 290964 318560
rect 290740 318436 290792 318442
rect 290740 318378 290792 318384
rect 290554 318064 290610 318073
rect 290554 317999 290610 318008
rect 290464 317484 290516 317490
rect 290464 317426 290516 317432
rect 290476 311250 290504 317426
rect 290476 311222 290596 311250
rect 290462 310448 290518 310457
rect 290462 310383 290518 310392
rect 290372 254584 290424 254590
rect 290372 254526 290424 254532
rect 289450 221776 289506 221785
rect 289450 221711 289506 221720
rect 290476 219230 290504 310383
rect 290568 306374 290596 311222
rect 290568 306346 290688 306374
rect 290554 294808 290610 294817
rect 290554 294743 290610 294752
rect 290464 219224 290516 219230
rect 290464 219166 290516 219172
rect 290568 216345 290596 294743
rect 290660 251870 290688 306346
rect 290752 295089 290780 318378
rect 290936 318374 290964 318532
rect 291028 318442 291056 319892
rect 291154 319874 291206 319880
rect 291106 319832 291162 319841
rect 291258 319818 291286 320076
rect 291350 319920 291378 320076
rect 291350 319892 291424 319920
rect 291396 319818 291424 319892
rect 291534 319818 291562 320076
rect 291626 319954 291654 320076
rect 292808 320104 292864 320113
rect 291704 320039 291760 320048
rect 291626 319926 291700 319954
rect 291258 319790 291332 319818
rect 291396 319790 291470 319818
rect 291534 319790 291608 319818
rect 291106 319767 291162 319776
rect 291016 318436 291068 318442
rect 291016 318378 291068 318384
rect 290924 318368 290976 318374
rect 290924 318310 290976 318316
rect 290936 318152 290964 318310
rect 290936 318124 291056 318152
rect 290922 318064 290978 318073
rect 290922 317999 290978 318008
rect 290936 311894 290964 317999
rect 290844 311866 290964 311894
rect 290844 307426 290872 311866
rect 290832 307420 290884 307426
rect 290832 307362 290884 307368
rect 291028 306374 291056 318124
rect 291120 311409 291148 319767
rect 291200 319660 291252 319666
rect 291200 319602 291252 319608
rect 291212 319394 291240 319602
rect 291200 319388 291252 319394
rect 291200 319330 291252 319336
rect 291304 317150 291332 319790
rect 291442 319716 291470 319790
rect 291442 319688 291516 319716
rect 291384 319524 291436 319530
rect 291384 319466 291436 319472
rect 291396 318646 291424 319466
rect 291384 318640 291436 318646
rect 291384 318582 291436 318588
rect 291488 318238 291516 319688
rect 291580 319598 291608 319790
rect 291568 319592 291620 319598
rect 291568 319534 291620 319540
rect 291568 319388 291620 319394
rect 291568 319330 291620 319336
rect 291476 318232 291528 318238
rect 291476 318174 291528 318180
rect 291292 317144 291344 317150
rect 291292 317086 291344 317092
rect 291384 315988 291436 315994
rect 291384 315930 291436 315936
rect 291106 311400 291162 311409
rect 291106 311335 291162 311344
rect 291106 311264 291162 311273
rect 291106 311199 291162 311208
rect 291120 310554 291148 311199
rect 291108 310548 291160 310554
rect 291108 310490 291160 310496
rect 291108 307556 291160 307562
rect 291108 307498 291160 307504
rect 291120 307426 291148 307498
rect 291108 307420 291160 307426
rect 291108 307362 291160 307368
rect 290936 306346 291056 306374
rect 290738 295080 290794 295089
rect 290738 295015 290794 295024
rect 290648 251864 290700 251870
rect 290648 251806 290700 251812
rect 290646 229800 290702 229809
rect 290646 229735 290702 229744
rect 290554 216336 290610 216345
rect 290554 216271 290610 216280
rect 290660 157321 290688 229735
rect 290752 216481 290780 295015
rect 290936 283626 290964 306346
rect 291016 305584 291068 305590
rect 291016 305526 291068 305532
rect 291028 294545 291056 305526
rect 291396 304842 291424 315930
rect 291580 311894 291608 319330
rect 291672 315178 291700 319926
rect 291810 319920 291838 320076
rect 291902 319954 291930 320076
rect 291902 319926 291976 319954
rect 291764 319892 291838 319920
rect 291764 319025 291792 319892
rect 291844 319796 291896 319802
rect 291844 319738 291896 319744
rect 291750 319016 291806 319025
rect 291750 318951 291806 318960
rect 291856 318794 291884 319738
rect 291948 319716 291976 319926
rect 292086 319818 292114 320076
rect 292166 319932 292218 319938
rect 292270 319920 292298 320076
rect 292362 319954 292390 320076
rect 292362 319926 292436 319954
rect 292218 319892 292298 319920
rect 292166 319874 292218 319880
rect 292302 319832 292358 319841
rect 292086 319790 292252 319818
rect 291948 319688 292068 319716
rect 291936 319592 291988 319598
rect 291936 319534 291988 319540
rect 291764 318766 291884 318794
rect 291660 315172 291712 315178
rect 291660 315114 291712 315120
rect 291488 311866 291608 311894
rect 291488 305794 291516 311866
rect 291476 305788 291528 305794
rect 291476 305730 291528 305736
rect 291488 305046 291516 305730
rect 291476 305040 291528 305046
rect 291476 304982 291528 304988
rect 291384 304836 291436 304842
rect 291384 304778 291436 304784
rect 291764 303006 291792 318766
rect 291844 318708 291896 318714
rect 291844 318650 291896 318656
rect 291856 318238 291884 318650
rect 291844 318232 291896 318238
rect 291844 318174 291896 318180
rect 291948 317694 291976 319534
rect 291936 317688 291988 317694
rect 291936 317630 291988 317636
rect 291936 315240 291988 315246
rect 291936 315182 291988 315188
rect 291842 309768 291898 309777
rect 291842 309703 291898 309712
rect 291752 303000 291804 303006
rect 291752 302942 291804 302948
rect 291014 294536 291070 294545
rect 291014 294471 291070 294480
rect 290924 283620 290976 283626
rect 290924 283562 290976 283568
rect 291856 234666 291884 309703
rect 291844 234660 291896 234666
rect 291844 234602 291896 234608
rect 291292 231804 291344 231810
rect 291292 231746 291344 231752
rect 291200 231464 291252 231470
rect 291200 231406 291252 231412
rect 291212 231334 291240 231406
rect 291200 231328 291252 231334
rect 291200 231270 291252 231276
rect 290738 216472 290794 216481
rect 290738 216407 290794 216416
rect 290646 157312 290702 157321
rect 290646 157247 290702 157256
rect 291106 157312 291162 157321
rect 291106 157247 291162 157256
rect 291120 156641 291148 157247
rect 291106 156632 291162 156641
rect 291106 156567 291162 156576
rect 289268 144900 289320 144906
rect 289268 144842 289320 144848
rect 289728 144900 289780 144906
rect 289728 144842 289780 144848
rect 289740 144294 289768 144842
rect 289728 144288 289780 144294
rect 289728 144230 289780 144236
rect 291212 128246 291240 231270
rect 291304 231266 291332 231746
rect 291292 231260 291344 231266
rect 291292 231202 291344 231208
rect 291304 150346 291332 231202
rect 291292 150340 291344 150346
rect 291292 150282 291344 150288
rect 291304 149734 291332 150282
rect 291292 149728 291344 149734
rect 291292 149670 291344 149676
rect 291200 128240 291252 128246
rect 291200 128182 291252 128188
rect 291660 128240 291712 128246
rect 291660 128182 291712 128188
rect 291672 127634 291700 128182
rect 291660 127628 291712 127634
rect 291660 127570 291712 127576
rect 291382 6760 291438 6769
rect 291382 6695 291438 6704
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 289176 3052 289228 3058
rect 289176 2994 289228 3000
rect 290200 480 290228 3470
rect 291396 480 291424 6695
rect 291856 2990 291884 234602
rect 291948 231810 291976 315182
rect 292040 311817 292068 319688
rect 292118 319424 292174 319433
rect 292118 319359 292174 319368
rect 292132 319326 292160 319359
rect 292120 319320 292172 319326
rect 292120 319262 292172 319268
rect 292224 318646 292252 319790
rect 292302 319767 292358 319776
rect 292316 319394 292344 319767
rect 292304 319388 292356 319394
rect 292304 319330 292356 319336
rect 292408 318968 292436 319926
rect 292546 319841 292574 320076
rect 292532 319832 292588 319841
rect 292532 319767 292588 319776
rect 292638 319682 292666 320076
rect 292730 319852 292758 320076
rect 293084 320104 293140 320113
rect 292808 320039 292864 320048
rect 292730 319824 292804 319852
rect 292638 319654 292712 319682
rect 292580 319592 292632 319598
rect 292578 319560 292580 319569
rect 292632 319560 292634 319569
rect 292578 319495 292634 319504
rect 292684 319444 292712 319654
rect 292592 319416 292712 319444
rect 292316 318940 292436 318968
rect 292486 319016 292542 319025
rect 292486 318951 292542 318960
rect 292212 318640 292264 318646
rect 292212 318582 292264 318588
rect 292224 317370 292252 318582
rect 292316 318050 292344 318940
rect 292500 318442 292528 318951
rect 292592 318782 292620 319416
rect 292670 319288 292726 319297
rect 292670 319223 292726 319232
rect 292684 319025 292712 319223
rect 292670 319016 292726 319025
rect 292670 318951 292726 318960
rect 292580 318776 292632 318782
rect 292580 318718 292632 318724
rect 292488 318436 292540 318442
rect 292488 318378 292540 318384
rect 292316 318022 292436 318050
rect 292304 317688 292356 317694
rect 292304 317630 292356 317636
rect 292132 317342 292252 317370
rect 292026 311808 292082 311817
rect 292026 311743 292082 311752
rect 292028 303136 292080 303142
rect 292028 303078 292080 303084
rect 291936 231804 291988 231810
rect 291936 231746 291988 231752
rect 292040 228449 292068 303078
rect 292132 246362 292160 317342
rect 292212 317144 292264 317150
rect 292212 317086 292264 317092
rect 292224 315602 292252 317086
rect 292316 315874 292344 317630
rect 292408 315994 292436 318022
rect 292396 315988 292448 315994
rect 292396 315930 292448 315936
rect 292316 315846 292436 315874
rect 292224 315574 292344 315602
rect 292212 315172 292264 315178
rect 292212 315114 292264 315120
rect 292224 295225 292252 315114
rect 292210 295216 292266 295225
rect 292210 295151 292266 295160
rect 292120 246356 292172 246362
rect 292120 246298 292172 246304
rect 292224 239698 292252 295151
rect 292316 279478 292344 315574
rect 292408 280838 292436 315846
rect 292500 282198 292528 318378
rect 292488 282192 292540 282198
rect 292488 282134 292540 282140
rect 292396 280832 292448 280838
rect 292396 280774 292448 280780
rect 292304 279472 292356 279478
rect 292304 279414 292356 279420
rect 292304 249144 292356 249150
rect 292304 249086 292356 249092
rect 292212 239692 292264 239698
rect 292212 239634 292264 239640
rect 292316 231470 292344 249086
rect 292304 231464 292356 231470
rect 292304 231406 292356 231412
rect 292026 228440 292082 228449
rect 292026 228375 292082 228384
rect 292592 219434 292620 318718
rect 292684 313562 292712 318951
rect 292776 318034 292804 319824
rect 292914 319784 292942 320076
rect 292868 319756 292942 319784
rect 293006 319784 293034 320076
rect 294004 320104 294060 320113
rect 293084 320039 293140 320048
rect 293190 319818 293218 320076
rect 293144 319790 293218 319818
rect 293006 319756 293080 319784
rect 292764 318028 292816 318034
rect 292764 317970 292816 317976
rect 292868 316520 292896 319756
rect 293052 319433 293080 319756
rect 293038 319424 293094 319433
rect 293038 319359 293094 319368
rect 292946 319288 293002 319297
rect 292946 319223 292948 319232
rect 293000 319223 293002 319232
rect 292948 319194 293000 319200
rect 293040 318028 293092 318034
rect 293040 317970 293092 317976
rect 292776 316492 292896 316520
rect 292776 313721 292804 316492
rect 292856 315988 292908 315994
rect 292856 315930 292908 315936
rect 292762 313712 292818 313721
rect 292762 313647 292818 313656
rect 292684 313534 292804 313562
rect 292672 313472 292724 313478
rect 292672 313414 292724 313420
rect 292684 239154 292712 313414
rect 292776 240786 292804 313534
rect 292868 305930 292896 315930
rect 292948 314900 293000 314906
rect 292948 314842 293000 314848
rect 292960 308310 292988 314842
rect 293052 311710 293080 317970
rect 293144 316034 293172 319790
rect 293282 319784 293310 320076
rect 293374 319954 293402 320076
rect 293374 319926 293448 319954
rect 293282 319756 293356 319784
rect 293144 316006 293264 316034
rect 293236 314401 293264 316006
rect 293222 314392 293278 314401
rect 293222 314327 293278 314336
rect 293328 314276 293356 319756
rect 293420 318073 293448 319926
rect 293558 319716 293586 320076
rect 293650 319954 293678 320076
rect 293650 319926 293724 319954
rect 293512 319688 293586 319716
rect 293406 318064 293462 318073
rect 293406 317999 293462 318008
rect 293236 314248 293356 314276
rect 293040 311704 293092 311710
rect 293040 311646 293092 311652
rect 293236 311370 293264 314248
rect 293420 313478 293448 317999
rect 293512 315994 293540 319688
rect 293696 319512 293724 319926
rect 293834 319852 293862 320076
rect 293604 319484 293724 319512
rect 293788 319824 293862 319852
rect 293500 315988 293552 315994
rect 293500 315930 293552 315936
rect 293604 314906 293632 319484
rect 293684 319388 293736 319394
rect 293684 319330 293736 319336
rect 293696 319025 293724 319330
rect 293682 319016 293738 319025
rect 293682 318951 293738 318960
rect 293684 317960 293736 317966
rect 293684 317902 293736 317908
rect 293696 317150 293724 317902
rect 293684 317144 293736 317150
rect 293684 317086 293736 317092
rect 293592 314900 293644 314906
rect 293592 314842 293644 314848
rect 293408 313472 293460 313478
rect 293408 313414 293460 313420
rect 293788 311894 293816 319824
rect 293926 319784 293954 320076
rect 295844 320104 295900 320113
rect 294004 320039 294060 320048
rect 294202 319954 294230 320076
rect 294386 319954 294414 320076
rect 294156 319926 294230 319954
rect 294340 319926 294414 319954
rect 294156 319802 294184 319926
rect 294234 319832 294290 319841
rect 293880 319756 293954 319784
rect 294144 319796 294196 319802
rect 293880 317762 293908 319756
rect 294234 319767 294290 319776
rect 294144 319738 294196 319744
rect 293960 319660 294012 319666
rect 293960 319602 294012 319608
rect 293972 318238 294000 319602
rect 294248 319530 294276 319767
rect 294236 319524 294288 319530
rect 294236 319466 294288 319472
rect 294234 319288 294290 319297
rect 294340 319258 294368 319926
rect 294478 319784 294506 320076
rect 294432 319756 294506 319784
rect 294234 319223 294290 319232
rect 294328 319252 294380 319258
rect 293960 318232 294012 318238
rect 293960 318174 294012 318180
rect 294144 318232 294196 318238
rect 294144 318174 294196 318180
rect 293868 317756 293920 317762
rect 293868 317698 293920 317704
rect 293328 311866 293816 311894
rect 293224 311364 293276 311370
rect 293224 311306 293276 311312
rect 292948 308304 293000 308310
rect 292948 308246 293000 308252
rect 292948 307896 293000 307902
rect 292948 307838 293000 307844
rect 292960 307630 292988 307838
rect 292948 307624 293000 307630
rect 292948 307566 293000 307572
rect 293236 307154 293264 311306
rect 293328 307630 293356 311866
rect 293408 311704 293460 311710
rect 293408 311646 293460 311652
rect 293316 307624 293368 307630
rect 293316 307566 293368 307572
rect 293224 307148 293276 307154
rect 293224 307090 293276 307096
rect 293224 306128 293276 306134
rect 293224 306070 293276 306076
rect 292856 305924 292908 305930
rect 292856 305866 292908 305872
rect 292868 305658 292896 305866
rect 292856 305652 292908 305658
rect 292856 305594 292908 305600
rect 292854 299296 292910 299305
rect 292854 299231 292910 299240
rect 292868 298761 292896 299231
rect 292854 298752 292910 298761
rect 292854 298687 292910 298696
rect 292764 240780 292816 240786
rect 292764 240722 292816 240728
rect 292672 239148 292724 239154
rect 292672 239090 292724 239096
rect 292672 227248 292724 227254
rect 292672 227190 292724 227196
rect 292684 227050 292712 227190
rect 292672 227044 292724 227050
rect 292672 226986 292724 226992
rect 292580 219428 292632 219434
rect 292580 219370 292632 219376
rect 292868 216646 292896 298687
rect 293236 234326 293264 306070
rect 293316 304496 293368 304502
rect 293316 304438 293368 304444
rect 293224 234320 293276 234326
rect 293224 234262 293276 234268
rect 293224 227044 293276 227050
rect 293224 226986 293276 226992
rect 292856 216640 292908 216646
rect 292856 216582 292908 216588
rect 293236 125497 293264 226986
rect 293328 224398 293356 304438
rect 293420 301510 293448 311646
rect 293960 308780 294012 308786
rect 293960 308722 294012 308728
rect 293972 308446 294000 308722
rect 294052 308712 294104 308718
rect 294052 308654 294104 308660
rect 293960 308440 294012 308446
rect 293960 308382 294012 308388
rect 293960 307828 294012 307834
rect 293960 307770 294012 307776
rect 293972 307222 294000 307770
rect 293960 307216 294012 307222
rect 293960 307158 294012 307164
rect 294064 307154 294092 308654
rect 294052 307148 294104 307154
rect 294052 307090 294104 307096
rect 294156 303142 294184 318174
rect 294248 307426 294276 319223
rect 294328 319194 294380 319200
rect 294340 318918 294368 319194
rect 294328 318912 294380 318918
rect 294328 318854 294380 318860
rect 294432 316282 294460 319756
rect 294570 319546 294598 320076
rect 294754 319954 294782 320076
rect 294708 319926 294782 319954
rect 294570 319518 294644 319546
rect 294510 319424 294566 319433
rect 294510 319359 294566 319368
rect 294340 316254 294460 316282
rect 294524 316266 294552 319359
rect 294616 318753 294644 319518
rect 294602 318744 294658 318753
rect 294602 318679 294658 318688
rect 294512 316260 294564 316266
rect 294340 308718 294368 316254
rect 294512 316202 294564 316208
rect 294708 316146 294736 319926
rect 294846 319852 294874 320076
rect 294432 316118 294736 316146
rect 294800 319824 294874 319852
rect 294432 308786 294460 316118
rect 294800 316062 294828 319824
rect 294938 319784 294966 320076
rect 295122 319784 295150 320076
rect 294892 319756 294966 319784
rect 295076 319756 295150 319784
rect 294788 316056 294840 316062
rect 294788 315998 294840 316004
rect 294512 315988 294564 315994
rect 294512 315930 294564 315936
rect 294524 309806 294552 315930
rect 294892 313002 294920 319756
rect 294970 319696 295026 319705
rect 294970 319631 295026 319640
rect 294984 319598 295012 319631
rect 294972 319592 295024 319598
rect 294972 319534 295024 319540
rect 294972 319456 295024 319462
rect 294972 319398 295024 319404
rect 294984 318918 295012 319398
rect 294972 318912 295024 318918
rect 294972 318854 295024 318860
rect 295076 316674 295104 319756
rect 295214 319716 295242 320076
rect 295306 319784 295334 320076
rect 295490 319852 295518 320076
rect 295444 319824 295518 319852
rect 295306 319756 295380 319784
rect 295168 319688 295242 319716
rect 295064 316668 295116 316674
rect 295064 316610 295116 316616
rect 294972 316260 295024 316266
rect 294972 316202 295024 316208
rect 294880 312996 294932 313002
rect 294880 312938 294932 312944
rect 294694 312624 294750 312633
rect 294694 312559 294750 312568
rect 294512 309800 294564 309806
rect 294512 309742 294564 309748
rect 294420 308780 294472 308786
rect 294420 308722 294472 308728
rect 294328 308712 294380 308718
rect 294328 308654 294380 308660
rect 294236 307420 294288 307426
rect 294236 307362 294288 307368
rect 294248 306374 294276 307362
rect 294248 306346 294644 306374
rect 294144 303136 294196 303142
rect 294144 303078 294196 303084
rect 293408 301504 293460 301510
rect 293408 301446 293460 301452
rect 294050 237008 294106 237017
rect 294050 236943 294106 236952
rect 294064 236065 294092 236943
rect 294050 236056 294106 236065
rect 294050 235991 294106 236000
rect 293316 224392 293368 224398
rect 293316 224334 293368 224340
rect 294064 146266 294092 235991
rect 294616 227458 294644 306346
rect 294604 227452 294656 227458
rect 294604 227394 294656 227400
rect 294604 221468 294656 221474
rect 294604 221410 294656 221416
rect 294052 146260 294104 146266
rect 294052 146202 294104 146208
rect 294616 132494 294644 221410
rect 294708 219162 294736 312559
rect 294892 311894 294920 312938
rect 294800 311866 294920 311894
rect 294800 237250 294828 311866
rect 294984 307222 295012 316202
rect 295064 316056 295116 316062
rect 295064 315998 295116 316004
rect 294972 307216 295024 307222
rect 294972 307158 295024 307164
rect 294878 305824 294934 305833
rect 294878 305759 294934 305768
rect 294788 237244 294840 237250
rect 294788 237186 294840 237192
rect 294892 231606 294920 305759
rect 295076 299334 295104 315998
rect 295168 315994 295196 319688
rect 295248 319320 295300 319326
rect 295248 319262 295300 319268
rect 295156 315988 295208 315994
rect 295156 315930 295208 315936
rect 295064 299328 295116 299334
rect 295064 299270 295116 299276
rect 295076 296714 295104 299270
rect 294984 296686 295104 296714
rect 294984 240922 295012 296686
rect 295064 260160 295116 260166
rect 295064 260102 295116 260108
rect 294972 240916 295024 240922
rect 294972 240858 295024 240864
rect 295076 236065 295104 260102
rect 295062 236056 295118 236065
rect 295062 235991 295118 236000
rect 294880 231600 294932 231606
rect 294880 231542 294932 231548
rect 295260 228546 295288 319262
rect 295352 318238 295380 319756
rect 295444 319734 295472 319824
rect 295582 319784 295610 320076
rect 295536 319756 295610 319784
rect 295432 319728 295484 319734
rect 295432 319670 295484 319676
rect 295432 319456 295484 319462
rect 295432 319398 295484 319404
rect 295444 318850 295472 319398
rect 295432 318844 295484 318850
rect 295432 318786 295484 318792
rect 295340 318232 295392 318238
rect 295340 318174 295392 318180
rect 295536 316146 295564 319756
rect 295674 319734 295702 320076
rect 295766 319784 295794 320076
rect 296212 320104 296268 320113
rect 295844 320039 295900 320048
rect 295950 319784 295978 320076
rect 295766 319756 295840 319784
rect 295662 319728 295714 319734
rect 295662 319670 295714 319676
rect 295812 319666 295840 319756
rect 295904 319756 295978 319784
rect 296134 319784 296162 320076
rect 297224 320104 297280 320113
rect 296212 320039 296268 320048
rect 296318 319818 296346 320076
rect 296272 319790 296346 319818
rect 296410 319818 296438 320076
rect 296410 319790 296484 319818
rect 296134 319756 296208 319784
rect 295800 319660 295852 319666
rect 295800 319602 295852 319608
rect 295708 319592 295760 319598
rect 295708 319534 295760 319540
rect 295616 319524 295668 319530
rect 295616 319466 295668 319472
rect 295444 316118 295564 316146
rect 295444 312934 295472 316118
rect 295524 315988 295576 315994
rect 295524 315930 295576 315936
rect 295432 312928 295484 312934
rect 295432 312870 295484 312876
rect 295340 311840 295392 311846
rect 295340 311782 295392 311788
rect 295352 310593 295380 311782
rect 295338 310584 295394 310593
rect 295338 310519 295394 310528
rect 295444 310078 295472 312870
rect 295432 310072 295484 310078
rect 295432 310014 295484 310020
rect 295340 304904 295392 304910
rect 295340 304846 295392 304852
rect 295352 304298 295380 304846
rect 295340 304292 295392 304298
rect 295340 304234 295392 304240
rect 295340 303204 295392 303210
rect 295340 303146 295392 303152
rect 295352 302938 295380 303146
rect 295536 303074 295564 315930
rect 295628 304910 295656 319466
rect 295720 319138 295748 319534
rect 295798 319424 295854 319433
rect 295798 319359 295854 319368
rect 295812 319326 295840 319359
rect 295800 319320 295852 319326
rect 295800 319262 295852 319268
rect 295720 319110 295840 319138
rect 295904 319122 295932 319756
rect 296074 319288 296130 319297
rect 296074 319223 296130 319232
rect 295706 319016 295762 319025
rect 295706 318951 295762 318960
rect 295720 309874 295748 318951
rect 295812 318617 295840 319110
rect 295892 319116 295944 319122
rect 295892 319058 295944 319064
rect 295984 319116 296036 319122
rect 295984 319058 296036 319064
rect 295996 318782 296024 319058
rect 295984 318776 296036 318782
rect 295984 318718 296036 318724
rect 295798 318608 295854 318617
rect 295798 318543 295854 318552
rect 295984 317552 296036 317558
rect 295984 317494 296036 317500
rect 295708 309868 295760 309874
rect 295708 309810 295760 309816
rect 295616 304904 295668 304910
rect 295616 304846 295668 304852
rect 295524 303068 295576 303074
rect 295524 303010 295576 303016
rect 295340 302932 295392 302938
rect 295340 302874 295392 302880
rect 295248 228540 295300 228546
rect 295248 228482 295300 228488
rect 295996 225690 296024 317494
rect 296088 316742 296116 319223
rect 296076 316736 296128 316742
rect 296076 316678 296128 316684
rect 296180 315994 296208 319756
rect 296272 318578 296300 319790
rect 296352 319728 296404 319734
rect 296352 319670 296404 319676
rect 296260 318572 296312 318578
rect 296260 318514 296312 318520
rect 296260 317620 296312 317626
rect 296260 317562 296312 317568
rect 296168 315988 296220 315994
rect 296168 315930 296220 315936
rect 296272 314430 296300 317562
rect 296260 314424 296312 314430
rect 296260 314366 296312 314372
rect 296076 305992 296128 305998
rect 296076 305934 296128 305940
rect 296258 305960 296314 305969
rect 296088 238921 296116 305934
rect 296258 305895 296314 305904
rect 296166 302152 296222 302161
rect 296166 302087 296222 302096
rect 296074 238912 296130 238921
rect 296074 238847 296130 238856
rect 296076 236836 296128 236842
rect 296076 236778 296128 236784
rect 295984 225684 296036 225690
rect 295984 225626 296036 225632
rect 294696 219156 294748 219162
rect 294696 219098 294748 219104
rect 295984 151088 296036 151094
rect 295984 151030 296036 151036
rect 295338 147656 295394 147665
rect 295338 147591 295394 147600
rect 295352 146985 295380 147591
rect 295338 146976 295394 146985
rect 295338 146911 295394 146920
rect 294880 146260 294932 146266
rect 294880 146202 294932 146208
rect 294892 145586 294920 146202
rect 294880 145580 294932 145586
rect 294880 145522 294932 145528
rect 294524 132466 294644 132494
rect 292578 125488 292634 125497
rect 292578 125423 292634 125432
rect 293222 125488 293278 125497
rect 293222 125423 293278 125432
rect 292592 124817 292620 125423
rect 292578 124808 292634 124817
rect 292578 124743 292634 124752
rect 294524 124166 294552 132466
rect 294512 124160 294564 124166
rect 294512 124102 294564 124108
rect 294524 123486 294552 124102
rect 294512 123480 294564 123486
rect 294512 123422 294564 123428
rect 294878 6624 294934 6633
rect 294878 6559 294934 6568
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 291844 2984 291896 2990
rect 291844 2926 291896 2932
rect 292592 480 292620 3538
rect 293684 2984 293736 2990
rect 293684 2926 293736 2932
rect 293696 480 293724 2926
rect 294892 480 294920 6559
rect 295996 3602 296024 151030
rect 296088 146985 296116 236778
rect 296180 218657 296208 302087
rect 296272 232966 296300 305895
rect 296364 302122 296392 319670
rect 296456 319530 296484 319790
rect 296594 319784 296622 320076
rect 296548 319756 296622 319784
rect 296444 319524 296496 319530
rect 296444 319466 296496 319472
rect 296444 318844 296496 318850
rect 296444 318786 296496 318792
rect 296456 303210 296484 318786
rect 296548 318510 296576 319756
rect 296686 319648 296714 320076
rect 296778 319716 296806 320076
rect 296870 319784 296898 320076
rect 297146 319954 297174 320076
rect 297592 320104 297648 320113
rect 297224 320039 297280 320048
rect 297330 319954 297358 320076
rect 297100 319926 297174 319954
rect 297284 319926 297358 319954
rect 296870 319756 296944 319784
rect 296778 319688 296852 319716
rect 296640 319620 296714 319648
rect 296640 318850 296668 319620
rect 296718 319288 296774 319297
rect 296718 319223 296774 319232
rect 296628 318844 296680 318850
rect 296628 318786 296680 318792
rect 296536 318504 296588 318510
rect 296536 318446 296588 318452
rect 296732 317626 296760 319223
rect 296720 317620 296772 317626
rect 296720 317562 296772 317568
rect 296536 316736 296588 316742
rect 296536 316678 296588 316684
rect 296626 316704 296682 316713
rect 296548 316538 296576 316678
rect 296626 316639 296682 316648
rect 296536 316532 296588 316538
rect 296536 316474 296588 316480
rect 296534 312488 296590 312497
rect 296534 312423 296590 312432
rect 296444 303204 296496 303210
rect 296444 303146 296496 303152
rect 296352 302116 296404 302122
rect 296352 302058 296404 302064
rect 296548 238814 296576 312423
rect 296640 238882 296668 316639
rect 296824 315994 296852 319688
rect 296916 319297 296944 319756
rect 296902 319288 296958 319297
rect 296902 319223 296958 319232
rect 296902 318880 296958 318889
rect 296902 318815 296958 318824
rect 296812 315988 296864 315994
rect 296812 315930 296864 315936
rect 296812 315784 296864 315790
rect 296812 315726 296864 315732
rect 296824 302258 296852 315726
rect 296916 304366 296944 318815
rect 296996 318776 297048 318782
rect 296996 318718 297048 318724
rect 297008 317898 297036 318718
rect 297100 318306 297128 319926
rect 297284 319716 297312 319926
rect 297422 319784 297450 320076
rect 297514 319920 297542 320076
rect 297776 320104 297832 320113
rect 297592 320039 297648 320048
rect 297698 319920 297726 320076
rect 298420 320104 298476 320113
rect 297776 320039 297832 320048
rect 297514 319892 297588 319920
rect 297422 319756 297496 319784
rect 297284 319688 297404 319716
rect 297272 319592 297324 319598
rect 297272 319534 297324 319540
rect 297284 319444 297312 319534
rect 297192 319416 297312 319444
rect 297088 318300 297140 318306
rect 297088 318242 297140 318248
rect 296996 317892 297048 317898
rect 296996 317834 297048 317840
rect 297192 310010 297220 319416
rect 297376 319025 297404 319688
rect 297468 319598 297496 319756
rect 297456 319592 297508 319598
rect 297456 319534 297508 319540
rect 297454 319288 297510 319297
rect 297454 319223 297510 319232
rect 297362 319016 297418 319025
rect 297362 318951 297418 318960
rect 297272 318708 297324 318714
rect 297272 318650 297324 318656
rect 297284 317898 297312 318650
rect 297362 318608 297418 318617
rect 297362 318543 297418 318552
rect 297376 318209 297404 318543
rect 297362 318200 297418 318209
rect 297362 318135 297418 318144
rect 297468 318034 297496 319223
rect 297560 319025 297588 319892
rect 297652 319892 297726 319920
rect 297652 319104 297680 319892
rect 297882 319818 297910 320076
rect 297744 319790 297910 319818
rect 297744 319433 297772 319790
rect 297974 319784 298002 320076
rect 298066 319954 298094 320076
rect 298066 319926 298140 319954
rect 297974 319756 298048 319784
rect 297730 319424 297786 319433
rect 297730 319359 297786 319368
rect 297652 319076 297956 319104
rect 297546 319016 297602 319025
rect 297546 318951 297602 318960
rect 297730 319016 297786 319025
rect 297730 318951 297786 318960
rect 297546 318472 297602 318481
rect 297546 318407 297602 318416
rect 297456 318028 297508 318034
rect 297456 317970 297508 317976
rect 297272 317892 297324 317898
rect 297272 317834 297324 317840
rect 297560 317354 297588 318407
rect 297548 317348 297600 317354
rect 297548 317290 297600 317296
rect 297548 315988 297600 315994
rect 297548 315930 297600 315936
rect 297364 310412 297416 310418
rect 297364 310354 297416 310360
rect 297180 310004 297232 310010
rect 297180 309946 297232 309952
rect 296904 304360 296956 304366
rect 296904 304302 296956 304308
rect 296812 302252 296864 302258
rect 296812 302194 296864 302200
rect 296628 238876 296680 238882
rect 296628 238818 296680 238824
rect 296536 238808 296588 238814
rect 296536 238754 296588 238756
rect 296364 238750 296588 238754
rect 296364 238726 296576 238750
rect 296260 232960 296312 232966
rect 296260 232902 296312 232908
rect 296364 227225 296392 238726
rect 296640 231577 296668 238818
rect 296626 231568 296682 231577
rect 296626 231503 296682 231512
rect 296350 227216 296406 227225
rect 296350 227151 296406 227160
rect 297376 225622 297404 310354
rect 297456 303748 297508 303754
rect 297456 303690 297508 303696
rect 296720 225616 296772 225622
rect 296720 225558 296772 225564
rect 297364 225616 297416 225622
rect 297364 225558 297416 225564
rect 296166 218648 296222 218657
rect 296166 218583 296222 218592
rect 296074 146976 296130 146985
rect 296074 146911 296130 146920
rect 296732 16574 296760 225558
rect 297468 224330 297496 303690
rect 297560 302190 297588 315930
rect 297744 315790 297772 318951
rect 297928 317948 297956 319076
rect 298020 318714 298048 319756
rect 298008 318708 298060 318714
rect 298008 318650 298060 318656
rect 298008 318504 298060 318510
rect 298008 318446 298060 318452
rect 298020 318102 298048 318446
rect 298008 318096 298060 318102
rect 298008 318038 298060 318044
rect 297928 317920 298048 317948
rect 297916 317484 297968 317490
rect 297916 317426 297968 317432
rect 297732 315784 297784 315790
rect 297732 315726 297784 315732
rect 297640 314492 297692 314498
rect 297640 314434 297692 314440
rect 297652 314226 297680 314434
rect 297640 314220 297692 314226
rect 297640 314162 297692 314168
rect 297548 302184 297600 302190
rect 297548 302126 297600 302132
rect 297560 301782 297588 302126
rect 297548 301776 297600 301782
rect 297548 301718 297600 301724
rect 297652 239018 297680 314162
rect 297928 311846 297956 317426
rect 298020 314498 298048 317920
rect 298008 314492 298060 314498
rect 298008 314434 298060 314440
rect 298008 314152 298060 314158
rect 298008 314094 298060 314100
rect 297916 311840 297968 311846
rect 297916 311782 297968 311788
rect 298020 311438 298048 314094
rect 298008 311432 298060 311438
rect 298008 311374 298060 311380
rect 297824 310140 297876 310146
rect 297824 310082 297876 310088
rect 297730 306232 297786 306241
rect 297730 306167 297786 306176
rect 297640 239012 297692 239018
rect 297640 238954 297692 238960
rect 297744 232898 297772 306167
rect 297836 239086 297864 310082
rect 298112 307358 298140 319926
rect 298250 319852 298278 320076
rect 298204 319824 298278 319852
rect 298204 317286 298232 319824
rect 298342 319784 298370 320076
rect 299064 320104 299120 320113
rect 298420 320039 298476 320048
rect 298618 319920 298646 320076
rect 298802 319954 298830 320076
rect 298572 319892 298646 319920
rect 298756 319926 298830 319954
rect 298342 319756 298416 319784
rect 298388 317490 298416 319756
rect 298376 317484 298428 317490
rect 298376 317426 298428 317432
rect 298192 317280 298244 317286
rect 298192 317222 298244 317228
rect 298284 316668 298336 316674
rect 298572 316656 298600 319892
rect 298756 319870 298784 319926
rect 298744 319864 298796 319870
rect 298664 319812 298744 319818
rect 298664 319806 298796 319812
rect 298894 319818 298922 320076
rect 298986 319954 299014 320076
rect 299432 320104 299488 320113
rect 299064 320039 299120 320048
rect 298986 319926 299060 319954
rect 299032 319920 299060 319926
rect 299032 319892 299244 319920
rect 298664 319790 298784 319806
rect 298894 319790 298968 319818
rect 298664 319666 298692 319790
rect 298744 319728 298796 319734
rect 298744 319670 298796 319676
rect 298836 319728 298888 319734
rect 298836 319670 298888 319676
rect 298652 319660 298704 319666
rect 298652 319602 298704 319608
rect 298756 319025 298784 319670
rect 298742 319016 298798 319025
rect 298742 318951 298798 318960
rect 298848 317422 298876 319670
rect 298940 318850 298968 319790
rect 299020 319796 299072 319802
rect 299020 319738 299072 319744
rect 298928 318844 298980 318850
rect 298928 318786 298980 318792
rect 298928 318708 298980 318714
rect 298928 318650 298980 318656
rect 298836 317416 298888 317422
rect 298836 317358 298888 317364
rect 298572 316628 298784 316656
rect 298284 316610 298336 316616
rect 298296 311234 298324 316610
rect 298650 316568 298706 316577
rect 298650 316503 298706 316512
rect 298374 316432 298430 316441
rect 298374 316367 298430 316376
rect 298284 311228 298336 311234
rect 298284 311170 298336 311176
rect 298284 308304 298336 308310
rect 298284 308246 298336 308252
rect 298100 307352 298152 307358
rect 298100 307294 298152 307300
rect 298008 302932 298060 302938
rect 298008 302874 298060 302880
rect 298020 302258 298048 302874
rect 298008 302252 298060 302258
rect 298008 302194 298060 302200
rect 297916 301776 297968 301782
rect 297916 301718 297968 301724
rect 297928 293321 297956 301718
rect 297914 293312 297970 293321
rect 297914 293247 297970 293256
rect 297824 239080 297876 239086
rect 297824 239022 297876 239028
rect 297732 232892 297784 232898
rect 297732 232834 297784 232840
rect 298020 224942 298048 302194
rect 298190 237144 298246 237153
rect 298190 237079 298246 237088
rect 298008 224936 298060 224942
rect 298008 224878 298060 224884
rect 297456 224324 297508 224330
rect 297456 224266 297508 224272
rect 298100 171148 298152 171154
rect 298100 171090 298152 171096
rect 296732 16546 297312 16574
rect 295984 3596 296036 3602
rect 295984 3538 296036 3544
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296088 480 296116 2994
rect 297284 480 297312 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 171090
rect 298204 150385 298232 237079
rect 298296 224806 298324 308246
rect 298388 301510 298416 316367
rect 298558 316296 298614 316305
rect 298558 316231 298614 316240
rect 298572 304026 298600 316231
rect 298664 304638 298692 316503
rect 298756 313682 298784 316628
rect 298836 316260 298888 316266
rect 298836 316202 298888 316208
rect 298744 313676 298796 313682
rect 298744 313618 298796 313624
rect 298652 304632 298704 304638
rect 298652 304574 298704 304580
rect 298560 304020 298612 304026
rect 298560 303962 298612 303968
rect 298664 303686 298692 304574
rect 298652 303680 298704 303686
rect 298652 303622 298704 303628
rect 298376 301504 298428 301510
rect 298376 301446 298428 301452
rect 298388 297537 298416 301446
rect 298374 297528 298430 297537
rect 298374 297463 298430 297472
rect 298284 224800 298336 224806
rect 298284 224742 298336 224748
rect 298756 224670 298784 313618
rect 298848 237153 298876 316202
rect 298940 310146 298968 318650
rect 299032 317218 299060 319738
rect 299112 318844 299164 318850
rect 299112 318786 299164 318792
rect 299020 317212 299072 317218
rect 299020 317154 299072 317160
rect 299124 311894 299152 318786
rect 299032 311866 299152 311894
rect 298928 310140 298980 310146
rect 298928 310082 298980 310088
rect 299032 309244 299060 311866
rect 299112 311772 299164 311778
rect 299112 311714 299164 311720
rect 299124 311234 299152 311714
rect 299112 311228 299164 311234
rect 299112 311170 299164 311176
rect 299112 310480 299164 310486
rect 299112 310422 299164 310428
rect 299124 309777 299152 310422
rect 299110 309768 299166 309777
rect 299110 309703 299166 309712
rect 299032 309216 299152 309244
rect 299124 304162 299152 309216
rect 299112 304156 299164 304162
rect 299112 304098 299164 304104
rect 299020 303680 299072 303686
rect 299020 303622 299072 303628
rect 298926 298888 298982 298897
rect 298926 298823 298982 298832
rect 298834 237144 298890 237153
rect 298834 237079 298890 237088
rect 298744 224664 298796 224670
rect 298744 224606 298796 224612
rect 298940 222873 298968 298823
rect 299032 228886 299060 303622
rect 299124 240854 299152 304098
rect 299216 302161 299244 319892
rect 299354 319784 299382 320076
rect 300076 320104 300132 320113
rect 299432 320039 299488 320048
rect 299538 319784 299566 320076
rect 299308 319756 299382 319784
rect 299492 319756 299566 319784
rect 299308 316674 299336 319756
rect 299492 319598 299520 319756
rect 299630 319682 299658 320076
rect 299722 319716 299750 320076
rect 299814 319784 299842 320076
rect 299906 319938 299934 320076
rect 300076 320039 300132 320048
rect 300260 320104 300316 320113
rect 300904 320104 300960 320113
rect 300260 320039 300316 320048
rect 299894 319932 299946 319938
rect 300366 319920 300394 320076
rect 299894 319874 299946 319880
rect 300320 319892 300394 319920
rect 299814 319756 300072 319784
rect 299722 319688 299796 319716
rect 299584 319654 299658 319682
rect 299480 319592 299532 319598
rect 299480 319534 299532 319540
rect 299584 319054 299612 319654
rect 299768 319648 299796 319688
rect 299768 319620 299888 319648
rect 299664 319592 299716 319598
rect 299716 319552 299796 319580
rect 299664 319534 299716 319540
rect 299572 319048 299624 319054
rect 299386 319016 299442 319025
rect 299572 318990 299624 318996
rect 299386 318951 299442 318960
rect 299296 316668 299348 316674
rect 299296 316610 299348 316616
rect 299294 316024 299350 316033
rect 299294 315959 299350 315968
rect 299202 302152 299258 302161
rect 299202 302087 299258 302096
rect 299112 240848 299164 240854
rect 299112 240790 299164 240796
rect 299308 239766 299336 315959
rect 299400 299441 299428 318951
rect 299662 318880 299718 318889
rect 299662 318815 299664 318824
rect 299716 318815 299718 318824
rect 299664 318786 299716 318792
rect 299664 318572 299716 318578
rect 299664 318514 299716 318520
rect 299572 317756 299624 317762
rect 299572 317698 299624 317704
rect 299480 317144 299532 317150
rect 299480 317086 299532 317092
rect 299492 316169 299520 317086
rect 299478 316160 299534 316169
rect 299478 316095 299534 316104
rect 299480 314356 299532 314362
rect 299480 314298 299532 314304
rect 299492 313993 299520 314298
rect 299478 313984 299534 313993
rect 299478 313919 299534 313928
rect 299584 311894 299612 317698
rect 299676 317558 299704 318514
rect 299664 317552 299716 317558
rect 299664 317494 299716 317500
rect 299664 315920 299716 315926
rect 299664 315862 299716 315868
rect 299492 311866 299612 311894
rect 299492 307494 299520 311866
rect 299480 307488 299532 307494
rect 299480 307430 299532 307436
rect 299676 304706 299704 315862
rect 299768 305454 299796 319552
rect 299860 317626 299888 319620
rect 299938 319424 299994 319433
rect 299938 319359 299994 319368
rect 299952 318170 299980 319359
rect 299940 318164 299992 318170
rect 299940 318106 299992 318112
rect 299848 317620 299900 317626
rect 299848 317562 299900 317568
rect 299940 316056 299992 316062
rect 299940 315998 299992 316004
rect 299848 315988 299900 315994
rect 299848 315930 299900 315936
rect 299860 311302 299888 315930
rect 299848 311296 299900 311302
rect 299848 311238 299900 311244
rect 299952 311234 299980 315998
rect 299940 311228 299992 311234
rect 299940 311170 299992 311176
rect 299952 307086 299980 311170
rect 299940 307080 299992 307086
rect 299940 307022 299992 307028
rect 299756 305448 299808 305454
rect 299756 305390 299808 305396
rect 299664 304700 299716 304706
rect 299664 304642 299716 304648
rect 299572 304292 299624 304298
rect 299572 304234 299624 304240
rect 299584 304026 299612 304234
rect 299572 304020 299624 304026
rect 299572 303962 299624 303968
rect 299386 299432 299442 299441
rect 299386 299367 299442 299376
rect 299296 239760 299348 239766
rect 299296 239702 299348 239708
rect 299020 228880 299072 228886
rect 299020 228822 299072 228828
rect 299584 224602 299612 303962
rect 299676 303686 299704 304642
rect 299664 303680 299716 303686
rect 299664 303622 299716 303628
rect 300044 302841 300072 319756
rect 300216 319048 300268 319054
rect 300214 319016 300216 319025
rect 300268 319016 300270 319025
rect 300214 318951 300270 318960
rect 300122 318880 300178 318889
rect 300122 318815 300178 318824
rect 300136 317529 300164 318815
rect 300228 318578 300256 318951
rect 300216 318572 300268 318578
rect 300216 318514 300268 318520
rect 300214 318064 300270 318073
rect 300214 317999 300270 318008
rect 300122 317520 300178 317529
rect 300122 317455 300178 317464
rect 300228 311166 300256 317999
rect 300320 314294 300348 319892
rect 300458 319852 300486 320076
rect 300642 319852 300670 320076
rect 300412 319824 300486 319852
rect 300596 319824 300670 319852
rect 300412 315994 300440 319824
rect 300490 319424 300546 319433
rect 300490 319359 300546 319368
rect 300400 315988 300452 315994
rect 300400 315930 300452 315936
rect 300308 314288 300360 314294
rect 300308 314230 300360 314236
rect 300216 311160 300268 311166
rect 300216 311102 300268 311108
rect 300308 309120 300360 309126
rect 300308 309062 300360 309068
rect 300216 308440 300268 308446
rect 300216 308382 300268 308388
rect 300124 303680 300176 303686
rect 300124 303622 300176 303628
rect 300030 302832 300086 302841
rect 300030 302767 300086 302776
rect 300044 302734 300072 302767
rect 300032 302728 300084 302734
rect 300032 302670 300084 302676
rect 299664 236700 299716 236706
rect 299664 236642 299716 236648
rect 299676 236026 299704 236642
rect 299664 236020 299716 236026
rect 299664 235962 299716 235968
rect 299572 224596 299624 224602
rect 299572 224538 299624 224544
rect 298926 222864 298982 222873
rect 298926 222799 298982 222808
rect 298190 150376 298246 150385
rect 298190 150311 298246 150320
rect 299386 150376 299442 150385
rect 299386 150311 299442 150320
rect 299400 149705 299428 150311
rect 299386 149696 299442 149705
rect 299386 149631 299442 149640
rect 299676 16574 299704 235962
rect 300136 224534 300164 303622
rect 300228 230314 300256 308382
rect 300320 233102 300348 309062
rect 300504 304230 300532 319359
rect 300596 318753 300624 319824
rect 300734 319784 300762 320076
rect 300826 319954 300854 320076
rect 302836 320104 302892 320113
rect 300904 320039 300960 320048
rect 300826 319926 300900 319954
rect 300688 319756 300762 319784
rect 300582 318744 300638 318753
rect 300582 318679 300638 318688
rect 300596 317801 300624 318679
rect 300582 317792 300638 317801
rect 300582 317727 300638 317736
rect 300584 317620 300636 317626
rect 300584 317562 300636 317568
rect 300596 314158 300624 317562
rect 300688 316062 300716 319756
rect 300872 319682 300900 319926
rect 301010 319920 301038 320076
rect 300780 319654 300900 319682
rect 300964 319892 301038 319920
rect 300676 316056 300728 316062
rect 300676 315998 300728 316004
rect 300780 315926 300808 319654
rect 300964 317762 300992 319892
rect 301102 319784 301130 320076
rect 301194 319938 301222 320076
rect 301182 319932 301234 319938
rect 301182 319874 301234 319880
rect 301378 319852 301406 320076
rect 301332 319824 301406 319852
rect 301332 319784 301360 319824
rect 301470 319784 301498 320076
rect 301056 319756 301130 319784
rect 301240 319756 301360 319784
rect 301424 319756 301498 319784
rect 301562 319784 301590 320076
rect 301654 319938 301682 320076
rect 301642 319932 301694 319938
rect 301642 319874 301694 319880
rect 301562 319756 301636 319784
rect 300952 317756 301004 317762
rect 300952 317698 301004 317704
rect 300952 317620 301004 317626
rect 300952 317562 301004 317568
rect 300860 316260 300912 316266
rect 300860 316202 300912 316208
rect 300768 315920 300820 315926
rect 300768 315862 300820 315868
rect 300872 314362 300900 316202
rect 300860 314356 300912 314362
rect 300860 314298 300912 314304
rect 300584 314152 300636 314158
rect 300584 314094 300636 314100
rect 300768 311432 300820 311438
rect 300768 311374 300820 311380
rect 300676 311296 300728 311302
rect 300676 311238 300728 311244
rect 300688 311030 300716 311238
rect 300780 311166 300808 311374
rect 300768 311160 300820 311166
rect 300768 311102 300820 311108
rect 300676 311024 300728 311030
rect 300676 310966 300728 310972
rect 300584 305448 300636 305454
rect 300584 305390 300636 305396
rect 300492 304224 300544 304230
rect 300492 304166 300544 304172
rect 300400 300688 300452 300694
rect 300400 300630 300452 300636
rect 300412 236026 300440 300630
rect 300400 236020 300452 236026
rect 300400 235962 300452 235968
rect 300308 233096 300360 233102
rect 300308 233038 300360 233044
rect 300504 231742 300532 304166
rect 300596 293185 300624 305390
rect 300964 304774 300992 317562
rect 300952 304768 301004 304774
rect 300952 304710 301004 304716
rect 300964 304502 300992 304710
rect 300952 304496 301004 304502
rect 300952 304438 301004 304444
rect 301056 304434 301084 319756
rect 301136 319660 301188 319666
rect 301136 319602 301188 319608
rect 301148 316266 301176 319602
rect 301136 316260 301188 316266
rect 301136 316202 301188 316208
rect 301240 315976 301268 319756
rect 301320 319660 301372 319666
rect 301320 319602 301372 319608
rect 301148 315948 301268 315976
rect 301148 304502 301176 315948
rect 301332 315874 301360 319602
rect 301424 317529 301452 319756
rect 301502 319424 301558 319433
rect 301502 319359 301558 319368
rect 301410 317520 301466 317529
rect 301410 317455 301466 317464
rect 301240 315846 301360 315874
rect 301240 304570 301268 315846
rect 301516 315772 301544 319359
rect 301332 315744 301544 315772
rect 301332 308802 301360 315744
rect 301504 312520 301556 312526
rect 301504 312462 301556 312468
rect 301410 308816 301466 308825
rect 301332 308774 301410 308802
rect 301410 308751 301466 308760
rect 301424 308417 301452 308751
rect 301410 308408 301466 308417
rect 301410 308343 301466 308352
rect 301228 304564 301280 304570
rect 301228 304506 301280 304512
rect 301136 304496 301188 304502
rect 301136 304438 301188 304444
rect 301044 304428 301096 304434
rect 301044 304370 301096 304376
rect 301056 303686 301084 304370
rect 301148 303754 301176 304438
rect 301136 303748 301188 303754
rect 301136 303690 301188 303696
rect 301044 303680 301096 303686
rect 301044 303622 301096 303628
rect 300768 301844 300820 301850
rect 300768 301786 300820 301792
rect 300780 301617 300808 301786
rect 300766 301608 300822 301617
rect 300766 301543 300822 301552
rect 300582 293176 300638 293185
rect 300582 293111 300638 293120
rect 300492 231736 300544 231742
rect 300492 231678 300544 231684
rect 301516 230450 301544 312462
rect 301608 311574 301636 319756
rect 301746 319648 301774 320076
rect 301838 319716 301866 320076
rect 301930 319852 301958 320076
rect 302022 319954 302050 320076
rect 302022 319926 302096 319954
rect 302206 319938 302234 320076
rect 302068 319920 302096 319926
rect 302194 319932 302246 319938
rect 302068 319892 302142 319920
rect 301930 319824 302004 319852
rect 301838 319688 301912 319716
rect 301746 319620 301820 319648
rect 301686 319016 301742 319025
rect 301686 318951 301742 318960
rect 301700 318918 301728 318951
rect 301688 318912 301740 318918
rect 301688 318854 301740 318860
rect 301792 317529 301820 319620
rect 301778 317520 301834 317529
rect 301778 317455 301834 317464
rect 301884 312526 301912 319688
rect 301872 312520 301924 312526
rect 301872 312462 301924 312468
rect 301596 311568 301648 311574
rect 301596 311510 301648 311516
rect 301688 308984 301740 308990
rect 301688 308926 301740 308932
rect 301596 303680 301648 303686
rect 301596 303622 301648 303628
rect 301504 230444 301556 230450
rect 301504 230386 301556 230392
rect 300216 230308 300268 230314
rect 300216 230250 300268 230256
rect 301608 224874 301636 303622
rect 301700 230178 301728 308926
rect 301976 306374 302004 319824
rect 302114 319818 302142 319892
rect 302194 319874 302246 319880
rect 302068 319790 302142 319818
rect 302068 317801 302096 319790
rect 302148 319728 302200 319734
rect 302298 319716 302326 320076
rect 302148 319670 302200 319676
rect 302252 319688 302326 319716
rect 302054 317792 302110 317801
rect 302054 317727 302110 317736
rect 302160 317626 302188 319670
rect 302252 318481 302280 319688
rect 302390 319648 302418 320076
rect 302482 319716 302510 320076
rect 302574 319818 302602 320076
rect 302666 319938 302694 320076
rect 303664 320104 303720 320113
rect 302836 320039 302892 320048
rect 302654 319932 302706 319938
rect 302654 319874 302706 319880
rect 302792 319932 302844 319938
rect 302792 319874 302844 319880
rect 302574 319790 302648 319818
rect 302482 319688 302556 319716
rect 302344 319620 302418 319648
rect 302344 318782 302372 319620
rect 302332 318776 302384 318782
rect 302332 318718 302384 318724
rect 302238 318472 302294 318481
rect 302238 318407 302294 318416
rect 302148 317620 302200 317626
rect 302148 317562 302200 317568
rect 302148 317484 302200 317490
rect 302148 317426 302200 317432
rect 302160 309126 302188 317426
rect 302528 315994 302556 319688
rect 302620 317529 302648 319790
rect 302700 319660 302752 319666
rect 302700 319602 302752 319608
rect 302606 317520 302662 317529
rect 302606 317455 302662 317464
rect 302712 316690 302740 319602
rect 302804 318209 302832 319874
rect 302942 319818 302970 320076
rect 302896 319790 302970 319818
rect 302790 318200 302846 318209
rect 302790 318135 302846 318144
rect 302620 316662 302740 316690
rect 302516 315988 302568 315994
rect 302516 315930 302568 315936
rect 302424 315784 302476 315790
rect 302424 315726 302476 315732
rect 302332 315716 302384 315722
rect 302332 315658 302384 315664
rect 302240 315444 302292 315450
rect 302240 315386 302292 315392
rect 302252 314770 302280 315386
rect 302240 314764 302292 314770
rect 302240 314706 302292 314712
rect 302148 309120 302200 309126
rect 302148 309062 302200 309068
rect 301792 306346 302004 306374
rect 301792 303482 301820 306346
rect 301780 303476 301832 303482
rect 301780 303418 301832 303424
rect 301688 230172 301740 230178
rect 301688 230114 301740 230120
rect 301792 226166 301820 303418
rect 301870 302832 301926 302841
rect 301870 302767 301926 302776
rect 301964 302796 302016 302802
rect 301884 228750 301912 302767
rect 301964 302738 302016 302744
rect 301976 235890 302004 302738
rect 302344 300558 302372 315658
rect 302436 304842 302464 315726
rect 302516 315444 302568 315450
rect 302516 315386 302568 315392
rect 302528 305862 302556 315386
rect 302620 309058 302648 316662
rect 302896 316146 302924 319790
rect 303034 319716 303062 320076
rect 303126 319818 303154 320076
rect 303218 319938 303246 320076
rect 303310 319938 303338 320076
rect 303206 319932 303258 319938
rect 303206 319874 303258 319880
rect 303298 319932 303350 319938
rect 303298 319874 303350 319880
rect 303402 319818 303430 320076
rect 303494 319938 303522 320076
rect 303482 319932 303534 319938
rect 303482 319874 303534 319880
rect 303586 319818 303614 320076
rect 305872 320104 305928 320113
rect 303664 320039 303720 320048
rect 303770 319920 303798 320076
rect 303126 319790 303200 319818
rect 302712 316118 302924 316146
rect 302988 319688 303062 319716
rect 302608 309052 302660 309058
rect 302608 308994 302660 309000
rect 302712 308446 302740 316118
rect 302792 316056 302844 316062
rect 302792 315998 302844 316004
rect 302804 309126 302832 315998
rect 302884 315988 302936 315994
rect 302884 315930 302936 315936
rect 302896 309874 302924 315930
rect 302988 315790 303016 319688
rect 303068 319592 303120 319598
rect 303068 319534 303120 319540
rect 302976 315784 303028 315790
rect 302976 315726 303028 315732
rect 303080 315722 303108 319534
rect 303172 317529 303200 319790
rect 303264 319790 303430 319818
rect 303540 319790 303614 319818
rect 303724 319892 303798 319920
rect 303158 317520 303214 317529
rect 303158 317455 303214 317464
rect 303068 315716 303120 315722
rect 303068 315658 303120 315664
rect 302884 309868 302936 309874
rect 302884 309810 302936 309816
rect 302792 309120 302844 309126
rect 302792 309062 302844 309068
rect 302700 308440 302752 308446
rect 302700 308382 302752 308388
rect 302516 305856 302568 305862
rect 302516 305798 302568 305804
rect 302424 304836 302476 304842
rect 302424 304778 302476 304784
rect 302436 304094 302464 304778
rect 302424 304088 302476 304094
rect 302424 304030 302476 304036
rect 302332 300552 302384 300558
rect 302332 300494 302384 300500
rect 302148 239420 302200 239426
rect 302148 239362 302200 239368
rect 302160 238241 302188 239362
rect 302146 238232 302202 238241
rect 302146 238167 302202 238176
rect 301964 235884 302016 235890
rect 301964 235826 302016 235832
rect 301872 228744 301924 228750
rect 301872 228686 301924 228692
rect 301780 226160 301832 226166
rect 301780 226102 301832 226108
rect 301596 224868 301648 224874
rect 301596 224810 301648 224816
rect 300124 224528 300176 224534
rect 300124 224470 300176 224476
rect 302896 224262 302924 309810
rect 302976 309120 303028 309126
rect 302976 309062 303028 309068
rect 302988 308922 303016 309062
rect 303160 309052 303212 309058
rect 303160 308994 303212 309000
rect 302976 308916 303028 308922
rect 302976 308858 303028 308864
rect 302988 306374 303016 308858
rect 303172 308854 303200 308994
rect 303160 308848 303212 308854
rect 303160 308790 303212 308796
rect 302988 306346 303108 306374
rect 302976 300552 303028 300558
rect 302976 300494 303028 300500
rect 302988 225758 303016 300494
rect 303080 234598 303108 306346
rect 303172 241126 303200 308790
rect 303264 298042 303292 319790
rect 303436 319728 303488 319734
rect 303436 319670 303488 319676
rect 303344 318028 303396 318034
rect 303344 317970 303396 317976
rect 303356 317801 303384 317970
rect 303342 317792 303398 317801
rect 303342 317727 303398 317736
rect 303344 317076 303396 317082
rect 303344 317018 303396 317024
rect 303356 316470 303384 317018
rect 303344 316464 303396 316470
rect 303344 316406 303396 316412
rect 303448 316062 303476 319670
rect 303436 316056 303488 316062
rect 303436 315998 303488 316004
rect 303540 315450 303568 319790
rect 303724 316402 303752 319892
rect 303862 319852 303890 320076
rect 303954 319920 303982 320076
rect 304138 319938 304166 320076
rect 304126 319932 304178 319938
rect 303954 319892 304028 319920
rect 303816 319824 303890 319852
rect 303816 317937 303844 319824
rect 303896 319728 303948 319734
rect 303896 319670 303948 319676
rect 303802 317928 303858 317937
rect 303802 317863 303858 317872
rect 303712 316396 303764 316402
rect 303712 316338 303764 316344
rect 303804 315920 303856 315926
rect 303804 315862 303856 315868
rect 303528 315444 303580 315450
rect 303528 315386 303580 315392
rect 303816 300286 303844 315862
rect 303908 302802 303936 319670
rect 304000 318034 304028 319892
rect 304126 319874 304178 319880
rect 304080 319796 304132 319802
rect 304080 319738 304132 319744
rect 303988 318028 304040 318034
rect 303988 317970 304040 317976
rect 303988 317756 304040 317762
rect 303988 317698 304040 317704
rect 304000 316130 304028 317698
rect 303988 316124 304040 316130
rect 303988 316066 304040 316072
rect 303988 315988 304040 315994
rect 303988 315930 304040 315936
rect 304000 307698 304028 315930
rect 304092 308650 304120 319738
rect 304230 319716 304258 320076
rect 304322 319870 304350 320076
rect 304310 319864 304362 319870
rect 304310 319806 304362 319812
rect 304414 319716 304442 320076
rect 304598 319920 304626 320076
rect 304690 319938 304718 320076
rect 304874 319954 304902 320076
rect 304184 319688 304258 319716
rect 304368 319688 304442 319716
rect 304552 319892 304626 319920
rect 304678 319932 304730 319938
rect 304184 316266 304212 319688
rect 304262 317792 304318 317801
rect 304262 317727 304318 317736
rect 304172 316260 304224 316266
rect 304172 316202 304224 316208
rect 304172 316056 304224 316062
rect 304172 315998 304224 316004
rect 304184 308990 304212 315998
rect 304172 308984 304224 308990
rect 304172 308926 304224 308932
rect 304080 308644 304132 308650
rect 304080 308586 304132 308592
rect 303988 307692 304040 307698
rect 303988 307634 304040 307640
rect 303896 302796 303948 302802
rect 303896 302738 303948 302744
rect 303804 300280 303856 300286
rect 303804 300222 303856 300228
rect 303252 298036 303304 298042
rect 303252 297978 303304 297984
rect 303264 289377 303292 297978
rect 303250 289368 303306 289377
rect 303250 289303 303306 289312
rect 303160 241120 303212 241126
rect 303160 241062 303212 241068
rect 303068 234592 303120 234598
rect 303068 234534 303120 234540
rect 302976 225752 303028 225758
rect 302976 225694 303028 225700
rect 302884 224256 302936 224262
rect 302884 224198 302936 224204
rect 303620 223032 303672 223038
rect 303620 222974 303672 222980
rect 303632 222902 303660 222974
rect 303620 222896 303672 222902
rect 303620 222838 303672 222844
rect 300860 160132 300912 160138
rect 300860 160074 300912 160080
rect 300872 16574 300900 160074
rect 302884 141636 302936 141642
rect 302884 141578 302936 141584
rect 299676 16546 300808 16574
rect 300872 16546 301544 16574
rect 299664 3596 299716 3602
rect 299664 3538 299716 3544
rect 299676 480 299704 3538
rect 300780 480 300808 16546
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 302896 3942 302924 141578
rect 303632 16574 303660 222838
rect 304276 219298 304304 317727
rect 304368 315994 304396 319688
rect 304552 319530 304580 319892
rect 304678 319874 304730 319880
rect 304828 319926 304902 319954
rect 304632 319796 304684 319802
rect 304632 319738 304684 319744
rect 304540 319524 304592 319530
rect 304540 319466 304592 319472
rect 304448 318708 304500 318714
rect 304448 318650 304500 318656
rect 304460 316606 304488 318650
rect 304448 316600 304500 316606
rect 304448 316542 304500 316548
rect 304448 316328 304500 316334
rect 304448 316270 304500 316276
rect 304460 316130 304488 316270
rect 304448 316124 304500 316130
rect 304448 316066 304500 316072
rect 304356 315988 304408 315994
rect 304356 315930 304408 315936
rect 304356 311500 304408 311506
rect 304356 311442 304408 311448
rect 304368 300150 304396 311442
rect 304448 308644 304500 308650
rect 304448 308586 304500 308592
rect 304356 300144 304408 300150
rect 304356 300086 304408 300092
rect 304368 223038 304396 300086
rect 304460 230382 304488 308586
rect 304538 307456 304594 307465
rect 304538 307391 304594 307400
rect 304552 233034 304580 307391
rect 304644 300626 304672 319738
rect 304724 319524 304776 319530
rect 304724 319466 304776 319472
rect 304736 317490 304764 319466
rect 304724 317484 304776 317490
rect 304724 317426 304776 317432
rect 304724 316668 304776 316674
rect 304724 316610 304776 316616
rect 304736 316402 304764 316610
rect 304724 316396 304776 316402
rect 304724 316338 304776 316344
rect 304724 316260 304776 316266
rect 304724 316202 304776 316208
rect 304632 300620 304684 300626
rect 304632 300562 304684 300568
rect 304644 234394 304672 300562
rect 304736 297906 304764 316202
rect 304828 316062 304856 319926
rect 304966 319818 304994 320076
rect 305058 319852 305086 320076
rect 305058 319824 305132 319852
rect 304920 319790 304994 319818
rect 304816 316056 304868 316062
rect 304816 315998 304868 316004
rect 304920 315926 304948 319790
rect 305104 319716 305132 319824
rect 305242 319784 305270 320076
rect 305426 319920 305454 320076
rect 305610 319920 305638 320076
rect 305702 319938 305730 320076
rect 305012 319688 305132 319716
rect 305196 319756 305270 319784
rect 305380 319892 305454 319920
rect 305564 319892 305638 319920
rect 305690 319932 305742 319938
rect 304908 315920 304960 315926
rect 304908 315862 304960 315868
rect 305012 314566 305040 319688
rect 305196 319648 305224 319756
rect 305104 319620 305224 319648
rect 305000 314560 305052 314566
rect 305000 314502 305052 314508
rect 305000 312452 305052 312458
rect 305000 312394 305052 312400
rect 305012 310418 305040 312394
rect 305104 310486 305132 319620
rect 305182 319560 305238 319569
rect 305182 319495 305238 319504
rect 305092 310480 305144 310486
rect 305092 310422 305144 310428
rect 305000 310412 305052 310418
rect 305000 310354 305052 310360
rect 305196 306338 305224 319495
rect 305380 318794 305408 319892
rect 305564 319444 305592 319892
rect 305690 319874 305742 319880
rect 305702 319784 305730 319874
rect 305794 319818 305822 320076
rect 306976 320104 307032 320113
rect 305872 320039 305928 320048
rect 305978 319920 306006 320076
rect 305932 319892 306006 319920
rect 305794 319790 305868 319818
rect 305288 318766 305408 318794
rect 305472 319416 305592 319444
rect 305656 319756 305730 319784
rect 305288 316470 305316 318766
rect 305276 316464 305328 316470
rect 305276 316406 305328 316412
rect 305276 316056 305328 316062
rect 305276 315998 305328 316004
rect 305288 308378 305316 315998
rect 305276 308372 305328 308378
rect 305276 308314 305328 308320
rect 305184 306332 305236 306338
rect 305184 306274 305236 306280
rect 305196 305046 305224 306274
rect 305184 305040 305236 305046
rect 305184 304982 305236 304988
rect 305366 302968 305422 302977
rect 305366 302903 305422 302912
rect 305380 302870 305408 302903
rect 305368 302864 305420 302870
rect 305368 302806 305420 302812
rect 304724 297900 304776 297906
rect 304724 297842 304776 297848
rect 304736 237998 304764 297842
rect 305380 296714 305408 302806
rect 305472 297838 305500 319416
rect 305550 319016 305606 319025
rect 305550 318951 305606 318960
rect 305564 316146 305592 318951
rect 305656 318510 305684 319756
rect 305734 319560 305790 319569
rect 305734 319495 305790 319504
rect 305644 318504 305696 318510
rect 305644 318446 305696 318452
rect 305564 316118 305684 316146
rect 305656 313206 305684 316118
rect 305644 313200 305696 313206
rect 305644 313142 305696 313148
rect 305656 312458 305684 313142
rect 305644 312452 305696 312458
rect 305644 312394 305696 312400
rect 305748 311894 305776 319495
rect 305564 311866 305776 311894
rect 305564 311250 305592 311866
rect 305840 311386 305868 319790
rect 305932 316062 305960 319892
rect 306070 319852 306098 320076
rect 306024 319824 306098 319852
rect 305920 316056 305972 316062
rect 305920 315998 305972 316004
rect 306024 311506 306052 319824
rect 306162 319818 306190 320076
rect 306346 319818 306374 320076
rect 306162 319790 306236 319818
rect 306104 319660 306156 319666
rect 306104 319602 306156 319608
rect 306116 319569 306144 319602
rect 306102 319560 306158 319569
rect 306102 319495 306158 319504
rect 306208 317801 306236 319790
rect 306300 319790 306374 319818
rect 306438 319818 306466 320076
rect 306530 319938 306558 320076
rect 306518 319932 306570 319938
rect 306518 319874 306570 319880
rect 306622 319818 306650 320076
rect 306438 319790 306512 319818
rect 306194 317792 306250 317801
rect 306194 317727 306250 317736
rect 306300 317529 306328 319790
rect 306484 319716 306512 319790
rect 306392 319688 306512 319716
rect 306576 319790 306650 319818
rect 306714 319818 306742 320076
rect 306806 319938 306834 320076
rect 306794 319932 306846 319938
rect 306794 319874 306846 319880
rect 306898 319818 306926 320076
rect 307344 320104 307400 320113
rect 306976 320039 307032 320048
rect 307024 319932 307076 319938
rect 307174 319920 307202 320076
rect 307024 319874 307076 319880
rect 307128 319892 307202 319920
rect 306714 319790 306788 319818
rect 306898 319790 306972 319818
rect 306392 318753 306420 319688
rect 306472 319524 306524 319530
rect 306472 319466 306524 319472
rect 306484 318918 306512 319466
rect 306472 318912 306524 318918
rect 306472 318854 306524 318860
rect 306378 318744 306434 318753
rect 306378 318679 306434 318688
rect 306392 317937 306420 318679
rect 306470 318472 306526 318481
rect 306470 318407 306526 318416
rect 306378 317928 306434 317937
rect 306378 317863 306434 317872
rect 306286 317520 306342 317529
rect 306286 317455 306342 317464
rect 306484 314770 306512 318407
rect 306472 314764 306524 314770
rect 306472 314706 306524 314712
rect 306378 314664 306434 314673
rect 306378 314599 306380 314608
rect 306432 314599 306434 314608
rect 306380 314570 306432 314576
rect 306012 311500 306064 311506
rect 306012 311442 306064 311448
rect 305840 311358 306052 311386
rect 305564 311222 305960 311250
rect 305828 308372 305880 308378
rect 305828 308314 305880 308320
rect 305644 305040 305696 305046
rect 305644 304982 305696 304988
rect 305460 297832 305512 297838
rect 305460 297774 305512 297780
rect 305196 296686 305408 296714
rect 304724 237992 304776 237998
rect 304724 237934 304776 237940
rect 304632 234388 304684 234394
rect 304632 234330 304684 234336
rect 304540 233028 304592 233034
rect 304540 232970 304592 232976
rect 305196 231538 305224 296686
rect 305656 234530 305684 304982
rect 305736 300212 305788 300218
rect 305736 300154 305788 300160
rect 305644 234524 305696 234530
rect 305644 234466 305696 234472
rect 305184 231532 305236 231538
rect 305184 231474 305236 231480
rect 305644 230444 305696 230450
rect 305644 230386 305696 230392
rect 304448 230376 304500 230382
rect 304448 230318 304500 230324
rect 305656 230246 305684 230386
rect 305644 230240 305696 230246
rect 305644 230182 305696 230188
rect 304356 223032 304408 223038
rect 304356 222974 304408 222980
rect 304264 219292 304316 219298
rect 304264 219234 304316 219240
rect 305000 176724 305052 176730
rect 305000 176666 305052 176672
rect 305012 16574 305040 176666
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 302884 3936 302936 3942
rect 302884 3878 302936 3884
rect 303160 3732 303212 3738
rect 303160 3674 303212 3680
rect 303172 480 303200 3674
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 305656 3874 305684 230182
rect 305748 226030 305776 300154
rect 305840 239494 305868 308314
rect 305932 301442 305960 311222
rect 305920 301436 305972 301442
rect 305920 301378 305972 301384
rect 305828 239488 305880 239494
rect 305828 239430 305880 239436
rect 305932 238950 305960 301378
rect 306024 300694 306052 311358
rect 306012 300688 306064 300694
rect 306012 300630 306064 300636
rect 306576 300218 306604 319790
rect 306760 319682 306788 319790
rect 306760 319654 306880 319682
rect 306746 319560 306802 319569
rect 306746 319495 306802 319504
rect 306654 319424 306710 319433
rect 306654 319359 306710 319368
rect 306668 318782 306696 319359
rect 306656 318776 306708 318782
rect 306656 318718 306708 318724
rect 306656 316260 306708 316266
rect 306656 316202 306708 316208
rect 306668 303385 306696 316202
rect 306760 305454 306788 319495
rect 306852 317529 306880 319654
rect 306838 317520 306894 317529
rect 306838 317455 306894 317464
rect 306840 316056 306892 316062
rect 306840 315998 306892 316004
rect 306852 306377 306880 315998
rect 306838 306368 306894 306377
rect 306838 306303 306894 306312
rect 306748 305448 306800 305454
rect 306748 305390 306800 305396
rect 306654 303376 306710 303385
rect 306654 303311 306710 303320
rect 306668 302297 306696 303311
rect 306654 302288 306710 302297
rect 306654 302223 306710 302232
rect 306944 300354 306972 319790
rect 307036 317150 307064 319874
rect 307128 319784 307156 319892
rect 307266 319852 307294 320076
rect 308080 320104 308136 320113
rect 307344 320039 307400 320048
rect 307266 319824 307340 319852
rect 307128 319756 307248 319784
rect 307116 319592 307168 319598
rect 307116 319534 307168 319540
rect 307024 317144 307076 317150
rect 307024 317086 307076 317092
rect 307128 316266 307156 319534
rect 307116 316260 307168 316266
rect 307116 316202 307168 316208
rect 307116 315988 307168 315994
rect 307116 315930 307168 315936
rect 307024 315444 307076 315450
rect 307024 315386 307076 315392
rect 307036 314702 307064 315386
rect 307024 314696 307076 314702
rect 307024 314638 307076 314644
rect 307036 304094 307064 314638
rect 307128 305017 307156 315930
rect 307220 311250 307248 319756
rect 307312 319598 307340 319824
rect 307450 319818 307478 320076
rect 307726 319954 307754 320076
rect 307404 319790 307478 319818
rect 307588 319926 307754 319954
rect 307300 319592 307352 319598
rect 307300 319534 307352 319540
rect 307298 319424 307354 319433
rect 307298 319359 307354 319368
rect 307312 316062 307340 319359
rect 307300 316056 307352 316062
rect 307300 315998 307352 316004
rect 307404 315994 307432 319790
rect 307484 319728 307536 319734
rect 307484 319670 307536 319676
rect 307496 317762 307524 319670
rect 307484 317756 307536 317762
rect 307484 317698 307536 317704
rect 307588 317608 307616 319926
rect 307818 319852 307846 320076
rect 307772 319824 307846 319852
rect 307668 319592 307720 319598
rect 307668 319534 307720 319540
rect 307680 318714 307708 319534
rect 307668 318708 307720 318714
rect 307668 318650 307720 318656
rect 307496 317580 307616 317608
rect 307392 315988 307444 315994
rect 307392 315930 307444 315936
rect 307496 315450 307524 317580
rect 307772 317529 307800 319824
rect 307910 319784 307938 320076
rect 308002 319818 308030 320076
rect 309828 320104 309884 320113
rect 308080 320039 308136 320048
rect 308186 319852 308214 320076
rect 308140 319824 308214 319852
rect 308002 319790 308076 319818
rect 307864 319756 307938 319784
rect 307864 319598 307892 319756
rect 307944 319660 307996 319666
rect 307944 319602 307996 319608
rect 307852 319592 307904 319598
rect 307956 319569 307984 319602
rect 307852 319534 307904 319540
rect 307942 319560 307998 319569
rect 307942 319495 307998 319504
rect 307942 319424 307998 319433
rect 307942 319359 307998 319368
rect 307852 318912 307904 318918
rect 307852 318854 307904 318860
rect 307758 317520 307814 317529
rect 307576 317484 307628 317490
rect 307758 317455 307814 317464
rect 307576 317426 307628 317432
rect 307484 315444 307536 315450
rect 307484 315386 307536 315392
rect 307220 311222 307432 311250
rect 307298 306368 307354 306377
rect 307404 306374 307432 311222
rect 307404 306346 307524 306374
rect 307298 306303 307354 306312
rect 307114 305008 307170 305017
rect 307114 304943 307170 304952
rect 307024 304088 307076 304094
rect 307024 304030 307076 304036
rect 307114 302288 307170 302297
rect 307114 302223 307170 302232
rect 306932 300348 306984 300354
rect 306932 300290 306984 300296
rect 306564 300212 306616 300218
rect 306564 300154 306616 300160
rect 306104 297832 306156 297838
rect 306104 297774 306156 297780
rect 306116 289105 306144 297774
rect 306944 296714 306972 300290
rect 306944 296686 307064 296714
rect 306102 289096 306158 289105
rect 306102 289031 306158 289040
rect 306012 288448 306064 288454
rect 306012 288390 306064 288396
rect 305920 238944 305972 238950
rect 305920 238886 305972 238892
rect 306024 230450 306052 288390
rect 306012 230444 306064 230450
rect 306012 230386 306064 230392
rect 307036 226098 307064 296686
rect 307024 226092 307076 226098
rect 307024 226034 307076 226040
rect 305736 226024 305788 226030
rect 305736 225966 305788 225972
rect 305644 3868 305696 3874
rect 305644 3810 305696 3816
rect 305748 3534 305776 225966
rect 306748 3936 306800 3942
rect 306748 3878 306800 3884
rect 305736 3528 305788 3534
rect 305736 3470 305788 3476
rect 306760 480 306788 3878
rect 307036 3058 307064 226034
rect 307128 220726 307156 302223
rect 307208 301912 307260 301918
rect 307208 301854 307260 301860
rect 307220 300082 307248 301854
rect 307208 300076 307260 300082
rect 307208 300018 307260 300024
rect 307208 292528 307260 292534
rect 307208 292470 307260 292476
rect 307220 221746 307248 292470
rect 307312 241194 307340 306303
rect 307392 305652 307444 305658
rect 307392 305594 307444 305600
rect 307404 305454 307432 305594
rect 307392 305448 307444 305454
rect 307392 305390 307444 305396
rect 307404 247722 307432 305390
rect 307496 300762 307524 306346
rect 307484 300756 307536 300762
rect 307484 300698 307536 300704
rect 307496 288454 307524 300698
rect 307588 297129 307616 317426
rect 307864 311894 307892 318854
rect 307956 317490 307984 319359
rect 307944 317484 307996 317490
rect 307944 317426 307996 317432
rect 307864 311866 307984 311894
rect 307666 305008 307722 305017
rect 307666 304943 307722 304952
rect 307680 301918 307708 304943
rect 307758 303648 307814 303657
rect 307758 303583 307814 303592
rect 307668 301912 307720 301918
rect 307668 301854 307720 301860
rect 307668 300484 307720 300490
rect 307668 300426 307720 300432
rect 307680 300218 307708 300426
rect 307772 300218 307800 303583
rect 307668 300212 307720 300218
rect 307668 300154 307720 300160
rect 307760 300212 307812 300218
rect 307760 300154 307812 300160
rect 307668 300076 307720 300082
rect 307668 300018 307720 300024
rect 307574 297120 307630 297129
rect 307574 297055 307630 297064
rect 307484 288448 307536 288454
rect 307484 288390 307536 288396
rect 307484 249756 307536 249762
rect 307484 249698 307536 249704
rect 307392 247716 307444 247722
rect 307392 247658 307444 247664
rect 307300 241188 307352 241194
rect 307300 241130 307352 241136
rect 307208 221740 307260 221746
rect 307208 221682 307260 221688
rect 307116 220720 307168 220726
rect 307116 220662 307168 220668
rect 307496 216578 307524 249698
rect 307680 236706 307708 300018
rect 307668 236700 307720 236706
rect 307668 236642 307720 236648
rect 307116 216572 307168 216578
rect 307116 216514 307168 216520
rect 307484 216572 307536 216578
rect 307484 216514 307536 216520
rect 307128 3806 307156 216514
rect 307208 152652 307260 152658
rect 307208 152594 307260 152600
rect 307116 3800 307168 3806
rect 307116 3742 307168 3748
rect 307220 3194 307248 152594
rect 307772 3482 307800 300154
rect 307956 297974 307984 311866
rect 308048 300830 308076 319790
rect 308140 319682 308168 319824
rect 308278 319784 308306 320076
rect 308370 319920 308398 320076
rect 308554 319920 308582 320076
rect 308370 319892 308490 319920
rect 308554 319892 308628 319920
rect 308462 319852 308490 319892
rect 308462 319824 308536 319852
rect 308278 319756 308444 319784
rect 308140 319654 308352 319682
rect 308126 319560 308182 319569
rect 308126 319495 308182 319504
rect 308140 306202 308168 319495
rect 308218 319016 308274 319025
rect 308218 318951 308274 318960
rect 308232 306270 308260 318951
rect 308324 318345 308352 319654
rect 308310 318336 308366 318345
rect 308310 318271 308366 318280
rect 308312 316056 308364 316062
rect 308312 315998 308364 316004
rect 308324 311030 308352 315998
rect 308416 314634 308444 319756
rect 308508 318918 308536 319824
rect 308496 318912 308548 318918
rect 308496 318854 308548 318860
rect 308494 318744 308550 318753
rect 308494 318679 308550 318688
rect 308404 314628 308456 314634
rect 308404 314570 308456 314576
rect 308312 311024 308364 311030
rect 308312 310966 308364 310972
rect 308220 306264 308272 306270
rect 308220 306206 308272 306212
rect 308128 306196 308180 306202
rect 308128 306138 308180 306144
rect 308140 305998 308168 306138
rect 308128 305992 308180 305998
rect 308128 305934 308180 305940
rect 308232 305046 308260 306206
rect 308220 305040 308272 305046
rect 308220 304982 308272 304988
rect 308036 300824 308088 300830
rect 308036 300766 308088 300772
rect 307944 297968 307996 297974
rect 307944 297910 307996 297916
rect 308416 217326 308444 314570
rect 308508 314090 308536 318679
rect 308600 315994 308628 319892
rect 308830 319852 308858 320076
rect 308922 319938 308950 320076
rect 308910 319932 308962 319938
rect 308910 319874 308962 319880
rect 308784 319824 308858 319852
rect 308680 319592 308732 319598
rect 308680 319534 308732 319540
rect 308588 315988 308640 315994
rect 308588 315930 308640 315936
rect 308496 314084 308548 314090
rect 308496 314026 308548 314032
rect 308692 306105 308720 319534
rect 308784 315178 308812 319824
rect 309014 319784 309042 320076
rect 308968 319756 309042 319784
rect 308864 319728 308916 319734
rect 308864 319670 308916 319676
rect 308876 317801 308904 319670
rect 308968 319598 308996 319756
rect 309106 319716 309134 320076
rect 309198 319784 309226 320076
rect 309290 319938 309318 320076
rect 309278 319932 309330 319938
rect 309278 319874 309330 319880
rect 309382 319818 309410 320076
rect 309566 319954 309594 320076
rect 309750 319954 309778 320076
rect 310288 320104 310344 320113
rect 309828 320039 309884 320048
rect 309566 319926 309640 319954
rect 309336 319790 309410 319818
rect 309508 319864 309560 319870
rect 309508 319806 309560 319812
rect 309198 319756 309272 319784
rect 309060 319688 309134 319716
rect 308956 319592 309008 319598
rect 308956 319534 309008 319540
rect 308956 319048 309008 319054
rect 308956 318990 309008 318996
rect 308968 318918 308996 318990
rect 308956 318912 309008 318918
rect 308956 318854 309008 318860
rect 308862 317792 308918 317801
rect 308862 317727 308918 317736
rect 309060 316062 309088 319688
rect 309244 319648 309272 319756
rect 309152 319620 309272 319648
rect 309152 318510 309180 319620
rect 309230 319560 309286 319569
rect 309230 319495 309286 319504
rect 309140 318504 309192 318510
rect 309140 318446 309192 318452
rect 309140 317212 309192 317218
rect 309140 317154 309192 317160
rect 309152 317014 309180 317154
rect 309140 317008 309192 317014
rect 309140 316950 309192 316956
rect 309048 316056 309100 316062
rect 309048 315998 309100 316004
rect 308864 315988 308916 315994
rect 308864 315930 308916 315936
rect 308772 315172 308824 315178
rect 308772 315114 308824 315120
rect 308678 306096 308734 306105
rect 308678 306031 308734 306040
rect 308588 305040 308640 305046
rect 308588 304982 308640 304988
rect 308496 297968 308548 297974
rect 308496 297910 308548 297916
rect 308508 297770 308536 297910
rect 308496 297764 308548 297770
rect 308496 297706 308548 297712
rect 308508 227361 308536 297706
rect 308600 241262 308628 304982
rect 308680 300824 308732 300830
rect 308680 300766 308732 300772
rect 308692 300082 308720 300766
rect 308680 300076 308732 300082
rect 308680 300018 308732 300024
rect 308692 249762 308720 300018
rect 308876 291990 308904 315930
rect 309140 315784 309192 315790
rect 309140 315726 309192 315732
rect 309046 298072 309102 298081
rect 309046 298007 309102 298016
rect 309060 297974 309088 298007
rect 309048 297968 309100 297974
rect 309048 297910 309100 297916
rect 309048 297696 309100 297702
rect 309046 297664 309048 297673
rect 309100 297664 309102 297673
rect 308956 297628 309008 297634
rect 309046 297599 309102 297608
rect 308956 297570 309008 297576
rect 308968 297129 308996 297570
rect 308954 297120 309010 297129
rect 308954 297055 309010 297064
rect 308864 291984 308916 291990
rect 308864 291926 308916 291932
rect 309152 291922 309180 315726
rect 309244 301782 309272 319495
rect 309232 301776 309284 301782
rect 309232 301718 309284 301724
rect 309336 301714 309364 319790
rect 309416 319728 309468 319734
rect 309416 319670 309468 319676
rect 309428 317218 309456 319670
rect 309416 317212 309468 317218
rect 309416 317154 309468 317160
rect 309416 316940 309468 316946
rect 309416 316882 309468 316888
rect 309428 316810 309456 316882
rect 309416 316804 309468 316810
rect 309416 316746 309468 316752
rect 309416 315988 309468 315994
rect 309416 315930 309468 315936
rect 309324 301708 309376 301714
rect 309324 301650 309376 301656
rect 309428 301646 309456 315930
rect 309520 305969 309548 319806
rect 309612 316810 309640 319926
rect 309704 319926 309778 319954
rect 309704 319433 309732 319926
rect 309934 319818 309962 320076
rect 309888 319790 309962 319818
rect 310026 319818 310054 320076
rect 310118 319938 310146 320076
rect 310106 319932 310158 319938
rect 310210 319920 310238 320076
rect 311668 320104 311724 320113
rect 310288 320039 310344 320048
rect 310210 319892 310284 319920
rect 310106 319874 310158 319880
rect 310026 319790 310100 319818
rect 309782 319560 309838 319569
rect 309782 319495 309838 319504
rect 309690 319424 309746 319433
rect 309690 319359 309746 319368
rect 309692 319048 309744 319054
rect 309692 318990 309744 318996
rect 309704 318889 309732 318990
rect 309690 318880 309746 318889
rect 309690 318815 309746 318824
rect 309796 317529 309824 319495
rect 309782 317520 309838 317529
rect 309782 317455 309838 317464
rect 309600 316804 309652 316810
rect 309600 316746 309652 316752
rect 309600 315920 309652 315926
rect 309600 315862 309652 315868
rect 309612 305998 309640 315862
rect 309888 313274 309916 319790
rect 310072 318794 310100 319790
rect 309980 318766 310100 318794
rect 309980 317529 310008 318766
rect 309966 317520 310022 317529
rect 309966 317455 310022 317464
rect 310256 315790 310284 319892
rect 310394 319818 310422 320076
rect 310348 319790 310422 319818
rect 310348 315926 310376 319790
rect 310486 319716 310514 320076
rect 310440 319688 310514 319716
rect 310578 319716 310606 320076
rect 310670 319870 310698 320076
rect 310762 319938 310790 320076
rect 310750 319932 310802 319938
rect 310854 319920 310882 320076
rect 310854 319892 310928 319920
rect 310750 319874 310802 319880
rect 310658 319864 310710 319870
rect 310658 319806 310710 319812
rect 310796 319796 310848 319802
rect 310796 319738 310848 319744
rect 310704 319728 310756 319734
rect 310578 319688 310652 319716
rect 310440 315994 310468 319688
rect 310428 315988 310480 315994
rect 310428 315930 310480 315936
rect 310624 315926 310652 319688
rect 310704 319670 310756 319676
rect 310716 318782 310744 319670
rect 310704 318776 310756 318782
rect 310704 318718 310756 318724
rect 310704 316056 310756 316062
rect 310704 315998 310756 316004
rect 310336 315920 310388 315926
rect 310336 315862 310388 315868
rect 310612 315920 310664 315926
rect 310612 315862 310664 315868
rect 310520 315852 310572 315858
rect 310520 315794 310572 315800
rect 310244 315784 310296 315790
rect 310058 315752 310114 315761
rect 310244 315726 310296 315732
rect 310058 315687 310114 315696
rect 309876 313268 309928 313274
rect 309876 313210 309928 313216
rect 309782 313168 309838 313177
rect 309782 313103 309838 313112
rect 309692 313064 309744 313070
rect 309692 313006 309744 313012
rect 309704 312361 309732 313006
rect 309690 312352 309746 312361
rect 309690 312287 309746 312296
rect 309796 306134 309824 313103
rect 310072 313070 310100 315687
rect 310532 315625 310560 315794
rect 310518 315616 310574 315625
rect 310518 315551 310574 315560
rect 310520 313880 310572 313886
rect 310520 313822 310572 313828
rect 310428 313268 310480 313274
rect 310428 313210 310480 313216
rect 310060 313064 310112 313070
rect 310060 313006 310112 313012
rect 310440 312254 310468 313210
rect 310532 312905 310560 313822
rect 310518 312896 310574 312905
rect 310518 312831 310574 312840
rect 310428 312248 310480 312254
rect 310428 312190 310480 312196
rect 309784 306128 309836 306134
rect 309784 306070 309836 306076
rect 309600 305992 309652 305998
rect 309506 305960 309562 305969
rect 309600 305934 309652 305940
rect 309506 305895 309562 305904
rect 309612 303090 309640 305934
rect 309612 303062 309916 303090
rect 309784 301980 309836 301986
rect 309784 301922 309836 301928
rect 309796 301714 309824 301922
rect 309784 301708 309836 301714
rect 309784 301650 309836 301656
rect 309416 301640 309468 301646
rect 309416 301582 309468 301588
rect 309140 291916 309192 291922
rect 309140 291858 309192 291864
rect 308680 249756 308732 249762
rect 308680 249698 308732 249704
rect 308588 241256 308640 241262
rect 308588 241198 308640 241204
rect 308494 227352 308550 227361
rect 308494 227287 308550 227296
rect 309796 220114 309824 301650
rect 309888 242350 309916 303062
rect 310152 301776 310204 301782
rect 310204 301724 310376 301730
rect 310152 301718 310376 301724
rect 310164 301702 310376 301718
rect 310164 299266 310192 301702
rect 310348 301646 310376 301702
rect 310244 301640 310296 301646
rect 310244 301582 310296 301588
rect 310336 301640 310388 301646
rect 310336 301582 310388 301588
rect 310152 299260 310204 299266
rect 310152 299202 310204 299208
rect 310060 299192 310112 299198
rect 310060 299134 310112 299140
rect 310072 298217 310100 299134
rect 310058 298208 310114 298217
rect 310058 298143 310114 298152
rect 310256 259486 310284 301582
rect 310336 299464 310388 299470
rect 310334 299432 310336 299441
rect 310388 299432 310390 299441
rect 310334 299367 310390 299376
rect 310336 299260 310388 299266
rect 310336 299202 310388 299208
rect 310244 259480 310296 259486
rect 310244 259422 310296 259428
rect 310256 258074 310284 259422
rect 309980 258046 310284 258074
rect 309876 242344 309928 242350
rect 309876 242286 309928 242292
rect 309980 225962 310008 258046
rect 310348 252754 310376 299202
rect 310336 252748 310388 252754
rect 310336 252690 310388 252696
rect 310060 245676 310112 245682
rect 310060 245618 310112 245624
rect 309968 225956 310020 225962
rect 309968 225898 310020 225904
rect 310072 225894 310100 245618
rect 310348 238754 310376 252690
rect 310440 245886 310468 312190
rect 310716 307698 310744 315998
rect 310808 315994 310836 319738
rect 310900 319666 310928 319892
rect 311038 319784 311066 320076
rect 311222 319920 311250 320076
rect 311176 319892 311250 319920
rect 311038 319756 311112 319784
rect 310888 319660 310940 319666
rect 310888 319602 310940 319608
rect 310978 319424 311034 319433
rect 310978 319359 311034 319368
rect 310888 318844 310940 318850
rect 310888 318786 310940 318792
rect 310796 315988 310848 315994
rect 310796 315930 310848 315936
rect 310796 315852 310848 315858
rect 310796 315794 310848 315800
rect 310808 309058 310836 315794
rect 310900 311166 310928 318786
rect 310992 318782 311020 319359
rect 310980 318776 311032 318782
rect 310980 318718 311032 318724
rect 311084 318458 311112 319756
rect 311176 318646 311204 319892
rect 311314 319818 311342 320076
rect 311268 319790 311342 319818
rect 311406 319818 311434 320076
rect 311590 319818 311618 320076
rect 312128 320104 312184 320113
rect 311668 320039 311724 320048
rect 311774 319954 311802 320076
rect 311406 319790 311480 319818
rect 311268 318850 311296 319790
rect 311348 319660 311400 319666
rect 311348 319602 311400 319608
rect 311256 318844 311308 318850
rect 311256 318786 311308 318792
rect 311164 318640 311216 318646
rect 311164 318582 311216 318588
rect 311084 318430 311204 318458
rect 311072 315988 311124 315994
rect 311072 315930 311124 315936
rect 310888 311160 310940 311166
rect 310888 311102 310940 311108
rect 311084 311098 311112 315930
rect 311176 315625 311204 318430
rect 311256 317756 311308 317762
rect 311256 317698 311308 317704
rect 311162 315616 311218 315625
rect 311162 315551 311218 315560
rect 311268 314090 311296 317698
rect 311256 314084 311308 314090
rect 311256 314026 311308 314032
rect 311360 313886 311388 319602
rect 311452 316266 311480 319790
rect 311544 319790 311618 319818
rect 311728 319926 311802 319954
rect 311440 316260 311492 316266
rect 311440 316202 311492 316208
rect 311348 313880 311400 313886
rect 311348 313822 311400 313828
rect 311544 311506 311572 319790
rect 311624 316260 311676 316266
rect 311624 316202 311676 316208
rect 311532 311500 311584 311506
rect 311532 311442 311584 311448
rect 311256 311160 311308 311166
rect 311256 311102 311308 311108
rect 311072 311092 311124 311098
rect 311072 311034 311124 311040
rect 311268 310962 311296 311102
rect 311256 310956 311308 310962
rect 311256 310898 311308 310904
rect 310980 309596 311032 309602
rect 310980 309538 311032 309544
rect 310796 309052 310848 309058
rect 310796 308994 310848 309000
rect 310704 307692 310756 307698
rect 310704 307634 310756 307640
rect 310992 306374 311020 309538
rect 310992 306346 311204 306374
rect 310520 291916 310572 291922
rect 310520 291858 310572 291864
rect 310428 245880 310480 245886
rect 310428 245822 310480 245828
rect 310440 245682 310468 245822
rect 310428 245676 310480 245682
rect 310428 245618 310480 245624
rect 310164 238726 310376 238754
rect 310164 236434 310192 238726
rect 310152 236428 310204 236434
rect 310152 236370 310204 236376
rect 310532 228721 310560 291858
rect 310518 228712 310574 228721
rect 310518 228647 310574 228656
rect 310060 225888 310112 225894
rect 310060 225830 310112 225836
rect 311176 223106 311204 306346
rect 311268 223174 311296 310898
rect 311544 309602 311572 311442
rect 311532 309596 311584 309602
rect 311532 309538 311584 309544
rect 311348 309052 311400 309058
rect 311348 308994 311400 309000
rect 311360 224913 311388 308994
rect 311440 307692 311492 307698
rect 311440 307634 311492 307640
rect 311452 307018 311480 307634
rect 311440 307012 311492 307018
rect 311440 306954 311492 306960
rect 311452 239562 311480 306954
rect 311636 298897 311664 316202
rect 311728 316062 311756 319926
rect 311866 319818 311894 320076
rect 311958 319870 311986 320076
rect 311820 319790 311894 319818
rect 311946 319864 311998 319870
rect 311946 319806 311998 319812
rect 311716 316056 311768 316062
rect 311716 315998 311768 316004
rect 311716 315920 311768 315926
rect 311716 315862 311768 315868
rect 311728 299062 311756 315862
rect 311820 315858 311848 319790
rect 312050 319784 312078 320076
rect 312772 320104 312828 320113
rect 312128 320039 312184 320048
rect 312234 319852 312262 320076
rect 312326 319938 312354 320076
rect 312314 319932 312366 319938
rect 312314 319874 312366 319880
rect 312188 319824 312262 319852
rect 312050 319756 312124 319784
rect 311900 319660 311952 319666
rect 312096 319648 312124 319756
rect 311900 319602 311952 319608
rect 312050 319620 312124 319648
rect 311912 317529 311940 319602
rect 312050 319580 312078 319620
rect 312004 319552 312078 319580
rect 311898 317520 311954 317529
rect 311898 317455 311954 317464
rect 312004 316878 312032 319552
rect 312082 319016 312138 319025
rect 312082 318951 312138 318960
rect 311992 316872 312044 316878
rect 311992 316814 312044 316820
rect 311992 316192 312044 316198
rect 311992 316134 312044 316140
rect 311808 315852 311860 315858
rect 311808 315794 311860 315800
rect 312004 314498 312032 316134
rect 312096 316062 312124 318951
rect 312188 316198 312216 319824
rect 312418 319818 312446 320076
rect 312418 319790 312492 319818
rect 312464 319784 312492 319790
rect 312694 319784 312722 320076
rect 313876 320104 313932 320113
rect 312772 320039 312828 320048
rect 312878 319784 312906 320076
rect 312464 319756 312584 319784
rect 312694 319756 312768 319784
rect 312452 319660 312504 319666
rect 312452 319602 312504 319608
rect 312266 319424 312322 319433
rect 312266 319359 312322 319368
rect 312176 316192 312228 316198
rect 312176 316134 312228 316140
rect 312084 316056 312136 316062
rect 312084 315998 312136 316004
rect 312176 315988 312228 315994
rect 312176 315930 312228 315936
rect 312084 315852 312136 315858
rect 312084 315794 312136 315800
rect 311992 314492 312044 314498
rect 311992 314434 312044 314440
rect 311808 311092 311860 311098
rect 311808 311034 311860 311040
rect 311716 299056 311768 299062
rect 311716 298998 311768 299004
rect 311622 298888 311678 298897
rect 311622 298823 311678 298832
rect 311728 287745 311756 298998
rect 311714 287736 311770 287745
rect 311714 287671 311770 287680
rect 311820 258074 311848 311034
rect 312096 301714 312124 315794
rect 312188 306241 312216 315930
rect 312280 307329 312308 319359
rect 312360 315920 312412 315926
rect 312360 315862 312412 315868
rect 312372 307465 312400 315862
rect 312464 315450 312492 319602
rect 312556 315858 312584 319756
rect 312740 316742 312768 319756
rect 312832 319756 312906 319784
rect 312970 319784 312998 320076
rect 313062 319938 313090 320076
rect 313050 319932 313102 319938
rect 313050 319874 313102 319880
rect 313154 319784 313182 320076
rect 312970 319756 313044 319784
rect 312728 316736 312780 316742
rect 312728 316678 312780 316684
rect 312832 315994 312860 319756
rect 312912 319660 312964 319666
rect 312912 319602 312964 319608
rect 312924 317801 312952 319602
rect 312910 317792 312966 317801
rect 312910 317727 312966 317736
rect 313016 316334 313044 319756
rect 313108 319756 313182 319784
rect 313004 316328 313056 316334
rect 313004 316270 313056 316276
rect 313004 316192 313056 316198
rect 313004 316134 313056 316140
rect 312912 316056 312964 316062
rect 312912 315998 312964 316004
rect 312820 315988 312872 315994
rect 312820 315930 312872 315936
rect 312544 315852 312596 315858
rect 312544 315794 312596 315800
rect 312452 315444 312504 315450
rect 312452 315386 312504 315392
rect 312450 314664 312506 314673
rect 312450 314599 312506 314608
rect 312464 313342 312492 314599
rect 312818 314528 312874 314537
rect 312818 314463 312874 314472
rect 312452 313336 312504 313342
rect 312452 313278 312504 313284
rect 312542 313168 312598 313177
rect 312542 313103 312598 313112
rect 312358 307456 312414 307465
rect 312358 307391 312414 307400
rect 312266 307320 312322 307329
rect 312266 307255 312322 307264
rect 312174 306232 312230 306241
rect 312174 306167 312230 306176
rect 312084 301708 312136 301714
rect 312084 301650 312136 301656
rect 312360 301708 312412 301714
rect 312360 301650 312412 301656
rect 311544 258046 311848 258074
rect 311544 254046 311572 258046
rect 311532 254040 311584 254046
rect 311532 253982 311584 253988
rect 311440 239556 311492 239562
rect 311440 239498 311492 239504
rect 311544 233753 311572 253982
rect 312372 244458 312400 301650
rect 312452 262880 312504 262886
rect 312452 262822 312504 262828
rect 312360 244452 312412 244458
rect 312360 244394 312412 244400
rect 312464 238678 312492 262822
rect 312452 238672 312504 238678
rect 312452 238614 312504 238620
rect 311530 233744 311586 233753
rect 311530 233679 311586 233688
rect 312556 226001 312584 313103
rect 312832 312662 312860 314463
rect 312820 312656 312872 312662
rect 312820 312598 312872 312604
rect 312832 312186 312860 312598
rect 312820 312180 312872 312186
rect 312820 312122 312872 312128
rect 312726 307320 312782 307329
rect 312726 307255 312782 307264
rect 312636 300756 312688 300762
rect 312636 300698 312688 300704
rect 312648 234161 312676 300698
rect 312740 245002 312768 307255
rect 312924 302054 312952 315998
rect 312912 302048 312964 302054
rect 312912 301990 312964 301996
rect 312924 248538 312952 301990
rect 313016 300762 313044 316134
rect 313108 315926 313136 319756
rect 313246 319682 313274 320076
rect 313338 319784 313366 320076
rect 313430 319954 313458 320076
rect 313430 319926 313504 319954
rect 313338 319756 313412 319784
rect 313200 319654 313274 319682
rect 313200 317490 313228 319654
rect 313188 317484 313240 317490
rect 313188 317426 313240 317432
rect 313188 316328 313240 316334
rect 313188 316270 313240 316276
rect 313096 315920 313148 315926
rect 313096 315862 313148 315868
rect 313200 314974 313228 316270
rect 313384 316062 313412 319756
rect 313476 318238 313504 319926
rect 313614 319818 313642 320076
rect 313706 319954 313734 320076
rect 313876 320039 313932 320048
rect 313706 319926 313780 319954
rect 313752 319920 313780 319926
rect 313752 319892 313826 319920
rect 313798 319818 313826 319892
rect 313614 319790 313688 319818
rect 313556 319728 313608 319734
rect 313556 319670 313608 319676
rect 313464 318232 313516 318238
rect 313464 318174 313516 318180
rect 313568 316282 313596 319670
rect 313660 318753 313688 319790
rect 313752 319790 313826 319818
rect 313646 318744 313702 318753
rect 313646 318679 313702 318688
rect 313476 316254 313596 316282
rect 313372 316056 313424 316062
rect 313372 315998 313424 316004
rect 313188 314968 313240 314974
rect 313188 314910 313240 314916
rect 313094 314664 313150 314673
rect 313094 314599 313150 314608
rect 313108 313138 313136 314599
rect 313096 313132 313148 313138
rect 313096 313074 313148 313080
rect 313108 312730 313136 313074
rect 313096 312724 313148 312730
rect 313096 312666 313148 312672
rect 313200 311894 313228 314910
rect 313108 311866 313228 311894
rect 313004 300756 313056 300762
rect 313004 300698 313056 300704
rect 313108 257378 313136 311866
rect 313476 307873 313504 316254
rect 313556 316192 313608 316198
rect 313556 316134 313608 316140
rect 313568 310282 313596 316134
rect 313660 315314 313688 318679
rect 313752 316266 313780 319790
rect 313982 319784 314010 320076
rect 313936 319756 314010 319784
rect 314074 319784 314102 320076
rect 314258 319938 314286 320076
rect 314246 319932 314298 319938
rect 314246 319874 314298 319880
rect 314350 319784 314378 320076
rect 314074 319756 314148 319784
rect 313832 319728 313884 319734
rect 313832 319670 313884 319676
rect 313844 317529 313872 319670
rect 313830 317520 313886 317529
rect 313830 317455 313886 317464
rect 313740 316260 313792 316266
rect 313740 316202 313792 316208
rect 313648 315308 313700 315314
rect 313648 315250 313700 315256
rect 313740 311636 313792 311642
rect 313740 311578 313792 311584
rect 313752 311506 313780 311578
rect 313740 311500 313792 311506
rect 313740 311442 313792 311448
rect 313556 310276 313608 310282
rect 313556 310218 313608 310224
rect 313462 307864 313518 307873
rect 313462 307799 313518 307808
rect 313568 306950 313596 310218
rect 313936 310078 313964 319756
rect 314014 319560 314070 319569
rect 314014 319495 314070 319504
rect 314028 317558 314056 319495
rect 314120 317626 314148 319756
rect 314304 319756 314378 319784
rect 314442 319784 314470 320076
rect 314534 319938 314562 320076
rect 314522 319932 314574 319938
rect 314522 319874 314574 319880
rect 314626 319870 314654 320076
rect 314614 319864 314666 319870
rect 314614 319806 314666 319812
rect 314442 319756 314516 319784
rect 314198 319424 314254 319433
rect 314198 319359 314254 319368
rect 314108 317620 314160 317626
rect 314108 317562 314160 317568
rect 314016 317552 314068 317558
rect 314016 317494 314068 317500
rect 314108 317484 314160 317490
rect 314108 317426 314160 317432
rect 313924 310072 313976 310078
rect 313924 310014 313976 310020
rect 313556 306944 313608 306950
rect 313556 306886 313608 306892
rect 313188 304088 313240 304094
rect 313188 304030 313240 304036
rect 313096 257372 313148 257378
rect 313096 257314 313148 257320
rect 312912 248532 312964 248538
rect 312912 248474 312964 248480
rect 312924 248414 312952 248474
rect 312832 248386 312952 248414
rect 312728 244996 312780 245002
rect 312728 244938 312780 244944
rect 312634 234152 312690 234161
rect 312634 234087 312690 234096
rect 312542 225992 312598 226001
rect 312542 225927 312598 225936
rect 311346 224904 311402 224913
rect 311346 224839 311402 224848
rect 312832 224738 312860 248386
rect 312912 244452 312964 244458
rect 312912 244394 312964 244400
rect 312820 224732 312872 224738
rect 312820 224674 312872 224680
rect 311256 223168 311308 223174
rect 311256 223110 311308 223116
rect 311164 223100 311216 223106
rect 311164 223042 311216 223048
rect 312924 222018 312952 244394
rect 312912 222012 312964 222018
rect 312912 221954 312964 221960
rect 309784 220108 309836 220114
rect 309784 220050 309836 220056
rect 308404 217320 308456 217326
rect 308404 217262 308456 217268
rect 307852 116680 307904 116686
rect 307852 116622 307904 116628
rect 307864 3602 307892 116622
rect 308416 3738 308444 217262
rect 308404 3732 308456 3738
rect 308404 3674 308456 3680
rect 307852 3596 307904 3602
rect 307852 3538 307904 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307772 3454 307984 3482
rect 307208 3188 307260 3194
rect 307208 3130 307260 3136
rect 307024 3052 307076 3058
rect 307024 2994 307076 3000
rect 307956 480 307984 3454
rect 309060 480 309088 3538
rect 309796 3330 309824 220050
rect 309876 142996 309928 143002
rect 309876 142938 309928 142944
rect 309888 3398 309916 142938
rect 311162 105496 311218 105505
rect 311162 105431 311218 105440
rect 311176 3534 311204 105431
rect 313200 4010 313228 304030
rect 313936 243710 313964 310014
rect 314014 308408 314070 308417
rect 314014 308343 314070 308352
rect 314028 307873 314056 308343
rect 314014 307864 314070 307873
rect 314014 307799 314070 307808
rect 314028 244934 314056 307799
rect 314120 305454 314148 317426
rect 314108 305448 314160 305454
rect 314108 305390 314160 305396
rect 314212 296714 314240 319359
rect 314304 316198 314332 319756
rect 314384 319660 314436 319666
rect 314384 319602 314436 319608
rect 314292 316192 314344 316198
rect 314292 316134 314344 316140
rect 314292 316056 314344 316062
rect 314292 315998 314344 316004
rect 314304 299198 314332 315998
rect 314396 315722 314424 319602
rect 314488 317529 314516 319756
rect 314718 319716 314746 320076
rect 314902 319954 314930 320076
rect 314672 319688 314746 319716
rect 314856 319926 314930 319954
rect 314672 318345 314700 319688
rect 314658 318336 314714 318345
rect 314658 318271 314714 318280
rect 314568 317620 314620 317626
rect 314568 317562 314620 317568
rect 314474 317520 314530 317529
rect 314474 317455 314530 317464
rect 314384 315716 314436 315722
rect 314384 315658 314436 315664
rect 314292 299192 314344 299198
rect 314292 299134 314344 299140
rect 314120 296686 314240 296714
rect 314120 292534 314148 296686
rect 314108 292528 314160 292534
rect 314108 292470 314160 292476
rect 314396 263702 314424 315658
rect 314580 315110 314608 317562
rect 314856 317121 314884 319926
rect 314994 319852 315022 320175
rect 315532 320104 315588 320113
rect 314948 319824 315022 319852
rect 314948 318073 314976 319824
rect 315086 319784 315114 320076
rect 315040 319756 315114 319784
rect 315178 319784 315206 320076
rect 315270 319938 315298 320076
rect 315258 319932 315310 319938
rect 315258 319874 315310 319880
rect 315362 319784 315390 320076
rect 315454 319852 315482 320076
rect 316636 320104 316692 320113
rect 315532 320039 315588 320048
rect 315454 319824 315528 319852
rect 315178 319756 315252 319784
rect 315040 318306 315068 319756
rect 315028 318300 315080 318306
rect 315028 318242 315080 318248
rect 314934 318064 314990 318073
rect 314934 317999 314990 318008
rect 314842 317112 314898 317121
rect 314842 317047 314898 317056
rect 315028 316192 315080 316198
rect 315028 316134 315080 316140
rect 314844 316056 314896 316062
rect 314844 315998 314896 316004
rect 314752 315920 314804 315926
rect 314752 315862 314804 315868
rect 314568 315104 314620 315110
rect 314568 315046 314620 315052
rect 314476 307148 314528 307154
rect 314476 307090 314528 307096
rect 314488 307057 314516 307090
rect 314474 307048 314530 307057
rect 314474 306983 314530 306992
rect 314476 306944 314528 306950
rect 314476 306886 314528 306892
rect 314108 263696 314160 263702
rect 314108 263638 314160 263644
rect 314384 263696 314436 263702
rect 314384 263638 314436 263644
rect 314016 244928 314068 244934
rect 314016 244870 314068 244876
rect 313924 243704 313976 243710
rect 313924 243646 313976 243652
rect 313924 242548 313976 242554
rect 313924 242490 313976 242496
rect 313936 218754 313964 242490
rect 314120 221882 314148 263638
rect 314200 249756 314252 249762
rect 314200 249698 314252 249704
rect 314212 248470 314240 249698
rect 314200 248464 314252 248470
rect 314488 248414 314516 306886
rect 314580 249762 314608 315046
rect 314764 305833 314792 315862
rect 314856 307057 314884 315998
rect 314936 315988 314988 315994
rect 314936 315930 314988 315936
rect 314948 307086 314976 315930
rect 315040 310554 315068 316134
rect 315224 312866 315252 319756
rect 315316 319756 315390 319784
rect 315316 316985 315344 319756
rect 315302 316976 315358 316985
rect 315302 316911 315358 316920
rect 315500 316198 315528 319824
rect 315638 319784 315666 320076
rect 315592 319756 315666 319784
rect 315730 319784 315758 320076
rect 315914 319954 315942 320076
rect 315868 319926 315942 319954
rect 315730 319756 315804 319784
rect 315488 316192 315540 316198
rect 315488 316134 315540 316140
rect 315592 315926 315620 319756
rect 315672 319660 315724 319666
rect 315672 319602 315724 319608
rect 315580 315920 315632 315926
rect 315580 315862 315632 315868
rect 315212 312860 315264 312866
rect 315212 312802 315264 312808
rect 315224 311894 315252 312802
rect 315224 311866 315436 311894
rect 315028 310548 315080 310554
rect 315028 310490 315080 310496
rect 314936 307080 314988 307086
rect 314842 307048 314898 307057
rect 314936 307022 314988 307028
rect 314842 306983 314898 306992
rect 314750 305824 314806 305833
rect 314750 305759 314806 305768
rect 315302 296848 315358 296857
rect 315302 296783 315358 296792
rect 314568 249756 314620 249762
rect 314568 249698 314620 249704
rect 314200 248406 314252 248412
rect 314108 221876 314160 221882
rect 314108 221818 314160 221824
rect 314212 221814 314240 248406
rect 314304 248386 314516 248414
rect 314304 247178 314332 248386
rect 314292 247172 314344 247178
rect 314292 247114 314344 247120
rect 314304 221950 314332 247114
rect 314292 221944 314344 221950
rect 314292 221886 314344 221892
rect 314200 221808 314252 221814
rect 314200 221750 314252 221756
rect 315316 219366 315344 296783
rect 315408 242554 315436 311866
rect 315580 307080 315632 307086
rect 315486 307048 315542 307057
rect 315580 307022 315632 307028
rect 315486 306983 315542 306992
rect 315500 243642 315528 306983
rect 315592 257417 315620 307022
rect 315684 304337 315712 319602
rect 315776 315790 315804 319756
rect 315868 316062 315896 319926
rect 316006 319784 316034 320076
rect 316098 319938 316126 320076
rect 316086 319932 316138 319938
rect 316086 319874 316138 319880
rect 316190 319818 316218 320076
rect 315960 319756 316034 319784
rect 316144 319790 316218 319818
rect 315856 316056 315908 316062
rect 315856 315998 315908 316004
rect 315960 315994 315988 319756
rect 316144 318782 316172 319790
rect 316282 319716 316310 320076
rect 316374 319784 316402 320076
rect 316466 319852 316494 320076
rect 316558 319954 316586 320076
rect 318292 320104 318348 320113
rect 316636 320039 316692 320048
rect 316742 319954 316770 320076
rect 316558 319926 316632 319954
rect 316466 319824 316540 319852
rect 316374 319756 316448 319784
rect 316282 319688 316356 319716
rect 316132 318776 316184 318782
rect 316132 318718 316184 318724
rect 316132 316260 316184 316266
rect 316132 316202 316184 316208
rect 315948 315988 316000 315994
rect 315948 315930 316000 315936
rect 315764 315784 315816 315790
rect 315764 315726 315816 315732
rect 315776 311894 315804 315726
rect 315776 311866 315896 311894
rect 315670 304328 315726 304337
rect 315670 304263 315726 304272
rect 315578 257408 315634 257417
rect 315578 257343 315634 257352
rect 315868 255338 315896 311866
rect 315948 311160 316000 311166
rect 315948 311102 316000 311108
rect 315960 310554 315988 311102
rect 315948 310548 316000 310554
rect 315948 310490 316000 310496
rect 315580 255332 315632 255338
rect 315580 255274 315632 255280
rect 315856 255332 315908 255338
rect 315856 255274 315908 255280
rect 315488 243636 315540 243642
rect 315488 243578 315540 243584
rect 315396 242548 315448 242554
rect 315396 242490 315448 242496
rect 315592 222057 315620 255274
rect 315960 251326 315988 310490
rect 316144 299402 316172 316202
rect 316328 316146 316356 319688
rect 316420 316266 316448 319756
rect 316512 318170 316540 319824
rect 316500 318164 316552 318170
rect 316500 318106 316552 318112
rect 316408 316260 316460 316266
rect 316408 316202 316460 316208
rect 316328 316118 316448 316146
rect 316224 316056 316276 316062
rect 316224 315998 316276 316004
rect 316236 309670 316264 315998
rect 316316 315988 316368 315994
rect 316316 315930 316368 315936
rect 316224 309664 316276 309670
rect 316224 309606 316276 309612
rect 316236 309194 316264 309606
rect 316328 309262 316356 315930
rect 316420 315586 316448 316118
rect 316408 315580 316460 315586
rect 316408 315522 316460 315528
rect 316604 311894 316632 319926
rect 316696 319926 316770 319954
rect 316696 316849 316724 319926
rect 316834 319784 316862 320076
rect 317018 319954 317046 320076
rect 316788 319756 316862 319784
rect 316972 319926 317046 319954
rect 316682 316840 316738 316849
rect 316682 316775 316738 316784
rect 316696 316402 316724 316775
rect 316684 316396 316736 316402
rect 316684 316338 316736 316344
rect 316788 315994 316816 319756
rect 316868 319660 316920 319666
rect 316868 319602 316920 319608
rect 316776 315988 316828 315994
rect 316776 315930 316828 315936
rect 316420 311866 316632 311894
rect 316420 311409 316448 311866
rect 316406 311400 316462 311409
rect 316406 311335 316462 311344
rect 316420 310593 316448 311335
rect 316406 310584 316462 310593
rect 316406 310519 316462 310528
rect 316316 309256 316368 309262
rect 316316 309198 316368 309204
rect 316224 309188 316276 309194
rect 316224 309130 316276 309136
rect 316684 309188 316736 309194
rect 316684 309130 316736 309136
rect 316132 299396 316184 299402
rect 316132 299338 316184 299344
rect 315672 251320 315724 251326
rect 315672 251262 315724 251268
rect 315948 251320 316000 251326
rect 315948 251262 316000 251268
rect 315684 225826 315712 251262
rect 316696 249150 316724 309130
rect 316776 299396 316828 299402
rect 316776 299338 316828 299344
rect 316788 299130 316816 299338
rect 316776 299124 316828 299130
rect 316776 299066 316828 299072
rect 316788 267073 316816 299066
rect 316880 297537 316908 319602
rect 316972 316062 317000 319926
rect 317110 319852 317138 320076
rect 317064 319824 317138 319852
rect 316960 316056 317012 316062
rect 317064 316033 317092 319824
rect 317202 319784 317230 320076
rect 317156 319756 317230 319784
rect 317294 319784 317322 320076
rect 317386 319938 317414 320076
rect 317374 319932 317426 319938
rect 317374 319874 317426 319880
rect 317478 319784 317506 320076
rect 317570 319938 317598 320076
rect 317558 319932 317610 319938
rect 317558 319874 317610 319880
rect 317662 319784 317690 320076
rect 317294 319756 317368 319784
rect 317156 319569 317184 319756
rect 317236 319660 317288 319666
rect 317236 319602 317288 319608
rect 317142 319560 317198 319569
rect 317142 319495 317198 319504
rect 317156 318073 317184 319495
rect 317142 318064 317198 318073
rect 317142 317999 317198 318008
rect 316960 315998 317012 316004
rect 317050 316024 317106 316033
rect 317050 315959 317106 315968
rect 316960 309732 317012 309738
rect 316960 309674 317012 309680
rect 316972 309262 317000 309674
rect 316960 309256 317012 309262
rect 316960 309198 317012 309204
rect 316866 297528 316922 297537
rect 316866 297463 316922 297472
rect 316880 296857 316908 297463
rect 316866 296848 316922 296857
rect 316866 296783 316922 296792
rect 316774 267064 316830 267073
rect 316774 266999 316830 267008
rect 316972 258126 317000 309198
rect 317064 264654 317092 315959
rect 317248 315042 317276 319602
rect 317340 317801 317368 319756
rect 317432 319756 317506 319784
rect 317616 319756 317690 319784
rect 317754 319784 317782 320076
rect 317938 319818 317966 320076
rect 317892 319790 317966 319818
rect 317754 319756 317828 319784
rect 317326 317792 317382 317801
rect 317326 317727 317382 317736
rect 317328 317552 317380 317558
rect 317328 317494 317380 317500
rect 317340 317082 317368 317494
rect 317328 317076 317380 317082
rect 317328 317018 317380 317024
rect 317328 315580 317380 315586
rect 317328 315522 317380 315528
rect 317236 315036 317288 315042
rect 317236 314978 317288 314984
rect 317142 312760 317198 312769
rect 317142 312695 317144 312704
rect 317196 312695 317198 312704
rect 317144 312666 317196 312672
rect 317142 310584 317198 310593
rect 317142 310519 317198 310528
rect 317052 264648 317104 264654
rect 317052 264590 317104 264596
rect 316960 258120 317012 258126
rect 316880 258068 316960 258074
rect 316880 258062 317012 258068
rect 316880 258046 317000 258062
rect 316776 253088 316828 253094
rect 316776 253030 316828 253036
rect 316684 249144 316736 249150
rect 316684 249086 316736 249092
rect 316684 245676 316736 245682
rect 316684 245618 316736 245624
rect 315672 225820 315724 225826
rect 315672 225762 315724 225768
rect 316696 223378 316724 245618
rect 316788 224641 316816 253030
rect 316880 231674 316908 258046
rect 317156 250510 317184 310519
rect 317248 253094 317276 314978
rect 317340 314838 317368 315522
rect 317328 314832 317380 314838
rect 317328 314774 317380 314780
rect 317236 253088 317288 253094
rect 317236 253030 317288 253036
rect 317248 252686 317276 253030
rect 317236 252680 317288 252686
rect 317236 252622 317288 252628
rect 317144 250504 317196 250510
rect 317144 250446 317196 250452
rect 317340 245682 317368 314774
rect 317432 299402 317460 319756
rect 317512 318504 317564 318510
rect 317512 318446 317564 318452
rect 317524 317014 317552 318446
rect 317512 317008 317564 317014
rect 317512 316950 317564 316956
rect 317512 316600 317564 316606
rect 317512 316542 317564 316548
rect 317524 315246 317552 316542
rect 317512 315240 317564 315246
rect 317512 315182 317564 315188
rect 317524 314906 317552 315182
rect 317512 314900 317564 314906
rect 317512 314842 317564 314848
rect 317616 311894 317644 319756
rect 317696 319660 317748 319666
rect 317696 319602 317748 319608
rect 317708 316606 317736 319602
rect 317800 317801 317828 319756
rect 317786 317792 317842 317801
rect 317786 317727 317842 317736
rect 317696 316600 317748 316606
rect 317696 316542 317748 316548
rect 317696 315988 317748 315994
rect 317696 315930 317748 315936
rect 317524 311866 317644 311894
rect 317524 310418 317552 311866
rect 317708 311681 317736 315930
rect 317892 314566 317920 319790
rect 318030 319784 318058 320076
rect 318122 319852 318150 320076
rect 318214 319954 318242 320076
rect 318844 320104 318900 320113
rect 318292 320039 318348 320048
rect 318398 319954 318426 320076
rect 318214 319926 318334 319954
rect 318398 319926 318472 319954
rect 318306 319852 318334 319926
rect 318122 319824 318196 319852
rect 318306 319824 318380 319852
rect 318030 319756 318104 319784
rect 318076 317529 318104 319756
rect 318168 317937 318196 319824
rect 318154 317928 318210 317937
rect 318154 317863 318210 317872
rect 318062 317520 318118 317529
rect 318062 317455 318118 317464
rect 318064 315920 318116 315926
rect 318064 315862 318116 315868
rect 317880 314560 317932 314566
rect 317880 314502 317932 314508
rect 317880 313812 317932 313818
rect 317880 313754 317932 313760
rect 317694 311672 317750 311681
rect 317694 311607 317750 311616
rect 317512 310412 317564 310418
rect 317512 310354 317564 310360
rect 317524 309194 317552 310354
rect 317512 309188 317564 309194
rect 317512 309130 317564 309136
rect 317512 303612 317564 303618
rect 317512 303554 317564 303560
rect 317524 303521 317552 303554
rect 317510 303512 317566 303521
rect 317510 303447 317566 303456
rect 317524 302841 317552 303447
rect 317510 302832 317566 302841
rect 317510 302767 317566 302776
rect 317892 302234 317920 313754
rect 318076 311545 318104 315862
rect 318352 315466 318380 319824
rect 318444 315994 318472 319926
rect 318582 319852 318610 320076
rect 318674 319938 318702 320076
rect 318662 319932 318714 319938
rect 318662 319874 318714 319880
rect 318536 319824 318610 319852
rect 318432 315988 318484 315994
rect 318432 315930 318484 315936
rect 318536 315926 318564 319824
rect 318766 319818 318794 320076
rect 319488 320104 319544 320113
rect 318844 320039 318900 320048
rect 318858 319870 318886 320039
rect 318674 319790 318794 319818
rect 318846 319864 318898 319870
rect 318846 319806 318898 319812
rect 318674 319784 318702 319790
rect 318628 319756 318702 319784
rect 318524 315920 318576 315926
rect 318524 315862 318576 315868
rect 318628 315602 318656 319756
rect 318950 319716 318978 320076
rect 319042 319784 319070 320076
rect 319226 319938 319254 320076
rect 319214 319932 319266 319938
rect 319214 319874 319266 319880
rect 319318 319818 319346 320076
rect 319410 319938 319438 320076
rect 320040 320104 320096 320113
rect 319488 320039 319544 320048
rect 319398 319932 319450 319938
rect 319398 319874 319450 319880
rect 319318 319790 319484 319818
rect 319042 319756 319208 319784
rect 318950 319688 319024 319716
rect 318708 319660 318760 319666
rect 318708 319602 318760 319608
rect 318800 319660 318852 319666
rect 318800 319602 318852 319608
rect 318720 318073 318748 319602
rect 318706 318064 318762 318073
rect 318706 317999 318762 318008
rect 318812 317937 318840 319602
rect 318996 319433 319024 319688
rect 318982 319424 319038 319433
rect 318982 319359 319038 319368
rect 318890 318336 318946 318345
rect 318890 318271 318946 318280
rect 318798 317928 318854 317937
rect 318798 317863 318854 317872
rect 318904 317801 318932 318271
rect 318890 317792 318946 317801
rect 318890 317727 318946 317736
rect 318628 315574 318748 315602
rect 318352 315438 318656 315466
rect 318432 314560 318484 314566
rect 318432 314502 318484 314508
rect 318444 314294 318472 314502
rect 318628 314498 318656 315438
rect 318616 314492 318668 314498
rect 318616 314434 318668 314440
rect 318432 314288 318484 314294
rect 318432 314230 318484 314236
rect 318062 311536 318118 311545
rect 318062 311471 318118 311480
rect 318076 311001 318104 311471
rect 318062 310992 318118 311001
rect 318062 310927 318118 310936
rect 317892 302206 318196 302234
rect 317420 299396 317472 299402
rect 317420 299338 317472 299344
rect 318064 299396 318116 299402
rect 318064 299338 318116 299344
rect 318076 299198 318104 299338
rect 318064 299192 318116 299198
rect 318064 299134 318116 299140
rect 317420 264648 317472 264654
rect 317420 264590 317472 264596
rect 317432 263634 317460 264590
rect 317420 263628 317472 263634
rect 317420 263570 317472 263576
rect 317328 245676 317380 245682
rect 317328 245618 317380 245624
rect 316868 231668 316920 231674
rect 316868 231610 316920 231616
rect 316774 224632 316830 224641
rect 316774 224567 316830 224576
rect 317432 223417 317460 263570
rect 317418 223408 317474 223417
rect 316684 223372 316736 223378
rect 317418 223343 317474 223352
rect 316684 223314 316736 223320
rect 315578 222048 315634 222057
rect 315578 221983 315634 221992
rect 318076 220182 318104 299134
rect 318168 260137 318196 302206
rect 318248 262744 318300 262750
rect 318248 262686 318300 262692
rect 318260 262274 318288 262686
rect 318248 262268 318300 262274
rect 318248 262210 318300 262216
rect 318154 260128 318210 260137
rect 318154 260063 318210 260072
rect 318156 247104 318208 247110
rect 318156 247046 318208 247052
rect 318168 223242 318196 247046
rect 318260 223446 318288 262210
rect 318444 248414 318472 314230
rect 318524 309188 318576 309194
rect 318524 309130 318576 309136
rect 318536 262750 318564 309130
rect 318524 262744 318576 262750
rect 318524 262686 318576 262692
rect 318352 248386 318472 248414
rect 318352 244390 318380 248386
rect 318628 247110 318656 314434
rect 318720 313818 318748 315574
rect 319180 314673 319208 319756
rect 319260 319660 319312 319666
rect 319260 319602 319312 319608
rect 319352 319660 319404 319666
rect 319352 319602 319404 319608
rect 319272 315353 319300 319602
rect 319364 318617 319392 319602
rect 319350 318608 319406 318617
rect 319350 318543 319406 318552
rect 319456 316606 319484 319790
rect 319594 319784 319622 320076
rect 319778 319784 319806 320076
rect 319962 319870 319990 320076
rect 320500 320104 320556 320113
rect 320040 320039 320096 320048
rect 319950 319864 320002 319870
rect 319950 319806 320002 319812
rect 319548 319756 319622 319784
rect 319732 319756 319806 319784
rect 319444 316600 319496 316606
rect 319444 316542 319496 316548
rect 319258 315344 319314 315353
rect 319258 315279 319314 315288
rect 319166 314664 319222 314673
rect 319166 314599 319222 314608
rect 319548 314129 319576 319756
rect 319732 319648 319760 319756
rect 320146 319716 320174 320076
rect 320238 319784 320266 320076
rect 320330 319938 320358 320076
rect 320318 319932 320370 319938
rect 320318 319874 320370 319880
rect 320422 319852 320450 320076
rect 321328 320104 321384 320113
rect 320500 320039 320556 320048
rect 320548 319932 320600 319938
rect 320698 319920 320726 320076
rect 320600 319892 320726 319920
rect 320548 319874 320600 319880
rect 320790 319852 320818 320076
rect 320422 319824 320496 319852
rect 320238 319756 320312 319784
rect 320100 319688 320174 319716
rect 319904 319660 319956 319666
rect 319732 319620 319806 319648
rect 319778 319546 319806 319620
rect 319904 319602 319956 319608
rect 319778 319518 319852 319546
rect 319626 319016 319682 319025
rect 319626 318951 319682 318960
rect 319534 314120 319590 314129
rect 319534 314055 319590 314064
rect 318708 313812 318760 313818
rect 318708 313754 318760 313760
rect 319444 313744 319496 313750
rect 319444 313686 319496 313692
rect 318706 300792 318762 300801
rect 318706 300727 318762 300736
rect 318720 300422 318748 300727
rect 318708 300416 318760 300422
rect 318708 300358 318760 300364
rect 318708 299396 318760 299402
rect 318708 299338 318760 299344
rect 318720 298897 318748 299338
rect 318706 298888 318762 298897
rect 318706 298823 318762 298832
rect 318720 297265 318748 298823
rect 318706 297256 318762 297265
rect 318706 297191 318762 297200
rect 318616 247104 318668 247110
rect 318616 247046 318668 247052
rect 318340 244384 318392 244390
rect 318340 244326 318392 244332
rect 318352 223514 318380 244326
rect 318340 223508 318392 223514
rect 318340 223450 318392 223456
rect 318248 223440 318300 223446
rect 318248 223382 318300 223388
rect 319456 223310 319484 313686
rect 319548 242457 319576 314055
rect 319640 308242 319668 318951
rect 319718 318880 319774 318889
rect 319718 318815 319774 318824
rect 319732 315654 319760 318815
rect 319824 315858 319852 319518
rect 319812 315852 319864 315858
rect 319812 315794 319864 315800
rect 319720 315648 319772 315654
rect 319720 315590 319772 315596
rect 319916 314786 319944 319602
rect 319994 319016 320050 319025
rect 319994 318951 320050 318960
rect 319824 314758 319944 314786
rect 319824 313750 319852 314758
rect 319902 314664 319958 314673
rect 319902 314599 319958 314608
rect 319916 313993 319944 314599
rect 319902 313984 319958 313993
rect 319902 313919 319958 313928
rect 319812 313744 319864 313750
rect 319812 313686 319864 313692
rect 319628 308236 319680 308242
rect 319628 308178 319680 308184
rect 319534 242448 319590 242457
rect 319534 242383 319590 242392
rect 319640 238202 319668 308178
rect 319916 258074 319944 313919
rect 320008 309602 320036 318951
rect 320100 318481 320128 319688
rect 320180 318844 320232 318850
rect 320180 318786 320232 318792
rect 320086 318472 320142 318481
rect 320086 318407 320142 318416
rect 320088 316600 320140 316606
rect 320088 316542 320140 316548
rect 319996 309596 320048 309602
rect 319996 309538 320048 309544
rect 319732 258046 319944 258074
rect 319732 256766 319760 258046
rect 319720 256760 319772 256766
rect 319720 256702 319772 256708
rect 319628 238196 319680 238202
rect 319628 238138 319680 238144
rect 319732 223582 319760 256702
rect 320008 242434 320036 309538
rect 320100 243030 320128 316542
rect 320192 303346 320220 318786
rect 320284 318073 320312 319756
rect 320364 319728 320416 319734
rect 320364 319670 320416 319676
rect 320376 318753 320404 319670
rect 320362 318744 320418 318753
rect 320362 318679 320418 318688
rect 320270 318064 320326 318073
rect 320270 317999 320326 318008
rect 320468 316198 320496 319824
rect 320744 319824 320818 319852
rect 320548 319796 320600 319802
rect 320548 319738 320600 319744
rect 320560 318850 320588 319738
rect 320638 319560 320694 319569
rect 320638 319495 320694 319504
rect 320548 318844 320600 318850
rect 320548 318786 320600 318792
rect 320548 318504 320600 318510
rect 320548 318446 320600 318452
rect 320456 316192 320508 316198
rect 320456 316134 320508 316140
rect 320456 315988 320508 315994
rect 320456 315930 320508 315936
rect 320468 304745 320496 315930
rect 320560 310049 320588 318446
rect 320652 317490 320680 319495
rect 320744 318510 320772 319824
rect 320882 319784 320910 320076
rect 320836 319756 320910 319784
rect 320732 318504 320784 318510
rect 320732 318446 320784 318452
rect 320730 318336 320786 318345
rect 320730 318271 320786 318280
rect 320640 317484 320692 317490
rect 320640 317426 320692 317432
rect 320744 315518 320772 318271
rect 320732 315512 320784 315518
rect 320732 315454 320784 315460
rect 320836 315466 320864 319756
rect 320974 319682 321002 320076
rect 321066 319784 321094 320076
rect 321158 319938 321186 320076
rect 321146 319932 321198 319938
rect 321146 319874 321198 319880
rect 321250 319784 321278 320076
rect 322800 320104 322856 320113
rect 321328 320039 321384 320048
rect 321434 319954 321462 320076
rect 321066 319756 321140 319784
rect 320928 319654 321002 319682
rect 320928 317529 320956 319654
rect 321112 319546 321140 319756
rect 321020 319518 321140 319546
rect 321204 319756 321278 319784
rect 321388 319926 321462 319954
rect 321020 317937 321048 319518
rect 321098 318744 321154 318753
rect 321098 318679 321154 318688
rect 321006 317928 321062 317937
rect 321006 317863 321062 317872
rect 321112 317529 321140 318679
rect 320914 317520 320970 317529
rect 320914 317455 320970 317464
rect 321098 317520 321154 317529
rect 321098 317455 321154 317464
rect 321100 316940 321152 316946
rect 321100 316882 321152 316888
rect 320836 315438 321048 315466
rect 321020 315382 321048 315438
rect 321008 315376 321060 315382
rect 321008 315318 321060 315324
rect 321112 314022 321140 316882
rect 321100 314016 321152 314022
rect 321100 313958 321152 313964
rect 320822 313304 320878 313313
rect 320822 313239 320878 313248
rect 320546 310040 320602 310049
rect 320546 309975 320602 309984
rect 320454 304736 320510 304745
rect 320454 304671 320510 304680
rect 320732 303544 320784 303550
rect 320732 303486 320784 303492
rect 320180 303340 320232 303346
rect 320180 303282 320232 303288
rect 320744 301374 320772 303486
rect 320732 301368 320784 301374
rect 320732 301310 320784 301316
rect 320088 243024 320140 243030
rect 320088 242966 320140 242972
rect 320100 242593 320128 242966
rect 320086 242584 320142 242593
rect 320086 242519 320142 242528
rect 320008 242406 320128 242434
rect 320100 241602 320128 242406
rect 320088 241596 320140 241602
rect 320088 241538 320140 241544
rect 320100 241058 320128 241538
rect 320088 241052 320140 241058
rect 320088 240994 320140 241000
rect 319720 223576 319772 223582
rect 319720 223518 319772 223524
rect 319444 223304 319496 223310
rect 319444 223246 319496 223252
rect 318156 223236 318208 223242
rect 318156 223178 318208 223184
rect 320836 221474 320864 313239
rect 321008 312452 321060 312458
rect 321008 312394 321060 312400
rect 320914 305008 320970 305017
rect 320914 304943 320970 304952
rect 320928 303550 320956 304943
rect 320916 303544 320968 303550
rect 320916 303486 320968 303492
rect 320916 303408 320968 303414
rect 320916 303350 320968 303356
rect 320928 242185 320956 303350
rect 321020 253201 321048 312394
rect 321098 310040 321154 310049
rect 321098 309975 321154 309984
rect 321112 303414 321140 309975
rect 321204 303414 321232 319756
rect 321284 319660 321336 319666
rect 321284 319602 321336 319608
rect 321296 316946 321324 319602
rect 321284 316940 321336 316946
rect 321284 316882 321336 316888
rect 321284 316328 321336 316334
rect 321284 316270 321336 316276
rect 321296 312458 321324 316270
rect 321388 315994 321416 319926
rect 321526 319784 321554 320076
rect 321480 319756 321554 319784
rect 321480 316334 321508 319756
rect 321618 319682 321646 320076
rect 321802 319954 321830 320076
rect 321572 319654 321646 319682
rect 321756 319926 321830 319954
rect 321468 316328 321520 316334
rect 321468 316270 321520 316276
rect 321468 316192 321520 316198
rect 321468 316134 321520 316140
rect 321376 315988 321428 315994
rect 321376 315930 321428 315936
rect 321284 312452 321336 312458
rect 321284 312394 321336 312400
rect 321282 304736 321338 304745
rect 321282 304671 321338 304680
rect 321100 303408 321152 303414
rect 321100 303350 321152 303356
rect 321192 303408 321244 303414
rect 321192 303350 321244 303356
rect 321100 303272 321152 303278
rect 321100 303214 321152 303220
rect 321112 253230 321140 303214
rect 321204 286346 321232 303350
rect 321296 303278 321324 304671
rect 321480 303346 321508 316134
rect 321572 315217 321600 319654
rect 321756 316713 321784 319926
rect 321894 319852 321922 320076
rect 321848 319824 321922 319852
rect 321742 316704 321798 316713
rect 321742 316639 321798 316648
rect 321848 316198 321876 319824
rect 321986 319784 322014 320076
rect 321940 319756 322014 319784
rect 321940 317558 321968 319756
rect 322078 319682 322106 320076
rect 322170 319870 322198 320076
rect 322158 319864 322210 319870
rect 322158 319806 322210 319812
rect 322262 319818 322290 320076
rect 322354 319920 322382 320076
rect 322538 319920 322566 320076
rect 322354 319892 322428 319920
rect 322262 319790 322336 319818
rect 322204 319728 322256 319734
rect 322078 319654 322152 319682
rect 322204 319670 322256 319676
rect 322018 318472 322074 318481
rect 322018 318407 322074 318416
rect 322032 317665 322060 318407
rect 322018 317656 322074 317665
rect 322018 317591 322074 317600
rect 321928 317552 321980 317558
rect 321928 317494 321980 317500
rect 321836 316192 321888 316198
rect 321836 316134 321888 316140
rect 322124 316010 322152 319654
rect 322216 317665 322244 319670
rect 322202 317656 322258 317665
rect 322202 317591 322258 317600
rect 321664 315982 322152 316010
rect 321558 315208 321614 315217
rect 321558 315143 321614 315152
rect 321572 313313 321600 315143
rect 321558 313304 321614 313313
rect 321558 313239 321614 313248
rect 321560 312180 321612 312186
rect 321560 312122 321612 312128
rect 321572 311506 321600 312122
rect 321560 311500 321612 311506
rect 321560 311442 321612 311448
rect 321664 305182 321692 315982
rect 322308 314922 322336 319790
rect 322400 316169 322428 319892
rect 322492 319892 322566 319920
rect 322492 317354 322520 319892
rect 322630 319852 322658 320076
rect 322584 319824 322658 319852
rect 322480 317348 322532 317354
rect 322480 317290 322532 317296
rect 322478 317248 322534 317257
rect 322478 317183 322534 317192
rect 322492 316713 322520 317183
rect 322478 316704 322534 316713
rect 322478 316639 322534 316648
rect 322584 316282 322612 319824
rect 322722 319784 322750 320076
rect 323352 320104 323408 320113
rect 322800 320039 322856 320048
rect 322906 319954 322934 320076
rect 322906 319926 322980 319954
rect 322676 319756 322750 319784
rect 322676 317529 322704 319756
rect 322848 319660 322900 319666
rect 322848 319602 322900 319608
rect 322860 318714 322888 319602
rect 322848 318708 322900 318714
rect 322848 318650 322900 318656
rect 322952 318594 322980 319926
rect 323090 319920 323118 320076
rect 323044 319892 323118 319920
rect 323044 319734 323072 319892
rect 323182 319818 323210 320076
rect 323274 319920 323302 320076
rect 324180 320104 324236 320113
rect 323352 320039 323408 320048
rect 323458 319954 323486 320076
rect 323458 319926 323532 319954
rect 323274 319892 323348 319920
rect 323136 319790 323210 319818
rect 323032 319728 323084 319734
rect 323032 319670 323084 319676
rect 322768 318566 322980 318594
rect 322662 317520 322718 317529
rect 322662 317455 322718 317464
rect 322664 317348 322716 317354
rect 322664 317290 322716 317296
rect 322492 316254 322612 316282
rect 322386 316160 322442 316169
rect 322386 316095 322442 316104
rect 322124 314894 322336 314922
rect 322124 313274 322152 314894
rect 322492 314786 322520 316254
rect 322572 316192 322624 316198
rect 322572 316134 322624 316140
rect 322216 314758 322520 314786
rect 322112 313268 322164 313274
rect 322112 313210 322164 313216
rect 322124 312390 322152 313210
rect 322112 312384 322164 312390
rect 322112 312326 322164 312332
rect 322216 311894 322244 314758
rect 322294 314664 322350 314673
rect 322294 314599 322350 314608
rect 321756 311866 322244 311894
rect 321756 310321 321784 311866
rect 321742 310312 321798 310321
rect 321742 310247 321798 310256
rect 322202 307592 322258 307601
rect 322202 307527 322258 307536
rect 321652 305176 321704 305182
rect 321652 305118 321704 305124
rect 321468 303340 321520 303346
rect 321468 303282 321520 303288
rect 321284 303272 321336 303278
rect 321284 303214 321336 303220
rect 321376 303272 321428 303278
rect 321376 303214 321428 303220
rect 321284 301368 321336 301374
rect 321284 301310 321336 301316
rect 321192 286340 321244 286346
rect 321192 286282 321244 286288
rect 321296 273290 321324 301310
rect 321284 273284 321336 273290
rect 321284 273226 321336 273232
rect 321100 253224 321152 253230
rect 321006 253192 321062 253201
rect 321100 253166 321152 253172
rect 321006 253127 321062 253136
rect 321388 251258 321416 303214
rect 321376 251252 321428 251258
rect 321376 251194 321428 251200
rect 320914 242176 320970 242185
rect 320914 242111 320970 242120
rect 321008 241528 321060 241534
rect 321008 241470 321060 241476
rect 321020 240990 321048 241470
rect 321008 240984 321060 240990
rect 321008 240926 321060 240932
rect 321388 238754 321416 251194
rect 321480 241534 321508 303282
rect 321652 273284 321704 273290
rect 321652 273226 321704 273232
rect 321560 244316 321612 244322
rect 321560 244258 321612 244264
rect 321572 243574 321600 244258
rect 321560 243568 321612 243574
rect 321560 243510 321612 243516
rect 321560 242956 321612 242962
rect 321560 242898 321612 242904
rect 321572 242282 321600 242898
rect 321560 242276 321612 242282
rect 321560 242218 321612 242224
rect 321468 241528 321520 241534
rect 321468 241470 321520 241476
rect 321020 238726 321416 238754
rect 321020 227730 321048 238726
rect 321560 236700 321612 236706
rect 321560 236642 321612 236648
rect 321008 227724 321060 227730
rect 321008 227666 321060 227672
rect 320824 221468 320876 221474
rect 320824 221410 320876 221416
rect 318064 220176 318116 220182
rect 318064 220118 318116 220124
rect 315304 219360 315356 219366
rect 315304 219302 315356 219308
rect 313924 218748 313976 218754
rect 313924 218690 313976 218696
rect 313188 4004 313240 4010
rect 313188 3946 313240 3952
rect 311440 3596 311492 3602
rect 311440 3538 311492 3544
rect 311164 3528 311216 3534
rect 311164 3470 311216 3476
rect 309876 3392 309928 3398
rect 309876 3334 309928 3340
rect 309784 3324 309836 3330
rect 309784 3266 309836 3272
rect 310244 3188 310296 3194
rect 310244 3130 310296 3136
rect 310256 480 310284 3130
rect 311452 480 311480 3538
rect 313936 3534 313964 218690
rect 316684 147008 316736 147014
rect 316684 146950 316736 146956
rect 314016 140140 314068 140146
rect 314016 140082 314068 140088
rect 314028 4078 314056 140082
rect 315302 113928 315358 113937
rect 315302 113863 315358 113872
rect 315316 4214 315344 113863
rect 315396 22772 315448 22778
rect 315396 22714 315448 22720
rect 315304 4208 315356 4214
rect 315304 4150 315356 4156
rect 315408 4146 315436 22714
rect 316696 4146 316724 146950
rect 320180 138780 320232 138786
rect 320180 138722 320232 138728
rect 318798 119504 318854 119513
rect 318798 119439 318854 119448
rect 318812 16574 318840 119439
rect 320192 16574 320220 138722
rect 321572 16574 321600 236642
rect 321664 227526 321692 273226
rect 322216 249121 322244 307527
rect 322308 260166 322336 314599
rect 322584 306374 322612 316134
rect 322676 314673 322704 317290
rect 322662 314664 322718 314673
rect 322662 314599 322718 314608
rect 322768 312390 322796 318566
rect 322846 317928 322902 317937
rect 322846 317863 322902 317872
rect 322860 312798 322888 317863
rect 323032 315988 323084 315994
rect 323032 315930 323084 315936
rect 322848 312792 322900 312798
rect 322848 312734 322900 312740
rect 322860 312594 322888 312734
rect 322848 312588 322900 312594
rect 322848 312530 322900 312536
rect 322756 312384 322808 312390
rect 322756 312326 322808 312332
rect 322768 311894 322796 312326
rect 322768 311866 322888 311894
rect 322662 310312 322718 310321
rect 322662 310247 322718 310256
rect 322400 306346 322612 306374
rect 322400 304609 322428 306346
rect 322386 304600 322442 304609
rect 322386 304535 322442 304544
rect 322296 260160 322348 260166
rect 322296 260102 322348 260108
rect 322400 258777 322428 304535
rect 322676 276078 322704 310247
rect 322756 305516 322808 305522
rect 322756 305458 322808 305464
rect 322768 305182 322796 305458
rect 322756 305176 322808 305182
rect 322756 305118 322808 305124
rect 322664 276072 322716 276078
rect 322664 276014 322716 276020
rect 322386 258768 322442 258777
rect 322386 258703 322442 258712
rect 322202 249112 322258 249121
rect 322202 249047 322258 249056
rect 322768 244322 322796 305118
rect 322756 244316 322808 244322
rect 322756 244258 322808 244264
rect 322860 242962 322888 311866
rect 323044 303249 323072 315930
rect 323136 313041 323164 319790
rect 323216 319728 323268 319734
rect 323216 319670 323268 319676
rect 323228 318646 323256 319670
rect 323216 318640 323268 318646
rect 323216 318582 323268 318588
rect 323122 313032 323178 313041
rect 323122 312967 323178 312976
rect 323320 311894 323348 319892
rect 323504 319784 323532 319926
rect 323642 319852 323670 320076
rect 323412 319756 323532 319784
rect 323596 319824 323670 319852
rect 323412 315994 323440 319756
rect 323490 319560 323546 319569
rect 323490 319495 323546 319504
rect 323504 317665 323532 319495
rect 323490 317656 323546 317665
rect 323490 317591 323546 317600
rect 323596 317370 323624 319824
rect 323734 319784 323762 320076
rect 323504 317342 323624 317370
rect 323688 319756 323762 319784
rect 323504 316130 323532 317342
rect 323584 317280 323636 317286
rect 323584 317222 323636 317228
rect 323492 316124 323544 316130
rect 323492 316066 323544 316072
rect 323596 316010 323624 317222
rect 323688 316305 323716 319756
rect 323826 319682 323854 320076
rect 323918 319818 323946 320076
rect 324010 319954 324038 320076
rect 324456 320104 324512 320113
rect 324180 320039 324236 320048
rect 324010 319938 324084 319954
rect 324010 319932 324096 319938
rect 324010 319926 324044 319932
rect 324286 319920 324314 320076
rect 324916 320104 324972 320113
rect 324456 320039 324512 320048
rect 324044 319874 324096 319880
rect 324240 319892 324314 319920
rect 323918 319790 324084 319818
rect 323780 319654 323854 319682
rect 323952 319728 324004 319734
rect 323952 319670 324004 319676
rect 323780 319569 323808 319654
rect 323766 319560 323822 319569
rect 323766 319495 323822 319504
rect 323860 318504 323912 318510
rect 323860 318446 323912 318452
rect 323674 316296 323730 316305
rect 323674 316231 323730 316240
rect 323766 316160 323822 316169
rect 323676 316124 323728 316130
rect 323766 316095 323822 316104
rect 323676 316066 323728 316072
rect 323400 315988 323452 315994
rect 323400 315930 323452 315936
rect 323504 315982 323624 316010
rect 323136 311866 323348 311894
rect 323136 309097 323164 311866
rect 323122 309088 323178 309097
rect 323122 309023 323178 309032
rect 323030 303240 323086 303249
rect 323030 303175 323086 303184
rect 323504 289134 323532 315982
rect 323582 313168 323638 313177
rect 323582 313103 323638 313112
rect 323596 312769 323624 313103
rect 323582 312760 323638 312769
rect 323582 312695 323638 312704
rect 323492 289128 323544 289134
rect 323492 289070 323544 289076
rect 322940 276072 322992 276078
rect 322940 276014 322992 276020
rect 322848 242956 322900 242962
rect 322848 242898 322900 242904
rect 322952 238134 322980 276014
rect 323032 249824 323084 249830
rect 323032 249766 323084 249772
rect 323044 249082 323072 249766
rect 323032 249076 323084 249082
rect 323032 249018 323084 249024
rect 323596 246265 323624 312695
rect 323688 309466 323716 316066
rect 323676 309460 323728 309466
rect 323676 309402 323728 309408
rect 323674 309088 323730 309097
rect 323674 309023 323730 309032
rect 323688 308689 323716 309023
rect 323674 308680 323730 308689
rect 323674 308615 323730 308624
rect 323688 247625 323716 308615
rect 323780 307698 323808 316095
rect 323872 313857 323900 318446
rect 323964 316282 323992 319670
rect 324056 318510 324084 319790
rect 324240 319410 324268 319892
rect 324562 319870 324590 320076
rect 324550 319864 324602 319870
rect 324746 319852 324774 320076
rect 324550 319806 324602 319812
rect 324700 319824 324774 319852
rect 324320 319796 324372 319802
rect 324320 319738 324372 319744
rect 324148 319382 324268 319410
rect 324044 318504 324096 318510
rect 324044 318446 324096 318452
rect 324042 318336 324098 318345
rect 324042 318271 324098 318280
rect 324056 316441 324084 318271
rect 324148 317286 324176 319382
rect 324228 318844 324280 318850
rect 324228 318786 324280 318792
rect 324240 318714 324268 318786
rect 324228 318708 324280 318714
rect 324228 318650 324280 318656
rect 324228 318232 324280 318238
rect 324228 318174 324280 318180
rect 324136 317280 324188 317286
rect 324136 317222 324188 317228
rect 324240 316946 324268 318174
rect 324228 316940 324280 316946
rect 324228 316882 324280 316888
rect 324136 316872 324188 316878
rect 324136 316814 324188 316820
rect 324042 316432 324098 316441
rect 324042 316367 324098 316376
rect 323964 316254 324084 316282
rect 324056 315058 324084 316254
rect 324148 315926 324176 316814
rect 324228 316804 324280 316810
rect 324228 316746 324280 316752
rect 324136 315920 324188 315926
rect 324136 315862 324188 315868
rect 324240 315489 324268 316746
rect 324226 315480 324282 315489
rect 324226 315415 324282 315424
rect 324056 315030 324268 315058
rect 323858 313848 323914 313857
rect 323858 313783 323914 313792
rect 324240 313177 324268 315030
rect 324226 313168 324282 313177
rect 324226 313103 324282 313112
rect 324134 313032 324190 313041
rect 324134 312967 324190 312976
rect 324148 312633 324176 312967
rect 324134 312624 324190 312633
rect 324134 312559 324190 312568
rect 323768 307692 323820 307698
rect 323768 307634 323820 307640
rect 323950 303512 324006 303521
rect 323950 303447 324006 303456
rect 323964 277438 323992 303447
rect 324042 303240 324098 303249
rect 324042 303175 324098 303184
rect 323952 277432 324004 277438
rect 323952 277374 324004 277380
rect 324056 258074 324084 303175
rect 323780 258046 324084 258074
rect 323780 253978 323808 258046
rect 323768 253972 323820 253978
rect 323768 253914 323820 253920
rect 323674 247616 323730 247625
rect 323674 247551 323730 247560
rect 323582 246256 323638 246265
rect 323582 246191 323638 246200
rect 322940 238128 322992 238134
rect 322940 238070 322992 238076
rect 323780 227594 323808 253914
rect 324148 252618 324176 312559
rect 323860 252612 323912 252618
rect 323860 252554 323912 252560
rect 324136 252612 324188 252618
rect 324136 252554 324188 252560
rect 323872 227662 323900 252554
rect 324240 249830 324268 313103
rect 324332 312497 324360 319738
rect 324594 319016 324650 319025
rect 324594 318951 324650 318960
rect 324502 318880 324558 318889
rect 324502 318815 324558 318824
rect 324412 318640 324464 318646
rect 324410 318608 324412 318617
rect 324464 318608 324466 318617
rect 324410 318543 324466 318552
rect 324412 315988 324464 315994
rect 324412 315930 324464 315936
rect 324318 312488 324374 312497
rect 324318 312423 324374 312432
rect 324424 308961 324452 315930
rect 324516 310185 324544 318815
rect 324608 318782 324636 318951
rect 324596 318776 324648 318782
rect 324596 318718 324648 318724
rect 324608 317762 324636 318718
rect 324700 318714 324728 319824
rect 324838 319784 324866 320076
rect 325560 320104 325616 320113
rect 324916 320039 324972 320048
rect 324792 319756 324866 319784
rect 324688 318708 324740 318714
rect 324688 318650 324740 318656
rect 324596 317756 324648 317762
rect 324596 317698 324648 317704
rect 324596 316056 324648 316062
rect 324596 315998 324648 316004
rect 324608 311681 324636 315998
rect 324792 315994 324820 319756
rect 324930 319716 324958 320039
rect 325114 319938 325142 320076
rect 325102 319932 325154 319938
rect 325102 319874 325154 319880
rect 325298 319784 325326 320076
rect 325390 319852 325418 320076
rect 326572 320104 326628 320113
rect 325560 320039 325616 320048
rect 325666 319938 325694 320076
rect 325654 319932 325706 319938
rect 325654 319874 325706 319880
rect 325758 319870 325786 320076
rect 325746 319864 325798 319870
rect 325390 319824 325464 319852
rect 325436 319818 325464 319824
rect 325436 319790 325648 319818
rect 325298 319756 325372 319784
rect 325148 319728 325200 319734
rect 324930 319688 325004 319716
rect 324976 317937 325004 319688
rect 325148 319670 325200 319676
rect 325054 318880 325110 318889
rect 325054 318815 325110 318824
rect 324962 317928 325018 317937
rect 324962 317863 325018 317872
rect 324964 317756 325016 317762
rect 324964 317698 325016 317704
rect 324872 316328 324924 316334
rect 324872 316270 324924 316276
rect 324780 315988 324832 315994
rect 324780 315930 324832 315936
rect 324884 311894 324912 316270
rect 324792 311866 324912 311894
rect 324594 311672 324650 311681
rect 324594 311607 324650 311616
rect 324502 310176 324558 310185
rect 324502 310111 324558 310120
rect 324410 308952 324466 308961
rect 324410 308887 324466 308896
rect 324792 306374 324820 311866
rect 324976 309369 325004 317698
rect 325068 317393 325096 318815
rect 325054 317384 325110 317393
rect 325054 317319 325110 317328
rect 325160 316062 325188 319670
rect 325344 319648 325372 319756
rect 325344 319620 325464 319648
rect 325330 319560 325386 319569
rect 325330 319495 325386 319504
rect 325148 316056 325200 316062
rect 325148 315998 325200 316004
rect 325344 314537 325372 319495
rect 325330 314528 325386 314537
rect 325330 314463 325386 314472
rect 325344 311894 325372 314463
rect 325436 314401 325464 319620
rect 325514 318744 325570 318753
rect 325514 318679 325570 318688
rect 325422 314392 325478 314401
rect 325422 314327 325478 314336
rect 325252 311866 325372 311894
rect 325146 311672 325202 311681
rect 325146 311607 325202 311616
rect 325054 310176 325110 310185
rect 325054 310111 325110 310120
rect 324962 309360 325018 309369
rect 324962 309295 325018 309304
rect 324792 306346 325004 306374
rect 324228 249824 324280 249830
rect 324228 249766 324280 249772
rect 324976 242214 325004 306346
rect 325068 250481 325096 310111
rect 325160 271153 325188 311607
rect 325252 284986 325280 311866
rect 325436 287706 325464 314327
rect 325424 287700 325476 287706
rect 325424 287642 325476 287648
rect 325240 284980 325292 284986
rect 325240 284922 325292 284928
rect 325146 271144 325202 271153
rect 325146 271079 325202 271088
rect 325148 266416 325200 266422
rect 325148 266358 325200 266364
rect 325054 250472 325110 250481
rect 325054 250407 325110 250416
rect 324964 242208 325016 242214
rect 324964 242150 325016 242156
rect 325160 228682 325188 266358
rect 325528 245041 325556 318679
rect 325620 317422 325648 319790
rect 325712 319812 325746 319818
rect 325712 319806 325798 319812
rect 325712 319790 325786 319806
rect 325608 317416 325660 317422
rect 325608 317358 325660 317364
rect 325620 316334 325648 317358
rect 325608 316328 325660 316334
rect 325608 316270 325660 316276
rect 325606 308952 325662 308961
rect 325606 308887 325662 308896
rect 325620 266422 325648 308887
rect 325608 266416 325660 266422
rect 325608 266358 325660 266364
rect 325712 246401 325740 319790
rect 325850 319716 325878 320076
rect 325804 319688 325878 319716
rect 325804 318794 325832 319688
rect 325942 319546 325970 320076
rect 326034 319716 326062 320076
rect 326126 319818 326154 320076
rect 326218 319920 326246 320076
rect 326218 319892 326292 319920
rect 326126 319790 326200 319818
rect 326034 319688 326108 319716
rect 325942 319518 326016 319546
rect 325804 318766 325924 318794
rect 325896 318209 325924 318766
rect 325882 318200 325938 318209
rect 325882 318135 325938 318144
rect 325882 317928 325938 317937
rect 325882 317863 325938 317872
rect 325792 317620 325844 317626
rect 325792 317562 325844 317568
rect 325804 311273 325832 317562
rect 325896 317529 325924 317863
rect 325882 317520 325938 317529
rect 325882 317455 325938 317464
rect 325988 316810 326016 319518
rect 325976 316804 326028 316810
rect 325976 316746 326028 316752
rect 326080 315897 326108 319688
rect 326172 317286 326200 319790
rect 326264 317529 326292 319892
rect 326402 319784 326430 320076
rect 326940 320104 326996 320113
rect 326572 320039 326628 320048
rect 326678 319920 326706 320076
rect 326678 319892 326752 319920
rect 326402 319756 326476 319784
rect 326250 317520 326306 317529
rect 326250 317455 326306 317464
rect 326160 317280 326212 317286
rect 326160 317222 326212 317228
rect 326066 315888 326122 315897
rect 326066 315823 326122 315832
rect 326080 311894 326108 315823
rect 326448 314265 326476 319756
rect 326724 319666 326752 319892
rect 326862 319852 326890 320076
rect 326940 320039 326996 320048
rect 326816 319824 326890 319852
rect 326528 319660 326580 319666
rect 326528 319602 326580 319608
rect 326712 319660 326764 319666
rect 326712 319602 326764 319608
rect 326540 317626 326568 319602
rect 326618 319560 326674 319569
rect 326618 319495 326674 319504
rect 326528 317620 326580 317626
rect 326528 317562 326580 317568
rect 326526 317384 326582 317393
rect 326526 317319 326582 317328
rect 326540 315761 326568 317319
rect 326526 315752 326582 315761
rect 326526 315687 326582 315696
rect 326434 314256 326490 314265
rect 326434 314191 326490 314200
rect 326526 313032 326582 313041
rect 326526 312967 326582 312976
rect 326080 311866 326384 311894
rect 325790 311264 325846 311273
rect 325790 311199 325846 311208
rect 325698 246392 325754 246401
rect 325698 246327 325754 246336
rect 325514 245032 325570 245041
rect 325514 244967 325570 244976
rect 326356 244905 326384 311866
rect 326434 310448 326490 310457
rect 326434 310383 326490 310392
rect 326448 247761 326476 310383
rect 326540 250617 326568 312967
rect 326632 312905 326660 319495
rect 326816 317529 326844 319824
rect 327046 319784 327074 320076
rect 327138 319938 327166 320076
rect 327126 319932 327178 319938
rect 327126 319874 327178 319880
rect 326908 319756 327074 319784
rect 326802 317520 326858 317529
rect 326802 317455 326858 317464
rect 326908 313041 326936 319756
rect 327138 319682 327166 319874
rect 327230 319784 327258 320076
rect 327552 320074 327580 330375
rect 327632 321904 327684 321910
rect 327632 321846 327684 321852
rect 327644 320793 327672 321846
rect 327736 321314 327764 359343
rect 327814 358048 327870 358057
rect 327814 357983 327870 357992
rect 327828 321570 327856 357983
rect 327906 351112 327962 351121
rect 327906 351047 327962 351056
rect 327816 321564 327868 321570
rect 327816 321506 327868 321512
rect 327920 321434 327948 351047
rect 327908 321428 327960 321434
rect 327908 321370 327960 321376
rect 327736 321286 327948 321314
rect 327724 321224 327776 321230
rect 327724 321166 327776 321172
rect 327630 320784 327686 320793
rect 327736 320754 327764 321166
rect 327630 320719 327686 320728
rect 327724 320748 327776 320754
rect 327724 320690 327776 320696
rect 327722 320648 327778 320657
rect 327644 320606 327722 320634
rect 327540 320068 327592 320074
rect 327540 320010 327592 320016
rect 327538 319968 327594 319977
rect 327538 319903 327594 319912
rect 327552 319818 327580 319903
rect 327644 319870 327672 320606
rect 327722 320583 327778 320592
rect 327722 320512 327778 320521
rect 327722 320447 327778 320456
rect 327736 320142 327764 320447
rect 327816 320272 327868 320278
rect 327816 320214 327868 320220
rect 327724 320136 327776 320142
rect 327724 320078 327776 320084
rect 327722 319968 327778 319977
rect 327722 319903 327778 319912
rect 327368 319790 327580 319818
rect 327632 319864 327684 319870
rect 327632 319806 327684 319812
rect 327230 319756 327304 319784
rect 327092 319654 327166 319682
rect 326986 319560 327042 319569
rect 326986 319495 327042 319504
rect 327000 316713 327028 319495
rect 326986 316704 327042 316713
rect 326986 316639 327042 316648
rect 326894 313032 326950 313041
rect 326894 312967 326950 312976
rect 326618 312896 326674 312905
rect 326618 312831 326674 312840
rect 326632 311894 326660 312831
rect 326632 311866 326752 311894
rect 326724 264217 326752 311866
rect 326986 311536 327042 311545
rect 326986 311471 327042 311480
rect 327000 311273 327028 311471
rect 326986 311264 327042 311273
rect 326986 311199 327042 311208
rect 326710 264208 326766 264217
rect 326710 264143 326766 264152
rect 327092 257281 327120 319654
rect 327276 318617 327304 319756
rect 327262 318608 327318 318617
rect 327262 318543 327318 318552
rect 327368 317937 327396 319790
rect 327446 319560 327502 319569
rect 327446 319495 327502 319504
rect 327354 317928 327410 317937
rect 327354 317863 327410 317872
rect 327460 317801 327488 319495
rect 327736 319433 327764 319903
rect 327828 319666 327856 320214
rect 327816 319660 327868 319666
rect 327816 319602 327868 319608
rect 327722 319424 327778 319433
rect 327722 319359 327778 319368
rect 327920 318374 327948 321286
rect 327908 318368 327960 318374
rect 327908 318310 327960 318316
rect 327540 318232 327592 318238
rect 327540 318174 327592 318180
rect 327446 317792 327502 317801
rect 327446 317727 327502 317736
rect 327446 317656 327502 317665
rect 327446 317591 327448 317600
rect 327500 317591 327502 317600
rect 327448 317562 327500 317568
rect 327262 316296 327318 316305
rect 327262 316231 327318 316240
rect 327172 309256 327224 309262
rect 327172 309198 327224 309204
rect 327078 257272 327134 257281
rect 327078 257207 327134 257216
rect 326526 250608 326582 250617
rect 326526 250543 326582 250552
rect 326434 247752 326490 247761
rect 326434 247687 326490 247696
rect 326342 244896 326398 244905
rect 326342 244831 326398 244840
rect 327184 229945 327212 309198
rect 327276 303521 327304 316231
rect 327460 308553 327488 317562
rect 327552 309262 327580 318174
rect 327816 317484 327868 317490
rect 327816 317426 327868 317432
rect 327828 315178 327856 317426
rect 327906 317384 327962 317393
rect 327906 317319 327962 317328
rect 327724 315172 327776 315178
rect 327724 315114 327776 315120
rect 327816 315172 327868 315178
rect 327816 315114 327868 315120
rect 327736 310418 327764 315114
rect 327816 314696 327868 314702
rect 327816 314638 327868 314644
rect 327724 310412 327776 310418
rect 327724 310354 327776 310360
rect 327540 309256 327592 309262
rect 327540 309198 327592 309204
rect 327446 308544 327502 308553
rect 327446 308479 327502 308488
rect 327262 303512 327318 303521
rect 327262 303447 327318 303456
rect 327264 277432 327316 277438
rect 327264 277374 327316 277380
rect 327170 229936 327226 229945
rect 327170 229871 327226 229880
rect 327276 228954 327304 277374
rect 327264 228948 327316 228954
rect 327264 228890 327316 228896
rect 325148 228676 325200 228682
rect 325148 228618 325200 228624
rect 323860 227656 323912 227662
rect 323860 227598 323912 227604
rect 323768 227588 323820 227594
rect 323768 227530 323820 227536
rect 321652 227520 321704 227526
rect 321652 227462 321704 227468
rect 327736 204270 327764 310354
rect 327828 225865 327856 314638
rect 327920 228818 327948 317319
rect 328012 309534 328040 395150
rect 329196 384396 329248 384402
rect 329196 384338 329248 384344
rect 328368 372088 328420 372094
rect 328368 372030 328420 372036
rect 328380 365673 328408 372030
rect 328366 365664 328422 365673
rect 328366 365599 328422 365608
rect 329104 363656 329156 363662
rect 329104 363598 329156 363604
rect 329012 329112 329064 329118
rect 329012 329054 329064 329060
rect 328182 323640 328238 323649
rect 328182 323575 328238 323584
rect 328092 321564 328144 321570
rect 328092 321506 328144 321512
rect 328104 318345 328132 321506
rect 328090 318336 328146 318345
rect 328090 318271 328146 318280
rect 328196 315858 328224 323575
rect 328366 321464 328422 321473
rect 328276 321428 328328 321434
rect 328366 321399 328422 321408
rect 328276 321370 328328 321376
rect 328288 318238 328316 321370
rect 328380 320521 328408 321399
rect 328366 320512 328422 320521
rect 328366 320447 328422 320456
rect 328368 320204 328420 320210
rect 328368 320146 328420 320152
rect 328380 319734 328408 320146
rect 328368 319728 328420 319734
rect 328368 319670 328420 319676
rect 328366 319016 328422 319025
rect 328366 318951 328422 318960
rect 328276 318232 328328 318238
rect 328276 318174 328328 318180
rect 328274 318064 328330 318073
rect 328274 317999 328330 318008
rect 328288 316878 328316 317999
rect 328276 316872 328328 316878
rect 328276 316814 328328 316820
rect 328184 315852 328236 315858
rect 328184 315794 328236 315800
rect 328288 314702 328316 316814
rect 328276 314696 328328 314702
rect 328276 314638 328328 314644
rect 328380 312662 328408 318951
rect 329024 318782 329052 329054
rect 329012 318776 329064 318782
rect 329012 318718 329064 318724
rect 328736 318368 328788 318374
rect 328736 318310 328788 318316
rect 328552 318300 328604 318306
rect 328552 318242 328604 318248
rect 328460 318232 328512 318238
rect 328460 318174 328512 318180
rect 328472 317218 328500 318174
rect 328460 317212 328512 317218
rect 328460 317154 328512 317160
rect 328564 317150 328592 318242
rect 328644 318164 328696 318170
rect 328644 318106 328696 318112
rect 328552 317144 328604 317150
rect 328552 317086 328604 317092
rect 328552 316940 328604 316946
rect 328552 316882 328604 316888
rect 328458 315752 328514 315761
rect 328458 315687 328514 315696
rect 328472 315314 328500 315687
rect 328460 315308 328512 315314
rect 328460 315250 328512 315256
rect 328368 312656 328420 312662
rect 328368 312598 328420 312604
rect 328458 311128 328514 311137
rect 328458 311063 328514 311072
rect 328000 309528 328052 309534
rect 328000 309470 328052 309476
rect 327908 228812 327960 228818
rect 327908 228754 327960 228760
rect 327814 225856 327870 225865
rect 327814 225791 327870 225800
rect 328472 223281 328500 311063
rect 328564 232558 328592 316882
rect 328656 315926 328684 318106
rect 328644 315920 328696 315926
rect 328644 315862 328696 315868
rect 328644 315172 328696 315178
rect 328644 315114 328696 315120
rect 328656 235414 328684 315114
rect 328748 314770 328776 318310
rect 329116 317626 329144 363598
rect 329104 317620 329156 317626
rect 329104 317562 329156 317568
rect 328828 317552 328880 317558
rect 328828 317494 328880 317500
rect 328840 317150 328868 317494
rect 329104 317348 329156 317354
rect 329104 317290 329156 317296
rect 328828 317144 328880 317150
rect 328828 317086 328880 317092
rect 328918 315752 328974 315761
rect 328918 315687 328974 315696
rect 328828 315308 328880 315314
rect 328828 315250 328880 315256
rect 328736 314764 328788 314770
rect 328736 314706 328788 314712
rect 328840 311894 328868 315250
rect 328932 315217 328960 315687
rect 328918 315208 328974 315217
rect 328918 315143 328974 315152
rect 328748 311866 328868 311894
rect 328748 237969 328776 311866
rect 328828 289128 328880 289134
rect 328828 289070 328880 289076
rect 328734 237960 328790 237969
rect 328734 237895 328790 237904
rect 328644 235408 328696 235414
rect 328644 235350 328696 235356
rect 328552 232552 328604 232558
rect 328552 232494 328604 232500
rect 328840 230489 328868 289070
rect 329116 235346 329144 317290
rect 329208 302870 329236 384338
rect 329300 314634 329328 395626
rect 330484 392556 330536 392562
rect 330484 392498 330536 392504
rect 329380 387524 329432 387530
rect 329380 387466 329432 387472
rect 329392 316470 329420 387466
rect 329472 387320 329524 387326
rect 329472 387262 329524 387268
rect 329380 316464 329432 316470
rect 329380 316406 329432 316412
rect 329484 316402 329512 387262
rect 329656 372156 329708 372162
rect 329656 372098 329708 372104
rect 329668 365702 329696 372098
rect 329748 367804 329800 367810
rect 329748 367746 329800 367752
rect 329656 365696 329708 365702
rect 329656 365638 329708 365644
rect 329564 334620 329616 334626
rect 329564 334562 329616 334568
rect 329576 317937 329604 334562
rect 329656 326392 329708 326398
rect 329656 326334 329708 326340
rect 329562 317928 329618 317937
rect 329562 317863 329618 317872
rect 329668 316946 329696 326334
rect 329760 318714 329788 367746
rect 330392 354000 330444 354006
rect 330392 353942 330444 353948
rect 330404 325694 330432 353942
rect 330220 325666 330432 325694
rect 330220 318782 330248 325666
rect 330392 322924 330444 322930
rect 330392 322866 330444 322872
rect 330404 321881 330432 322866
rect 330390 321872 330446 321881
rect 330390 321807 330446 321816
rect 329840 318776 329892 318782
rect 330208 318776 330260 318782
rect 329840 318718 329892 318724
rect 330114 318744 330170 318753
rect 329748 318708 329800 318714
rect 329748 318650 329800 318656
rect 329852 318646 329880 318718
rect 330208 318718 330260 318724
rect 330114 318679 330170 318688
rect 329840 318640 329892 318646
rect 329840 318582 329892 318588
rect 330024 318640 330076 318646
rect 330024 318582 330076 318588
rect 329930 318200 329986 318209
rect 329930 318135 329986 318144
rect 329838 318064 329894 318073
rect 329838 317999 329894 318008
rect 329748 317144 329800 317150
rect 329748 317086 329800 317092
rect 329656 316940 329708 316946
rect 329656 316882 329708 316888
rect 329472 316396 329524 316402
rect 329472 316338 329524 316344
rect 329288 314628 329340 314634
rect 329288 314570 329340 314576
rect 329760 313698 329788 317086
rect 329852 313886 329880 317999
rect 329840 313880 329892 313886
rect 329840 313822 329892 313828
rect 329760 313670 329880 313698
rect 329852 312882 329880 313670
rect 329944 313070 329972 318135
rect 330036 318102 330064 318582
rect 330024 318096 330076 318102
rect 330024 318038 330076 318044
rect 330128 317354 330156 318679
rect 330116 317348 330168 317354
rect 330116 317290 330168 317296
rect 330114 316704 330170 316713
rect 330114 316639 330170 316648
rect 330022 314256 330078 314265
rect 330022 314191 330078 314200
rect 330036 314022 330064 314191
rect 330024 314016 330076 314022
rect 330024 313958 330076 313964
rect 329932 313064 329984 313070
rect 329932 313006 329984 313012
rect 329852 312854 329972 312882
rect 329840 312792 329892 312798
rect 329840 312734 329892 312740
rect 329196 302864 329248 302870
rect 329196 302806 329248 302812
rect 329104 235340 329156 235346
rect 329104 235282 329156 235288
rect 329852 230994 329880 312734
rect 329944 235958 329972 312854
rect 330036 236638 330064 313958
rect 330128 307193 330156 316639
rect 330206 314528 330262 314537
rect 330206 314463 330262 314472
rect 330220 314265 330248 314463
rect 330206 314256 330262 314265
rect 330206 314191 330262 314200
rect 330392 310208 330444 310214
rect 330392 310150 330444 310156
rect 330404 309466 330432 310150
rect 330392 309460 330444 309466
rect 330392 309402 330444 309408
rect 330114 307184 330170 307193
rect 330114 307119 330170 307128
rect 330496 305726 330524 392498
rect 330588 313206 330616 395694
rect 330680 313682 330708 397190
rect 330772 319598 330800 398618
rect 330942 398440 330998 398449
rect 330942 398375 330998 398384
rect 330852 397588 330904 397594
rect 330852 397530 330904 397536
rect 330760 319592 330812 319598
rect 330760 319534 330812 319540
rect 330864 319530 330892 397530
rect 330852 319524 330904 319530
rect 330852 319466 330904 319472
rect 330956 318850 330984 398375
rect 331036 387592 331088 387598
rect 331036 387534 331088 387540
rect 330944 318844 330996 318850
rect 330944 318786 330996 318792
rect 330760 318096 330812 318102
rect 330760 318038 330812 318044
rect 330668 313676 330720 313682
rect 330668 313618 330720 313624
rect 330576 313200 330628 313206
rect 330576 313142 330628 313148
rect 330772 311001 330800 318038
rect 330850 314664 330906 314673
rect 330850 314599 330906 314608
rect 330864 313857 330892 314599
rect 330850 313848 330906 313857
rect 330850 313783 330906 313792
rect 330956 312798 330984 318786
rect 331048 312934 331076 387534
rect 331220 372020 331272 372026
rect 331220 371962 331272 371968
rect 331232 371278 331260 371962
rect 331220 371272 331272 371278
rect 331220 371214 331272 371220
rect 331680 371272 331732 371278
rect 331680 371214 331732 371220
rect 331128 359508 331180 359514
rect 331128 359450 331180 359456
rect 331140 318646 331168 359450
rect 331220 323604 331272 323610
rect 331220 323546 331272 323552
rect 331232 322969 331260 323546
rect 331218 322960 331274 322969
rect 331218 322895 331274 322904
rect 331312 322856 331364 322862
rect 331312 322798 331364 322804
rect 331324 322153 331352 322798
rect 331310 322144 331366 322153
rect 331310 322079 331366 322088
rect 331220 318776 331272 318782
rect 331220 318718 331272 318724
rect 331128 318640 331180 318646
rect 331128 318582 331180 318588
rect 331036 312928 331088 312934
rect 331036 312870 331088 312876
rect 330944 312792 330996 312798
rect 330944 312734 330996 312740
rect 330758 310992 330814 311001
rect 330758 310927 330814 310936
rect 330484 305720 330536 305726
rect 330484 305662 330536 305668
rect 330024 236632 330076 236638
rect 330024 236574 330076 236580
rect 329932 235952 329984 235958
rect 329932 235894 329984 235900
rect 329840 230988 329892 230994
rect 329840 230930 329892 230936
rect 328826 230480 328882 230489
rect 328826 230415 328882 230424
rect 331232 229809 331260 318718
rect 331324 235249 331352 322079
rect 331496 318708 331548 318714
rect 331496 318650 331548 318656
rect 331402 318608 331458 318617
rect 331402 318543 331458 318552
rect 331416 318034 331444 318543
rect 331404 318028 331456 318034
rect 331404 317970 331456 317976
rect 331416 235929 331444 317970
rect 331402 235920 331458 235929
rect 331402 235855 331458 235864
rect 331508 235482 331536 318650
rect 331588 315376 331640 315382
rect 331588 315318 331640 315324
rect 331496 235476 331548 235482
rect 331496 235418 331548 235424
rect 331600 235278 331628 315318
rect 331692 291854 331720 371214
rect 331772 323604 331824 323610
rect 331772 323546 331824 323552
rect 331784 300121 331812 323546
rect 331876 307290 331904 399638
rect 331954 395992 332010 396001
rect 331954 395927 332010 395936
rect 331968 308310 331996 395927
rect 332060 371210 332088 455738
rect 332048 371204 332100 371210
rect 332048 371146 332100 371152
rect 332152 370802 332180 455806
rect 333336 455728 333388 455734
rect 333336 455670 333388 455676
rect 332232 455660 332284 455666
rect 332232 455602 332284 455608
rect 332244 371958 332272 455602
rect 333244 397792 333296 397798
rect 333244 397734 333296 397740
rect 333256 397662 333284 397734
rect 333244 397656 333296 397662
rect 333244 397598 333296 397604
rect 332324 397316 332376 397322
rect 332324 397258 332376 397264
rect 332232 371952 332284 371958
rect 332232 371894 332284 371900
rect 332140 370796 332192 370802
rect 332140 370738 332192 370744
rect 332048 349852 332100 349858
rect 332048 349794 332100 349800
rect 332060 318442 332088 349794
rect 332140 348424 332192 348430
rect 332140 348366 332192 348372
rect 332048 318436 332100 318442
rect 332048 318378 332100 318384
rect 332152 317898 332180 348366
rect 332232 342916 332284 342922
rect 332232 342858 332284 342864
rect 332140 317892 332192 317898
rect 332140 317834 332192 317840
rect 332244 317830 332272 342858
rect 332232 317824 332284 317830
rect 332232 317766 332284 317772
rect 332336 314158 332364 397258
rect 333242 397216 333298 397225
rect 333242 397151 333298 397160
rect 332416 387388 332468 387394
rect 332416 387330 332468 387336
rect 332428 314906 332456 387330
rect 332692 372088 332744 372094
rect 332692 372030 332744 372036
rect 332600 371952 332652 371958
rect 332600 371894 332652 371900
rect 332612 371346 332640 371894
rect 332704 371414 332732 372030
rect 332692 371408 332744 371414
rect 332692 371350 332744 371356
rect 332600 371340 332652 371346
rect 332600 371282 332652 371288
rect 332704 354674 332732 371350
rect 332968 371340 333020 371346
rect 332968 371282 333020 371288
rect 332612 354646 332732 354674
rect 332416 314900 332468 314906
rect 332416 314842 332468 314848
rect 332324 314152 332376 314158
rect 332324 314094 332376 314100
rect 332612 308514 332640 354646
rect 332692 322244 332744 322250
rect 332692 322186 332744 322192
rect 332704 322017 332732 322186
rect 332690 322008 332746 322017
rect 332746 321966 332824 321994
rect 332690 321943 332746 321952
rect 332692 321292 332744 321298
rect 332692 321234 332744 321240
rect 332704 320210 332732 321234
rect 332692 320204 332744 320210
rect 332692 320146 332744 320152
rect 332600 308508 332652 308514
rect 332600 308450 332652 308456
rect 331956 308304 332008 308310
rect 331956 308246 332008 308252
rect 331864 307284 331916 307290
rect 331864 307226 331916 307232
rect 331770 300112 331826 300121
rect 331770 300047 331826 300056
rect 331680 291848 331732 291854
rect 331680 291790 331732 291796
rect 331588 235272 331640 235278
rect 331310 235240 331366 235249
rect 331588 235214 331640 235220
rect 331310 235175 331366 235184
rect 332704 231130 332732 320146
rect 332796 238785 332824 321966
rect 332876 317280 332928 317286
rect 332876 317222 332928 317228
rect 332782 238776 332838 238785
rect 332782 238711 332838 238720
rect 332888 236774 332916 317222
rect 332980 308582 333008 371282
rect 333060 318640 333112 318646
rect 333060 318582 333112 318588
rect 332968 308576 333020 308582
rect 332968 308518 333020 308524
rect 332876 236768 332928 236774
rect 332876 236710 332928 236716
rect 332692 231124 332744 231130
rect 332692 231066 332744 231072
rect 331218 229800 331274 229809
rect 331218 229735 331274 229744
rect 333072 227118 333100 318582
rect 333152 312656 333204 312662
rect 333152 312598 333204 312604
rect 333164 237289 333192 312598
rect 333256 311846 333284 397151
rect 333348 370938 333376 455670
rect 333428 455592 333480 455598
rect 333428 455534 333480 455540
rect 333440 372094 333468 455534
rect 333886 450256 333942 450265
rect 333886 450191 333942 450200
rect 333520 388748 333572 388754
rect 333520 388690 333572 388696
rect 333428 372088 333480 372094
rect 333428 372030 333480 372036
rect 333336 370932 333388 370938
rect 333336 370874 333388 370880
rect 333336 358080 333388 358086
rect 333336 358022 333388 358028
rect 333348 318578 333376 358022
rect 333428 355360 333480 355366
rect 333428 355302 333480 355308
rect 333336 318572 333388 318578
rect 333336 318514 333388 318520
rect 333440 317694 333468 355302
rect 333428 317688 333480 317694
rect 333428 317630 333480 317636
rect 333244 311840 333296 311846
rect 333244 311782 333296 311788
rect 333532 310486 333560 388690
rect 333612 387456 333664 387462
rect 333612 387398 333664 387404
rect 333624 314566 333652 387398
rect 333900 369034 333928 450191
rect 334162 398576 334218 398585
rect 334162 398511 334218 398520
rect 334176 398313 334204 398511
rect 334162 398304 334218 398313
rect 334162 398239 334218 398248
rect 334636 370666 334664 455874
rect 334728 401606 334756 457234
rect 355336 456794 355364 484366
rect 356704 472660 356756 472666
rect 356704 472602 356756 472608
rect 355968 456816 356020 456822
rect 355336 456766 355548 456794
rect 355520 455938 355548 456766
rect 355968 456758 356020 456764
rect 355508 455932 355560 455938
rect 355508 455874 355560 455880
rect 351920 454980 351972 454986
rect 351920 454922 351972 454928
rect 337936 454776 337988 454782
rect 337936 454718 337988 454724
rect 337292 454708 337344 454714
rect 337292 454650 337344 454656
rect 336464 454164 336516 454170
rect 336464 454106 336516 454112
rect 335268 453484 335320 453490
rect 335268 453426 335320 453432
rect 335176 453280 335228 453286
rect 335176 453222 335228 453228
rect 334806 452704 334862 452713
rect 334806 452639 334862 452648
rect 334820 405618 334848 452639
rect 334808 405612 334860 405618
rect 334808 405554 334860 405560
rect 334716 401600 334768 401606
rect 334716 401542 334768 401548
rect 334992 399084 335044 399090
rect 334992 399026 335044 399032
rect 334716 397452 334768 397458
rect 334716 397394 334768 397400
rect 334624 370660 334676 370666
rect 334624 370602 334676 370608
rect 333888 369028 333940 369034
rect 333888 368970 333940 368976
rect 334624 369028 334676 369034
rect 334624 368970 334676 368976
rect 333900 368801 333928 368970
rect 333886 368792 333942 368801
rect 333886 368727 333942 368736
rect 333704 333260 333756 333266
rect 333704 333202 333756 333208
rect 333716 317286 333744 333202
rect 333980 325100 334032 325106
rect 333980 325042 334032 325048
rect 333992 319977 334020 325042
rect 333978 319968 334034 319977
rect 333978 319903 334034 319912
rect 333704 317280 333756 317286
rect 333704 317222 333756 317228
rect 333612 314560 333664 314566
rect 333612 314502 333664 314508
rect 333520 310480 333572 310486
rect 333520 310422 333572 310428
rect 333150 237280 333206 237289
rect 333150 237215 333206 237224
rect 333992 227633 334020 319903
rect 334072 307692 334124 307698
rect 334072 307634 334124 307640
rect 334084 233073 334112 307634
rect 334070 233064 334126 233073
rect 334070 232999 334126 233008
rect 333978 227624 334034 227633
rect 333978 227559 334034 227568
rect 333060 227112 333112 227118
rect 333060 227054 333112 227060
rect 328458 223272 328514 223281
rect 328458 223207 328514 223216
rect 327724 204264 327776 204270
rect 327724 204206 327776 204212
rect 327080 149796 327132 149802
rect 327080 149738 327132 149744
rect 323584 141500 323636 141506
rect 323584 141442 323636 141448
rect 322938 68232 322994 68241
rect 322938 68167 322994 68176
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 315396 4140 315448 4146
rect 315396 4082 315448 4088
rect 316040 4140 316092 4146
rect 316040 4082 316092 4088
rect 316684 4140 316736 4146
rect 316684 4082 316736 4088
rect 314016 4072 314068 4078
rect 314016 4014 314068 4020
rect 314016 3868 314068 3874
rect 314016 3810 314068 3816
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 313924 3528 313976 3534
rect 313924 3470 313976 3476
rect 312648 480 312676 3470
rect 313832 3392 313884 3398
rect 313832 3334 313884 3340
rect 313844 480 313872 3334
rect 314028 3262 314056 3810
rect 314016 3256 314068 3262
rect 314016 3198 314068 3204
rect 315028 3052 315080 3058
rect 315028 2994 315080 3000
rect 315040 480 315068 2994
rect 316052 2122 316080 4082
rect 317328 4004 317380 4010
rect 317328 3946 317380 3952
rect 316052 2094 316264 2122
rect 316236 480 316264 2094
rect 317340 480 317368 3946
rect 318524 3256 318576 3262
rect 318524 3198 318576 3204
rect 318536 480 318564 3198
rect 319732 480 319760 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 320824 3596 320876 3602
rect 320824 3538 320876 3544
rect 320836 3398 320864 3538
rect 320824 3392 320876 3398
rect 320824 3334 320876 3340
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 68167
rect 323596 3874 323624 141442
rect 327092 16574 327120 149738
rect 327092 16546 327672 16574
rect 323676 4140 323728 4146
rect 323676 4082 323728 4088
rect 323688 3942 323716 4082
rect 326804 4072 326856 4078
rect 326804 4014 326856 4020
rect 325608 4004 325660 4010
rect 325608 3946 325660 3952
rect 323676 3936 323728 3942
rect 323676 3878 323728 3884
rect 323584 3868 323636 3874
rect 323584 3810 323636 3816
rect 324412 3664 324464 3670
rect 324412 3606 324464 3612
rect 324424 480 324452 3606
rect 325620 480 325648 3946
rect 326816 480 326844 4014
rect 327644 3482 327672 16546
rect 327736 3670 327764 204206
rect 332690 102776 332746 102785
rect 332690 102711 332746 102720
rect 331864 72480 331916 72486
rect 331864 72422 331916 72428
rect 330392 4820 330444 4826
rect 330392 4762 330444 4768
rect 329196 3800 329248 3806
rect 329196 3742 329248 3748
rect 327724 3664 327776 3670
rect 327724 3606 327776 3612
rect 327644 3454 328040 3482
rect 328012 480 328040 3454
rect 329208 480 329236 3742
rect 330404 480 330432 4762
rect 331588 3936 331640 3942
rect 331588 3878 331640 3884
rect 331600 480 331628 3878
rect 331876 3194 331904 72422
rect 332600 3732 332652 3738
rect 332600 3674 332652 3680
rect 331864 3188 331916 3194
rect 331864 3130 331916 3136
rect 332612 762 332640 3674
rect 332704 3398 332732 102711
rect 334636 20670 334664 368970
rect 334728 304162 334756 397394
rect 334806 395856 334862 395865
rect 334806 395791 334862 395800
rect 334716 304156 334768 304162
rect 334716 304098 334768 304104
rect 334820 304094 334848 395791
rect 334900 394596 334952 394602
rect 334900 394538 334952 394544
rect 334912 305590 334940 394538
rect 335004 315382 335032 399026
rect 335084 396024 335136 396030
rect 335084 395966 335136 395972
rect 334992 315376 335044 315382
rect 334992 315318 335044 315324
rect 335096 312526 335124 395966
rect 335188 370870 335216 453222
rect 335176 370864 335228 370870
rect 335176 370806 335228 370812
rect 335280 370734 335308 453426
rect 335818 452160 335874 452169
rect 335818 452095 335874 452104
rect 335832 451761 335860 452095
rect 335818 451752 335874 451761
rect 335818 451687 335874 451696
rect 336002 449304 336058 449313
rect 336002 449239 336058 449248
rect 336016 448905 336044 449239
rect 336002 448896 336058 448905
rect 336002 448831 336058 448840
rect 336094 402248 336150 402257
rect 336094 402183 336150 402192
rect 336004 396568 336056 396574
rect 336004 396510 336056 396516
rect 335268 370728 335320 370734
rect 335268 370670 335320 370676
rect 335176 356720 335228 356726
rect 335176 356662 335228 356668
rect 335188 318481 335216 356662
rect 335912 331900 335964 331906
rect 335912 331842 335964 331848
rect 335266 329216 335322 329225
rect 335266 329151 335322 329160
rect 335174 318472 335230 318481
rect 335174 318407 335230 318416
rect 335084 312520 335136 312526
rect 335084 312462 335136 312468
rect 335280 307698 335308 329151
rect 335818 321328 335874 321337
rect 335818 321263 335874 321272
rect 335832 320249 335860 321263
rect 335450 320240 335506 320249
rect 335450 320175 335506 320184
rect 335818 320240 335874 320249
rect 335818 320175 335874 320184
rect 335358 316568 335414 316577
rect 335358 316503 335414 316512
rect 335268 307692 335320 307698
rect 335268 307634 335320 307640
rect 334900 305584 334952 305590
rect 334900 305526 334952 305532
rect 334808 304088 334860 304094
rect 334808 304030 334860 304036
rect 335372 229022 335400 316503
rect 335464 233170 335492 320175
rect 335924 316577 335952 331842
rect 335910 316568 335966 316577
rect 335910 316503 335966 316512
rect 336016 305794 336044 396510
rect 336108 311370 336136 402183
rect 336278 397624 336334 397633
rect 336278 397559 336334 397568
rect 336188 397112 336240 397118
rect 336188 397054 336240 397060
rect 336200 312594 336228 397054
rect 336292 313954 336320 397559
rect 336372 395820 336424 395826
rect 336372 395762 336424 395768
rect 336280 313948 336332 313954
rect 336280 313890 336332 313896
rect 336188 312588 336240 312594
rect 336188 312530 336240 312536
rect 336384 312322 336412 395762
rect 336476 371890 336504 454106
rect 336556 394528 336608 394534
rect 336556 394470 336608 394476
rect 336464 371884 336516 371890
rect 336464 371826 336516 371832
rect 336462 326496 336518 326505
rect 336462 326431 336518 326440
rect 336372 312316 336424 312322
rect 336372 312258 336424 312264
rect 336096 311364 336148 311370
rect 336096 311306 336148 311312
rect 336004 305788 336056 305794
rect 336004 305730 336056 305736
rect 336476 304337 336504 326431
rect 336568 315450 336596 394470
rect 336648 393100 336700 393106
rect 336648 393042 336700 393048
rect 336660 316674 336688 393042
rect 337304 377466 337332 454650
rect 337384 454640 337436 454646
rect 337384 454582 337436 454588
rect 337292 377460 337344 377466
rect 337292 377402 337344 377408
rect 337396 372570 337424 454582
rect 337476 454096 337528 454102
rect 337476 454038 337528 454044
rect 337488 413982 337516 454038
rect 337568 451512 337620 451518
rect 337568 451454 337620 451460
rect 337580 418810 337608 451454
rect 337568 418804 337620 418810
rect 337568 418746 337620 418752
rect 337476 413976 337528 413982
rect 337476 413918 337528 413924
rect 337752 399220 337804 399226
rect 337752 399162 337804 399168
rect 337474 397352 337530 397361
rect 337474 397287 337530 397296
rect 337384 372564 337436 372570
rect 337384 372506 337436 372512
rect 337382 368520 337438 368529
rect 337382 368455 337438 368464
rect 337292 326460 337344 326466
rect 337292 326402 337344 326408
rect 337200 325032 337252 325038
rect 337200 324974 337252 324980
rect 337212 320521 337240 324974
rect 336830 320512 336886 320521
rect 336830 320447 336886 320456
rect 337198 320512 337254 320521
rect 337198 320447 337254 320456
rect 336738 317112 336794 317121
rect 336738 317047 336794 317056
rect 336648 316668 336700 316674
rect 336648 316610 336700 316616
rect 336556 315444 336608 315450
rect 336556 315386 336608 315392
rect 335542 304328 335598 304337
rect 335542 304263 335598 304272
rect 336462 304328 336518 304337
rect 336462 304263 336518 304272
rect 335556 238066 335584 304263
rect 336372 291984 336424 291990
rect 336372 291926 336424 291932
rect 336384 291174 336412 291926
rect 336004 291168 336056 291174
rect 336004 291110 336056 291116
rect 336372 291168 336424 291174
rect 336372 291110 336424 291116
rect 335544 238060 335596 238066
rect 335544 238002 335596 238008
rect 335452 233164 335504 233170
rect 335452 233106 335504 233112
rect 335360 229016 335412 229022
rect 335360 228958 335412 228964
rect 336016 213246 336044 291110
rect 336752 222086 336780 317047
rect 336844 227322 336872 320447
rect 337304 316034 337332 326402
rect 336936 316006 337332 316034
rect 336936 315353 336964 316006
rect 336922 315344 336978 315353
rect 336922 315279 336978 315288
rect 336832 227316 336884 227322
rect 336832 227258 336884 227264
rect 336936 227050 336964 315279
rect 336924 227044 336976 227050
rect 336924 226986 336976 226992
rect 336740 222080 336792 222086
rect 336740 222022 336792 222028
rect 335360 213240 335412 213246
rect 335360 213182 335412 213188
rect 336004 213240 336056 213246
rect 336004 213182 336056 213188
rect 334624 20664 334676 20670
rect 334624 20606 334676 20612
rect 335372 16574 335400 213182
rect 337396 100706 337424 368455
rect 337488 302938 337516 397287
rect 337660 395276 337712 395282
rect 337660 395218 337712 395224
rect 337568 390244 337620 390250
rect 337568 390186 337620 390192
rect 337476 302932 337528 302938
rect 337476 302874 337528 302880
rect 337580 298994 337608 390186
rect 337672 307222 337700 395218
rect 337764 315586 337792 399162
rect 337844 397180 337896 397186
rect 337844 397122 337896 397128
rect 337752 315580 337804 315586
rect 337752 315522 337804 315528
rect 337856 315178 337884 397122
rect 337948 373454 337976 454718
rect 340696 454232 340748 454238
rect 340696 454174 340748 454180
rect 340052 452668 340104 452674
rect 340052 452610 340104 452616
rect 339408 451376 339460 451382
rect 339408 451318 339460 451324
rect 338856 451308 338908 451314
rect 338856 451250 338908 451256
rect 338764 450152 338816 450158
rect 338764 450094 338816 450100
rect 338028 399152 338080 399158
rect 338028 399094 338080 399100
rect 337936 373448 337988 373454
rect 337936 373390 337988 373396
rect 337934 327720 337990 327729
rect 337934 327655 337990 327664
rect 337948 317121 337976 327655
rect 338040 322862 338068 399094
rect 338672 384464 338724 384470
rect 338672 384406 338724 384412
rect 338118 325272 338174 325281
rect 338118 325207 338174 325216
rect 338028 322856 338080 322862
rect 338028 322798 338080 322804
rect 337934 317112 337990 317121
rect 337934 317047 337990 317056
rect 338132 316849 338160 325207
rect 338210 321736 338266 321745
rect 338210 321671 338266 321680
rect 338118 316840 338174 316849
rect 338118 316775 338174 316784
rect 337844 315172 337896 315178
rect 337844 315114 337896 315120
rect 337660 307216 337712 307222
rect 337660 307158 337712 307164
rect 337568 298988 337620 298994
rect 337568 298930 337620 298936
rect 338132 220794 338160 316775
rect 338224 229090 338252 321671
rect 338684 307766 338712 384406
rect 338776 368665 338804 450094
rect 338868 406502 338896 451250
rect 338856 406496 338908 406502
rect 338856 406438 338908 406444
rect 339132 398812 339184 398818
rect 339132 398754 339184 398760
rect 338948 397656 339000 397662
rect 338948 397598 339000 397604
rect 338854 394768 338910 394777
rect 338854 394703 338910 394712
rect 338762 368656 338818 368665
rect 338762 368591 338818 368600
rect 338672 307760 338724 307766
rect 338672 307702 338724 307708
rect 338212 229084 338264 229090
rect 338212 229026 338264 229032
rect 338120 220788 338172 220794
rect 338120 220730 338172 220736
rect 338776 193186 338804 368591
rect 338868 295186 338896 394703
rect 338960 309806 338988 397598
rect 339040 393440 339092 393446
rect 339040 393382 339092 393388
rect 338948 309800 339000 309806
rect 338948 309742 339000 309748
rect 339052 306066 339080 393382
rect 339144 311234 339172 398754
rect 339316 395616 339368 395622
rect 339316 395558 339368 395564
rect 339224 394460 339276 394466
rect 339224 394402 339276 394408
rect 339132 311228 339184 311234
rect 339132 311170 339184 311176
rect 339236 308242 339264 394402
rect 339328 317150 339356 395558
rect 339420 370666 339448 451318
rect 339868 400104 339920 400110
rect 339868 400046 339920 400052
rect 339880 396982 339908 400046
rect 339868 396976 339920 396982
rect 339868 396918 339920 396924
rect 339866 396264 339922 396273
rect 339866 396199 339922 396208
rect 339880 394262 339908 396199
rect 339868 394256 339920 394262
rect 339868 394198 339920 394204
rect 340064 373318 340092 452610
rect 340144 452056 340196 452062
rect 340144 451998 340196 452004
rect 340156 407794 340184 451998
rect 340234 451480 340290 451489
rect 340234 451415 340290 451424
rect 340248 409154 340276 451415
rect 340328 450016 340380 450022
rect 340328 449958 340380 449964
rect 340340 411262 340368 449958
rect 340328 411256 340380 411262
rect 340328 411198 340380 411204
rect 340236 409148 340288 409154
rect 340236 409090 340288 409096
rect 340144 407788 340196 407794
rect 340144 407730 340196 407736
rect 340328 399764 340380 399770
rect 340328 399706 340380 399712
rect 340340 398614 340368 399706
rect 340512 398948 340564 398954
rect 340512 398890 340564 398896
rect 340420 398880 340472 398886
rect 340420 398822 340472 398828
rect 340328 398608 340380 398614
rect 340328 398550 340380 398556
rect 340234 398304 340290 398313
rect 340234 398239 340290 398248
rect 340144 395888 340196 395894
rect 340144 395830 340196 395836
rect 340052 373312 340104 373318
rect 340052 373254 340104 373260
rect 339408 370660 339460 370666
rect 339408 370602 339460 370608
rect 339420 369986 339448 370602
rect 339408 369980 339460 369986
rect 339408 369922 339460 369928
rect 340050 365664 340106 365673
rect 340050 365599 340106 365608
rect 340064 364993 340092 365599
rect 340050 364984 340106 364993
rect 340050 364919 340106 364928
rect 339316 317144 339368 317150
rect 339316 317086 339368 317092
rect 339498 317112 339554 317121
rect 339498 317047 339554 317056
rect 339224 308236 339276 308242
rect 339224 308178 339276 308184
rect 339040 306060 339092 306066
rect 339040 306002 339092 306008
rect 338856 295180 338908 295186
rect 338856 295122 338908 295128
rect 339512 223553 339540 317047
rect 339592 305448 339644 305454
rect 339592 305390 339644 305396
rect 339604 305046 339632 305390
rect 339592 305040 339644 305046
rect 339592 304982 339644 304988
rect 339498 223544 339554 223553
rect 339498 223479 339554 223488
rect 339604 222193 339632 304982
rect 340156 300082 340184 395830
rect 340248 303006 340276 398239
rect 340326 396536 340382 396545
rect 340326 396471 340382 396480
rect 340340 304366 340368 396471
rect 340432 308378 340460 398822
rect 340524 309942 340552 398890
rect 340604 396772 340656 396778
rect 340604 396714 340656 396720
rect 340512 309936 340564 309942
rect 340512 309878 340564 309884
rect 340616 308446 340644 396714
rect 340708 373386 340736 454174
rect 350722 454064 350778 454073
rect 350722 453999 350778 454008
rect 341984 452736 342036 452742
rect 341984 452678 342036 452684
rect 341524 451716 341576 451722
rect 341524 451658 341576 451664
rect 340972 451648 341024 451654
rect 340972 451590 341024 451596
rect 340878 451344 340934 451353
rect 340878 451279 340934 451288
rect 340788 449948 340840 449954
rect 340788 449890 340840 449896
rect 340696 373380 340748 373386
rect 340696 373322 340748 373328
rect 340800 364993 340828 449890
rect 340892 435402 340920 451279
rect 340984 445058 341012 451590
rect 340972 445052 341024 445058
rect 340972 444994 341024 445000
rect 341536 441614 341564 451658
rect 341708 451444 341760 451450
rect 341708 451386 341760 451392
rect 341444 441586 341564 441614
rect 340970 438288 341026 438297
rect 340970 438223 341026 438232
rect 340984 438190 341012 438223
rect 340972 438184 341024 438190
rect 340972 438126 341024 438132
rect 340880 435396 340932 435402
rect 340880 435338 340932 435344
rect 341444 431954 341472 441586
rect 341720 438297 341748 451386
rect 341706 438288 341762 438297
rect 341706 438223 341762 438232
rect 341444 431926 341564 431954
rect 341536 412634 341564 431926
rect 340984 412606 341564 412634
rect 340984 404326 341012 412606
rect 340972 404320 341024 404326
rect 340972 404262 341024 404268
rect 341338 401840 341394 401849
rect 341338 401775 341394 401784
rect 341352 400178 341380 401775
rect 341800 400988 341852 400994
rect 341800 400930 341852 400936
rect 341432 400852 341484 400858
rect 341432 400794 341484 400800
rect 341524 400852 341576 400858
rect 341524 400794 341576 400800
rect 341444 400761 341472 400794
rect 341430 400752 341486 400761
rect 341430 400687 341486 400696
rect 341432 400376 341484 400382
rect 341432 400318 341484 400324
rect 341340 400172 341392 400178
rect 341340 400114 341392 400120
rect 341248 399696 341300 399702
rect 341248 399638 341300 399644
rect 341156 398132 341208 398138
rect 341156 398074 341208 398080
rect 340972 397520 341024 397526
rect 340972 397462 341024 397468
rect 340984 391513 341012 397462
rect 340970 391504 341026 391513
rect 340970 391439 341026 391448
rect 341168 390561 341196 398074
rect 341154 390552 341210 390561
rect 341154 390487 341210 390496
rect 341260 387258 341288 399638
rect 341444 398993 341472 400318
rect 341536 399974 341564 400794
rect 341614 400344 341670 400353
rect 341614 400279 341670 400288
rect 341628 400110 341656 400279
rect 341616 400104 341668 400110
rect 341616 400046 341668 400052
rect 341524 399968 341576 399974
rect 341524 399910 341576 399916
rect 341812 399634 341840 400930
rect 341892 400580 341944 400586
rect 341892 400522 341944 400528
rect 341904 400314 341932 400522
rect 341892 400308 341944 400314
rect 341892 400250 341944 400256
rect 341890 400208 341946 400217
rect 341890 400143 341946 400152
rect 341904 399809 341932 400143
rect 341890 399800 341946 399809
rect 341890 399735 341946 399744
rect 341800 399628 341852 399634
rect 341800 399570 341852 399576
rect 341430 398984 341486 398993
rect 341430 398919 341486 398928
rect 341890 398848 341946 398857
rect 341890 398783 341946 398792
rect 341904 398342 341932 398783
rect 341892 398336 341944 398342
rect 341892 398278 341944 398284
rect 341892 398064 341944 398070
rect 341892 398006 341944 398012
rect 341524 397860 341576 397866
rect 341524 397802 341576 397808
rect 341338 395720 341394 395729
rect 341338 395655 341394 395664
rect 341248 387252 341300 387258
rect 341248 387194 341300 387200
rect 340880 369844 340932 369850
rect 340880 369786 340932 369792
rect 340892 369170 340920 369786
rect 340880 369164 340932 369170
rect 340880 369106 340932 369112
rect 340786 364984 340842 364993
rect 340786 364919 340842 364928
rect 340694 337376 340750 337385
rect 340694 337311 340750 337320
rect 340708 317121 340736 337311
rect 340970 323776 341026 323785
rect 340788 323740 340840 323746
rect 340970 323711 341026 323720
rect 340788 323682 340840 323688
rect 340694 317112 340750 317121
rect 340694 317047 340750 317056
rect 340604 308440 340656 308446
rect 340604 308382 340656 308388
rect 340420 308372 340472 308378
rect 340420 308314 340472 308320
rect 340800 305046 340828 323682
rect 340880 317280 340932 317286
rect 340880 317222 340932 317228
rect 340892 317014 340920 317222
rect 340984 317082 341012 323711
rect 340972 317076 341024 317082
rect 340972 317018 341024 317024
rect 340880 317008 340932 317014
rect 340880 316950 340932 316956
rect 340788 305040 340840 305046
rect 340788 304982 340840 304988
rect 340328 304360 340380 304366
rect 340328 304302 340380 304308
rect 340236 303000 340288 303006
rect 340236 302942 340288 302948
rect 340144 300076 340196 300082
rect 340144 300018 340196 300024
rect 339590 222184 339646 222193
rect 339590 222119 339646 222128
rect 340892 220833 340920 316950
rect 340984 222154 341012 317018
rect 341352 316878 341380 395655
rect 341432 393168 341484 393174
rect 341432 393110 341484 393116
rect 341340 316872 341392 316878
rect 341340 316814 341392 316820
rect 341444 314090 341472 393110
rect 341432 314084 341484 314090
rect 341432 314026 341484 314032
rect 341536 295322 341564 397802
rect 341800 396160 341852 396166
rect 341800 396102 341852 396108
rect 341708 395956 341760 395962
rect 341708 395898 341760 395904
rect 341616 394664 341668 394670
rect 341616 394606 341668 394612
rect 341628 304230 341656 394606
rect 341720 310418 341748 395898
rect 341812 395350 341840 396102
rect 341800 395344 341852 395350
rect 341800 395286 341852 395292
rect 341800 393236 341852 393242
rect 341800 393178 341852 393184
rect 341812 392057 341840 393178
rect 341798 392048 341854 392057
rect 341798 391983 341854 391992
rect 341800 391060 341852 391066
rect 341800 391002 341852 391008
rect 341812 313002 341840 391002
rect 341904 314226 341932 398006
rect 341996 379030 342024 452678
rect 348516 452192 348568 452198
rect 344466 452160 344522 452169
rect 348516 452134 348568 452140
rect 344466 452095 344522 452104
rect 342168 451852 342220 451858
rect 342168 451794 342220 451800
rect 342076 449336 342128 449342
rect 342076 449278 342128 449284
rect 341984 379024 342036 379030
rect 341984 378966 342036 378972
rect 342088 378876 342116 449278
rect 341996 378848 342116 378876
rect 341996 369170 342024 378848
rect 342076 378752 342128 378758
rect 342076 378694 342128 378700
rect 342088 372638 342116 378694
rect 342076 372632 342128 372638
rect 342076 372574 342128 372580
rect 342088 370598 342116 372574
rect 342076 370592 342128 370598
rect 342076 370534 342128 370540
rect 341984 369164 342036 369170
rect 341984 369106 342036 369112
rect 342180 365702 342208 451794
rect 342352 451784 342404 451790
rect 342352 451726 342404 451732
rect 344098 451752 344154 451761
rect 342364 447134 342392 451726
rect 344098 451687 344154 451696
rect 344112 449970 344140 451687
rect 344480 449970 344508 452095
rect 345202 452024 345258 452033
rect 345202 451959 345258 451968
rect 345064 450256 345120 450265
rect 345064 450191 345120 450200
rect 344112 449942 344356 449970
rect 344480 449942 344724 449970
rect 345078 449956 345106 450191
rect 345216 449970 345244 451959
rect 347778 451888 347834 451897
rect 347778 451823 347834 451832
rect 345938 451480 345994 451489
rect 345938 451415 345994 451424
rect 345952 449970 345980 451415
rect 347042 451344 347098 451353
rect 347042 451279 347098 451288
rect 347056 449970 347084 451279
rect 347792 449970 347820 451823
rect 348528 449970 348556 452134
rect 350632 452124 350684 452130
rect 350632 452066 350684 452072
rect 349252 451512 349304 451518
rect 349252 451454 349304 451460
rect 349114 450152 349166 450158
rect 349114 450094 349166 450100
rect 345216 449942 345460 449970
rect 345952 449942 346196 449970
rect 347056 449942 347300 449970
rect 347792 449942 348036 449970
rect 348160 449954 348404 449970
rect 348148 449948 348404 449954
rect 348200 449942 348404 449948
rect 348528 449942 348772 449970
rect 349126 449956 349154 450094
rect 349264 449970 349292 451454
rect 349264 449942 349508 449970
rect 348148 449890 348200 449896
rect 350644 449834 350672 452066
rect 350736 449970 350764 453999
rect 351460 451308 351512 451314
rect 351460 451250 351512 451256
rect 351472 449970 351500 451250
rect 351932 449970 351960 454922
rect 354680 454844 354732 454850
rect 354680 454786 354732 454792
rect 353300 454436 353352 454442
rect 353300 454378 353352 454384
rect 353024 452736 353076 452742
rect 353024 452678 353076 452684
rect 352194 451616 352250 451625
rect 352194 451551 352250 451560
rect 352656 451580 352708 451586
rect 352208 449970 352236 451551
rect 352656 451522 352708 451528
rect 352668 451382 352696 451522
rect 352564 451376 352616 451382
rect 352564 451318 352616 451324
rect 352656 451376 352708 451382
rect 352656 451318 352708 451324
rect 352576 449970 352604 451318
rect 352930 450256 352986 450265
rect 352930 450191 352986 450200
rect 352944 449993 352972 450191
rect 352930 449984 352986 449993
rect 350736 449942 350980 449970
rect 351472 449942 351716 449970
rect 351932 449942 352084 449970
rect 352208 449942 352452 449970
rect 352576 449942 352820 449970
rect 353036 449970 353064 452678
rect 353312 449970 353340 454378
rect 354128 452940 354180 452946
rect 354128 452882 354180 452888
rect 353668 451852 353720 451858
rect 353668 451794 353720 451800
rect 353680 449970 353708 451794
rect 354140 450158 354168 452882
rect 354588 451580 354640 451586
rect 354588 451522 354640 451528
rect 354600 450566 354628 451522
rect 354588 450560 354640 450566
rect 354588 450502 354640 450508
rect 354128 450152 354180 450158
rect 354128 450094 354180 450100
rect 353036 449942 353188 449970
rect 353312 449942 353556 449970
rect 353680 449942 353924 449970
rect 352930 449919 352986 449928
rect 350612 449806 350672 449834
rect 354140 449834 354168 450094
rect 354692 449970 354720 454786
rect 355048 454164 355100 454170
rect 355048 454106 355100 454112
rect 355060 451314 355088 454106
rect 355416 452600 355468 452606
rect 355416 452542 355468 452548
rect 355428 451926 355456 452542
rect 355416 451920 355468 451926
rect 355416 451862 355468 451868
rect 355048 451308 355100 451314
rect 355048 451250 355100 451256
rect 355060 449970 355088 451250
rect 355428 449970 355456 451862
rect 354660 449954 354904 449970
rect 354660 449948 354916 449954
rect 354660 449942 354864 449948
rect 355028 449942 355088 449970
rect 355396 449942 355456 449970
rect 355520 449970 355548 455874
rect 355980 452606 356008 456758
rect 356152 455864 356204 455870
rect 356152 455806 356204 455812
rect 355968 452600 356020 452606
rect 355968 452542 356020 452548
rect 355520 449942 355764 449970
rect 354864 449890 354916 449896
rect 356164 449834 356192 455806
rect 356244 453348 356296 453354
rect 356244 453290 356296 453296
rect 356256 452674 356284 453290
rect 356244 452668 356296 452674
rect 356244 452610 356296 452616
rect 356256 449970 356284 452610
rect 356716 451353 356744 472602
rect 357716 468512 357768 468518
rect 357716 468454 357768 468460
rect 356796 463004 356848 463010
rect 356796 462946 356848 462952
rect 356808 456794 356836 462946
rect 357348 460284 357400 460290
rect 357348 460226 357400 460232
rect 356808 456766 356928 456794
rect 356702 451344 356758 451353
rect 356702 451279 356758 451288
rect 356900 450294 356928 456766
rect 357360 455870 357388 460226
rect 357624 456136 357676 456142
rect 357624 456078 357676 456084
rect 357348 455864 357400 455870
rect 357348 455806 357400 455812
rect 357440 454844 357492 454850
rect 357440 454786 357492 454792
rect 357452 454238 357480 454786
rect 357636 454782 357664 456078
rect 357624 454776 357676 454782
rect 357624 454718 357676 454724
rect 357440 454232 357492 454238
rect 357440 454174 357492 454180
rect 357452 451466 357480 454174
rect 357452 451438 357572 451466
rect 356978 451344 357034 451353
rect 356978 451279 357034 451288
rect 357440 451308 357492 451314
rect 356888 450288 356940 450294
rect 356888 450230 356940 450236
rect 356256 449942 356500 449970
rect 356900 449834 356928 450230
rect 356992 449970 357020 451279
rect 357440 451250 357492 451256
rect 357452 450566 357480 451250
rect 357440 450560 357492 450566
rect 357440 450502 357492 450508
rect 357544 450242 357572 451438
rect 357728 450838 357756 468454
rect 357716 450832 357768 450838
rect 357716 450774 357768 450780
rect 357544 450214 357618 450242
rect 356992 449942 357236 449970
rect 357590 449956 357618 450214
rect 357728 449970 357756 450774
rect 357728 449942 357972 449970
rect 354140 449806 354292 449834
rect 356132 449806 356192 449834
rect 356868 449806 356928 449834
rect 346536 449576 346592 449585
rect 346536 449511 346592 449520
rect 342444 449472 342496 449478
rect 349620 449472 349672 449478
rect 342444 449414 342496 449420
rect 343822 449440 343878 449449
rect 342456 448594 342484 449414
rect 345800 449440 345856 449449
rect 343878 449398 343988 449426
rect 343822 449375 343878 449384
rect 351092 449472 351144 449478
rect 349986 449440 350042 449449
rect 349672 449420 349876 449426
rect 349620 449414 349876 449420
rect 349632 449398 349876 449414
rect 345800 449375 345856 449384
rect 350042 449398 350244 449426
rect 358096 449426 358124 576846
rect 359476 460934 359504 643078
rect 359556 630692 359608 630698
rect 359556 630634 359608 630640
rect 359108 460906 359504 460934
rect 358452 454776 358504 454782
rect 358452 454718 358504 454724
rect 358464 449970 358492 454718
rect 359108 453490 359136 460906
rect 359568 455802 359596 630634
rect 360120 456794 360148 670686
rect 361488 511284 361540 511290
rect 361488 511226 361540 511232
rect 360844 469872 360896 469878
rect 360844 469814 360896 469820
rect 360028 456766 360148 456794
rect 360856 456794 360884 469814
rect 361120 458856 361172 458862
rect 361120 458798 361172 458804
rect 360856 456766 361068 456794
rect 359556 455796 359608 455802
rect 359556 455738 359608 455744
rect 359096 453484 359148 453490
rect 359096 453426 359148 453432
rect 359108 449970 359136 453426
rect 359568 449970 359596 455738
rect 358464 449942 358708 449970
rect 359076 449942 359136 449970
rect 359444 449942 359596 449970
rect 359784 449440 359840 449449
rect 351144 449420 351348 449426
rect 351092 449414 351348 449420
rect 351104 449398 351348 449414
rect 358096 449410 358340 449426
rect 358084 449404 358340 449410
rect 349986 449375 350042 449384
rect 358136 449398 358340 449404
rect 360028 449426 360056 456766
rect 360934 451480 360990 451489
rect 360934 451415 360990 451424
rect 360750 451344 360806 451353
rect 360750 451279 360806 451288
rect 360200 450764 360252 450770
rect 360200 450706 360252 450712
rect 360212 449970 360240 450706
rect 360180 449942 360240 449970
rect 360382 449984 360438 449993
rect 360764 449970 360792 451279
rect 360948 449970 360976 451415
rect 361040 450362 361068 456766
rect 361132 451489 361160 458798
rect 361396 453484 361448 453490
rect 361396 453426 361448 453432
rect 361118 451480 361174 451489
rect 361118 451415 361174 451424
rect 361408 450770 361436 453426
rect 361500 451353 361528 511226
rect 362224 465724 362276 465730
rect 362224 465666 362276 465672
rect 361672 456000 361724 456006
rect 361672 455942 361724 455948
rect 361684 455734 361712 455942
rect 361672 455728 361724 455734
rect 361672 455670 361724 455676
rect 361486 451344 361542 451353
rect 361486 451279 361542 451288
rect 361396 450764 361448 450770
rect 361396 450706 361448 450712
rect 361028 450356 361080 450362
rect 361028 450298 361080 450304
rect 360438 449942 360792 449970
rect 360916 449956 360976 449970
rect 360902 449942 360976 449956
rect 361040 449970 361068 450298
rect 361684 449970 361712 455670
rect 362236 455530 362264 465666
rect 362316 464364 362368 464370
rect 362316 464306 362368 464312
rect 362328 456006 362356 464306
rect 363144 460216 363196 460222
rect 363144 460158 363196 460164
rect 362868 456068 362920 456074
rect 362868 456010 362920 456016
rect 362316 456000 362368 456006
rect 362316 455942 362368 455948
rect 362224 455524 362276 455530
rect 362224 455466 362276 455472
rect 362040 454708 362092 454714
rect 362040 454650 362092 454656
rect 362052 449970 362080 454650
rect 362236 453914 362264 455466
rect 362236 453886 362540 453914
rect 362408 453280 362460 453286
rect 362408 453222 362460 453228
rect 362420 449970 362448 453222
rect 361040 449942 361284 449970
rect 361652 449942 361712 449970
rect 362020 449942 362080 449970
rect 362388 449942 362448 449970
rect 362512 449970 362540 453886
rect 362880 453286 362908 456010
rect 363156 454646 363184 460158
rect 363144 454640 363196 454646
rect 363144 454582 363196 454588
rect 362868 453280 362920 453286
rect 362868 453222 362920 453228
rect 363156 449970 363184 454582
rect 363328 451920 363380 451926
rect 363328 451862 363380 451868
rect 362512 449942 362756 449970
rect 363124 449942 363184 449970
rect 360382 449919 360438 449928
rect 360658 449848 360714 449857
rect 360902 449834 360930 449942
rect 360714 449820 360930 449834
rect 360714 449806 360916 449820
rect 360658 449783 360714 449792
rect 363340 449614 363368 451862
rect 363616 451858 363644 698634
rect 363972 474020 364024 474026
rect 363972 473962 364024 473968
rect 363604 451852 363656 451858
rect 363604 451794 363656 451800
rect 363510 451344 363566 451353
rect 363510 451279 363566 451288
rect 363524 449970 363552 451279
rect 363492 449942 363552 449970
rect 363602 449984 363658 449993
rect 363984 449970 364012 473962
rect 364156 461712 364208 461718
rect 364156 461654 364208 461660
rect 364064 451852 364116 451858
rect 364064 451794 364116 451800
rect 363658 449942 364012 449970
rect 364076 449970 364104 451794
rect 364168 451353 364196 461654
rect 364444 455666 364472 700266
rect 364536 456794 364564 700334
rect 364996 698698 365024 703520
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 364984 698692 365036 698698
rect 364984 698634 365036 698640
rect 378784 696992 378836 696998
rect 378784 696934 378836 696940
rect 369860 683188 369912 683194
rect 369860 683130 369912 683136
rect 367744 590708 367796 590714
rect 367744 590650 367796 590656
rect 367756 468518 367784 590650
rect 367836 470620 367888 470626
rect 367836 470562 367888 470568
rect 367744 468512 367796 468518
rect 367744 468454 367796 468460
rect 367284 463752 367336 463758
rect 367284 463694 367336 463700
rect 365720 461644 365772 461650
rect 365720 461586 365772 461592
rect 364536 456766 364748 456794
rect 364432 455660 364484 455666
rect 364432 455602 364484 455608
rect 364154 451344 364210 451353
rect 364154 451279 364210 451288
rect 364444 449970 364472 455602
rect 364720 451382 364748 456766
rect 365076 453416 365128 453422
rect 365076 453358 365128 453364
rect 364708 451376 364760 451382
rect 364708 451318 364760 451324
rect 364720 449970 364748 451318
rect 365088 449993 365116 453358
rect 365732 451926 365760 461586
rect 367100 453212 367152 453218
rect 367100 453154 367152 453160
rect 365720 451920 365772 451926
rect 365720 451862 365772 451868
rect 366180 451920 366232 451926
rect 366180 451862 366232 451868
rect 365812 451784 365864 451790
rect 365812 451726 365864 451732
rect 365720 451308 365772 451314
rect 365720 451250 365772 451256
rect 365732 450537 365760 451250
rect 365718 450528 365774 450537
rect 365718 450463 365774 450472
rect 365444 450084 365496 450090
rect 365444 450026 365496 450032
rect 365074 449984 365130 449993
rect 364076 449942 364228 449970
rect 364444 449942 364596 449970
rect 364720 449942 364964 449970
rect 363602 449919 363658 449928
rect 363328 449608 363380 449614
rect 363328 449550 363380 449556
rect 364076 449426 364104 449942
rect 365456 449970 365484 450026
rect 365824 449970 365852 451726
rect 366192 449970 366220 451862
rect 366548 451512 366600 451518
rect 366548 451454 366600 451460
rect 366560 449970 366588 451454
rect 367112 451382 367140 453154
rect 367192 451988 367244 451994
rect 367192 451930 367244 451936
rect 367100 451376 367152 451382
rect 367100 451318 367152 451324
rect 367204 449970 367232 451930
rect 365130 449942 365332 449970
rect 365456 449942 365700 449970
rect 365824 449942 366068 449970
rect 366192 449942 366436 449970
rect 366560 449942 366804 449970
rect 367172 449942 367232 449970
rect 367296 449970 367324 463694
rect 367848 460290 367876 470562
rect 368572 467152 368624 467158
rect 368572 467094 368624 467100
rect 368480 465112 368532 465118
rect 368480 465054 368532 465060
rect 367836 460284 367888 460290
rect 367836 460226 367888 460232
rect 368018 454200 368074 454209
rect 368018 454135 368074 454144
rect 367882 450220 367934 450226
rect 367882 450162 367934 450168
rect 367296 449942 367540 449970
rect 367894 449956 367922 450162
rect 368032 449970 368060 454135
rect 368492 449970 368520 465054
rect 368584 451353 368612 467094
rect 369122 452704 369178 452713
rect 369122 452639 369178 452648
rect 368570 451344 368626 451353
rect 368570 451279 368626 451288
rect 368984 450256 369040 450265
rect 368984 450191 369040 450200
rect 368032 449942 368276 449970
rect 368492 449942 368644 449970
rect 368998 449956 369026 450191
rect 369136 449970 369164 452639
rect 369490 451344 369546 451353
rect 369490 451279 369546 451288
rect 369504 449970 369532 451279
rect 369136 449942 369380 449970
rect 369504 449942 369748 449970
rect 365074 449919 365130 449928
rect 365088 449859 365116 449919
rect 369872 449478 369900 683130
rect 371240 632120 371292 632126
rect 371240 632062 371292 632068
rect 369952 451308 370004 451314
rect 369952 451250 370004 451256
rect 369964 449970 369992 451250
rect 371252 450226 371280 632062
rect 372620 579692 372672 579698
rect 372620 579634 372672 579640
rect 372632 460934 372660 579634
rect 376024 563100 376076 563106
rect 376024 563042 376076 563048
rect 374000 527196 374052 527202
rect 374000 527138 374052 527144
rect 372632 460906 372844 460934
rect 372712 456952 372764 456958
rect 372712 456894 372764 456900
rect 371424 456884 371476 456890
rect 371424 456826 371476 456832
rect 371332 453144 371384 453150
rect 371332 453086 371384 453092
rect 371344 451994 371372 453086
rect 371332 451988 371384 451994
rect 371332 451930 371384 451936
rect 371436 451274 371464 456826
rect 371344 451246 371464 451274
rect 371240 450220 371292 450226
rect 371240 450162 371292 450168
rect 370456 450120 370512 450129
rect 370456 450055 370512 450064
rect 369964 449942 370116 449970
rect 370470 449956 370498 450055
rect 371344 449970 371372 451246
rect 371700 450220 371752 450226
rect 371700 450162 371752 450168
rect 371344 449942 371588 449970
rect 371712 449834 371740 450162
rect 372068 450016 372120 450022
rect 372724 449970 372752 456894
rect 372120 449964 372324 449970
rect 372068 449958 372324 449964
rect 372080 449942 372324 449958
rect 372692 449942 372752 449970
rect 371712 449806 372016 449834
rect 370608 449478 370636 449509
rect 359840 449398 360056 449426
rect 363984 449410 364104 449426
rect 369860 449472 369912 449478
rect 370596 449472 370648 449478
rect 369860 449414 369912 449420
rect 370594 449440 370596 449449
rect 370648 449440 370650 449449
rect 363972 449404 364104 449410
rect 359784 449375 359840 449384
rect 358084 449346 358136 449352
rect 364024 449398 364104 449404
rect 370650 449398 370852 449426
rect 371988 449392 372016 449806
rect 372816 449426 372844 460906
rect 373540 457292 373592 457298
rect 373540 457234 373592 457240
rect 373172 450424 373224 450430
rect 373172 450366 373224 450372
rect 373184 449970 373212 450366
rect 373552 449970 373580 457234
rect 373184 449942 373428 449970
rect 373552 449942 373796 449970
rect 373170 449440 373226 449449
rect 372816 449398 373170 449426
rect 370594 449375 370650 449384
rect 363972 449346 364024 449352
rect 371942 449364 372016 449392
rect 374012 449426 374040 527138
rect 374460 474768 374512 474774
rect 374460 474710 374512 474716
rect 374276 454096 374328 454102
rect 374276 454038 374328 454044
rect 374288 449970 374316 454038
rect 374472 452577 374500 474710
rect 375748 457088 375800 457094
rect 375748 457030 375800 457036
rect 374458 452568 374514 452577
rect 374458 452503 374514 452512
rect 374644 451716 374696 451722
rect 374644 451658 374696 451664
rect 374656 449970 374684 451658
rect 375380 451376 375432 451382
rect 375380 451318 375432 451324
rect 375392 449970 375420 451318
rect 375760 449970 375788 457030
rect 376036 454850 376064 563042
rect 377404 536852 377456 536858
rect 377404 536794 377456 536800
rect 377416 463010 377444 536794
rect 377404 463004 377456 463010
rect 377404 462946 377456 462952
rect 376024 454844 376076 454850
rect 376024 454786 376076 454792
rect 376760 454572 376812 454578
rect 376760 454514 376812 454520
rect 376116 453008 376168 453014
rect 376116 452950 376168 452956
rect 376128 449970 376156 452950
rect 376772 452606 376800 454514
rect 378692 454504 378744 454510
rect 378692 454446 378744 454452
rect 378324 454368 378376 454374
rect 378324 454310 378376 454316
rect 376944 454300 376996 454306
rect 376944 454242 376996 454248
rect 376760 452600 376812 452606
rect 376760 452542 376812 452548
rect 376760 451988 376812 451994
rect 376760 451930 376812 451936
rect 376772 449970 376800 451930
rect 374288 449942 374532 449970
rect 374656 449942 374900 449970
rect 375392 449942 375636 449970
rect 375760 449942 376004 449970
rect 376128 449942 376372 449970
rect 376740 449942 376800 449970
rect 376956 449970 376984 454242
rect 377220 453076 377272 453082
rect 377220 453018 377272 453024
rect 377232 449970 377260 453018
rect 377586 451344 377642 451353
rect 377586 451279 377642 451288
rect 377600 449970 377628 451279
rect 378336 449970 378364 454310
rect 378416 453552 378468 453558
rect 378416 453494 378468 453500
rect 376956 449942 377108 449970
rect 377232 449942 377476 449970
rect 377600 449942 377844 449970
rect 378212 449942 378364 449970
rect 378428 449970 378456 453494
rect 378704 449970 378732 454446
rect 378796 453490 378824 696934
rect 382924 616888 382976 616894
rect 382924 616830 382976 616836
rect 381084 457156 381136 457162
rect 381084 457098 381136 457104
rect 380164 455592 380216 455598
rect 380164 455534 380216 455540
rect 379796 454912 379848 454918
rect 379796 454854 379848 454860
rect 378784 453484 378836 453490
rect 378784 453426 378836 453432
rect 379060 452600 379112 452606
rect 379060 452542 379112 452548
rect 379072 449970 379100 452542
rect 379428 450628 379480 450634
rect 379428 450570 379480 450576
rect 379440 449970 379468 450570
rect 379808 449970 379836 454854
rect 380176 449970 380204 455534
rect 380532 450696 380584 450702
rect 380532 450638 380584 450644
rect 380544 449970 380572 450638
rect 381096 450242 381124 457098
rect 381268 457020 381320 457026
rect 381268 456962 381320 456968
rect 381096 450214 381170 450242
rect 378428 449942 378580 449970
rect 378704 449942 378948 449970
rect 379072 449942 379316 449970
rect 379440 449942 379684 449970
rect 379808 449942 380052 449970
rect 380176 449942 380420 449970
rect 380544 449942 380788 449970
rect 381142 449956 381170 450214
rect 381280 449970 381308 456962
rect 382936 456142 382964 616830
rect 392584 524476 392636 524482
rect 392584 524418 392636 524424
rect 392596 472666 392624 524418
rect 392584 472660 392636 472666
rect 392584 472602 392636 472608
rect 396736 461718 396764 699654
rect 412652 474026 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 412640 474020 412692 474026
rect 412640 473962 412692 473968
rect 396724 461712 396776 461718
rect 396724 461654 396776 461660
rect 429212 460222 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 460216 429252 460222
rect 429200 460158 429252 460164
rect 384212 457224 384264 457230
rect 384212 457166 384264 457172
rect 382924 456136 382976 456142
rect 382924 456078 382976 456084
rect 383108 455456 383160 455462
rect 383108 455398 383160 455404
rect 381636 452872 381688 452878
rect 381636 452814 381688 452820
rect 381648 449970 381676 452814
rect 382372 451444 382424 451450
rect 382372 451386 382424 451392
rect 382384 449970 382412 451386
rect 382740 450492 382792 450498
rect 382740 450434 382792 450440
rect 382752 449970 382780 450434
rect 383120 449970 383148 455398
rect 383844 453620 383896 453626
rect 383844 453562 383896 453568
rect 383856 449970 383884 453562
rect 384224 449970 384252 457166
rect 462332 456074 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 465730 477540 702406
rect 477500 465724 477552 465730
rect 477500 465666 477552 465672
rect 462320 456068 462372 456074
rect 462320 456010 462372 456016
rect 494072 454714 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 469878 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 527180 469872 527232 469878
rect 527180 469814 527232 469820
rect 542372 464370 542400 702406
rect 542360 464364 542412 464370
rect 542360 464306 542412 464312
rect 558932 458862 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580276 511290 580304 683839
rect 580354 511320 580410 511329
rect 580264 511284 580316 511290
rect 580354 511255 580410 511264
rect 580264 511226 580316 511232
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580078 471472 580134 471481
rect 580078 471407 580134 471416
rect 580092 470626 580120 471407
rect 580080 470620 580132 470626
rect 580080 470562 580132 470568
rect 558920 458856 558972 458862
rect 558920 458798 558972 458804
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 494060 454708 494112 454714
rect 494060 454650 494112 454656
rect 580368 453354 580396 511255
rect 580356 453348 580408 453354
rect 580356 453290 580408 453296
rect 385040 452804 385092 452810
rect 385040 452746 385092 452752
rect 384580 451580 384632 451586
rect 384580 451522 384632 451528
rect 384592 449970 384620 451522
rect 385052 449970 385080 452746
rect 385684 452056 385736 452062
rect 385684 451998 385736 452004
rect 385696 449970 385724 451998
rect 580264 450560 580316 450566
rect 580264 450502 580316 450508
rect 388444 450152 388496 450158
rect 388444 450094 388496 450100
rect 381280 449942 381524 449970
rect 381648 449942 381892 449970
rect 382384 449942 382628 449970
rect 382752 449942 382996 449970
rect 383120 449942 383364 449970
rect 383856 449942 384100 449970
rect 384224 449942 384468 449970
rect 384592 449942 384836 449970
rect 385052 449942 385204 449970
rect 385696 449942 385940 449970
rect 375010 449576 375066 449585
rect 375066 449534 375268 449562
rect 375010 449511 375066 449520
rect 374274 449440 374330 449449
rect 374012 449398 374274 449426
rect 373170 449375 373226 449384
rect 374274 449375 374330 449384
rect 385314 449440 385370 449449
rect 385370 449398 385572 449426
rect 385314 449375 385370 449384
rect 371942 449313 371970 449364
rect 346904 449304 346960 449313
rect 346904 449239 346960 449248
rect 347640 449304 347696 449313
rect 347640 449239 347696 449248
rect 359784 449304 359840 449313
rect 359784 449239 359840 449248
rect 371192 449304 371248 449313
rect 371192 449239 371248 449248
rect 371928 449304 371984 449313
rect 371928 449239 371984 449248
rect 382232 449304 382288 449313
rect 382232 449239 382288 449248
rect 383704 449304 383760 449313
rect 383704 449239 383760 449248
rect 342444 448588 342496 448594
rect 342444 448530 342496 448536
rect 342364 447106 342484 447134
rect 342456 439521 342484 447106
rect 342442 439512 342498 439521
rect 342442 439447 342498 439456
rect 388456 422294 388484 450094
rect 389824 449948 389876 449954
rect 389824 449890 389876 449896
rect 389836 431934 389864 449890
rect 389824 431928 389876 431934
rect 389824 431870 389876 431876
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 388456 422266 389036 422294
rect 389008 405686 389036 422266
rect 580276 418305 580304 450502
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 388996 405680 389048 405686
rect 388996 405622 389048 405628
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 342258 401976 342314 401985
rect 342258 401911 342314 401920
rect 342272 400858 342300 401911
rect 342260 400852 342312 400858
rect 342260 400794 342312 400800
rect 342258 400616 342314 400625
rect 342258 400551 342314 400560
rect 342272 400518 342300 400551
rect 342260 400512 342312 400518
rect 342260 400454 342312 400460
rect 387800 400512 387852 400518
rect 387800 400454 387852 400460
rect 392124 400512 392176 400518
rect 392124 400454 392176 400460
rect 342260 400376 342312 400382
rect 387812 400353 387840 400454
rect 390192 400376 390244 400382
rect 387798 400344 387854 400353
rect 342260 400318 342312 400324
rect 342272 399566 342300 400318
rect 387412 400302 387748 400330
rect 342352 399900 342404 399906
rect 342352 399842 342404 399848
rect 342260 399560 342312 399566
rect 342260 399502 342312 399508
rect 342364 398834 342392 399842
rect 342502 399786 342530 400044
rect 342594 399906 342622 400044
rect 342582 399900 342634 399906
rect 342582 399842 342634 399848
rect 342502 399758 342576 399786
rect 342272 398806 342392 398834
rect 342272 391406 342300 398806
rect 342444 397996 342496 398002
rect 342444 397938 342496 397944
rect 342456 394126 342484 397938
rect 342548 397746 342576 399758
rect 342686 399684 342714 400044
rect 342778 399906 342806 400044
rect 342766 399900 342818 399906
rect 342766 399842 342818 399848
rect 342870 399684 342898 400044
rect 342962 399809 342990 400044
rect 343054 399945 343082 400044
rect 343040 399936 343096 399945
rect 343040 399871 343096 399880
rect 342948 399800 343004 399809
rect 343146 399752 343174 400044
rect 343238 399809 343266 400044
rect 342948 399735 343004 399744
rect 343100 399724 343174 399752
rect 343224 399800 343280 399809
rect 343224 399735 343280 399744
rect 342686 399656 342760 399684
rect 342870 399656 342944 399684
rect 342548 397718 342668 397746
rect 342444 394120 342496 394126
rect 342444 394062 342496 394068
rect 342536 393916 342588 393922
rect 342536 393858 342588 393864
rect 342444 393848 342496 393854
rect 342444 393790 342496 393796
rect 342260 391400 342312 391406
rect 342260 391342 342312 391348
rect 342456 389910 342484 393790
rect 342444 389904 342496 389910
rect 342444 389846 342496 389852
rect 342168 365696 342220 365702
rect 342168 365638 342220 365644
rect 341982 329352 342038 329361
rect 341982 329287 342038 329296
rect 341996 317286 342024 329287
rect 342260 323672 342312 323678
rect 342260 323614 342312 323620
rect 342272 320385 342300 323614
rect 342258 320376 342314 320385
rect 342258 320311 342314 320320
rect 341984 317280 342036 317286
rect 341984 317222 342036 317228
rect 341892 314220 341944 314226
rect 341892 314162 341944 314168
rect 341800 312996 341852 313002
rect 341800 312938 341852 312944
rect 341708 310412 341760 310418
rect 341708 310354 341760 310360
rect 341616 304224 341668 304230
rect 341616 304166 341668 304172
rect 341524 295316 341576 295322
rect 341524 295258 341576 295264
rect 342272 226234 342300 320311
rect 342548 319297 342576 393858
rect 342640 389978 342668 397718
rect 342732 392970 342760 399656
rect 342812 399560 342864 399566
rect 342812 399502 342864 399508
rect 342720 392964 342772 392970
rect 342720 392906 342772 392912
rect 342628 389972 342680 389978
rect 342628 389914 342680 389920
rect 342824 387190 342852 399502
rect 342916 398546 342944 399656
rect 342904 398540 342956 398546
rect 342904 398482 342956 398488
rect 342904 398268 342956 398274
rect 342904 398210 342956 398216
rect 342812 387184 342864 387190
rect 342812 387126 342864 387132
rect 342534 319288 342590 319297
rect 342534 319223 342590 319232
rect 342916 311302 342944 398210
rect 343100 397866 343128 399724
rect 343330 399684 343358 400044
rect 343284 399656 343358 399684
rect 343178 398712 343234 398721
rect 343178 398647 343234 398656
rect 343088 397860 343140 397866
rect 343088 397802 343140 397808
rect 342996 394052 343048 394058
rect 342996 393994 343048 394000
rect 342904 311296 342956 311302
rect 342904 311238 342956 311244
rect 342352 311024 342404 311030
rect 342352 310966 342404 310972
rect 342364 309942 342392 310966
rect 342352 309936 342404 309942
rect 342352 309878 342404 309884
rect 342904 309936 342956 309942
rect 342904 309878 342956 309884
rect 342260 226228 342312 226234
rect 342260 226170 342312 226176
rect 340972 222148 341024 222154
rect 340972 222090 341024 222096
rect 340878 220824 340934 220833
rect 340878 220759 340934 220768
rect 342260 200116 342312 200122
rect 342260 200058 342312 200064
rect 342272 199510 342300 200058
rect 342916 199510 342944 309878
rect 343008 296614 343036 393994
rect 343088 389972 343140 389978
rect 343088 389914 343140 389920
rect 343100 305658 343128 389914
rect 343192 388618 343220 398647
rect 343284 393922 343312 399656
rect 343422 399616 343450 400044
rect 343514 399684 343542 400044
rect 343606 399786 343634 400044
rect 343698 399906 343726 400044
rect 343790 399945 343818 400044
rect 343776 399936 343832 399945
rect 343686 399900 343738 399906
rect 343776 399871 343832 399880
rect 343686 399842 343738 399848
rect 343606 399758 343680 399786
rect 343514 399656 343588 399684
rect 343376 399588 343450 399616
rect 343376 398002 343404 399588
rect 343364 397996 343416 398002
rect 343364 397938 343416 397944
rect 343560 395214 343588 399656
rect 343652 396642 343680 399758
rect 343882 399752 343910 400044
rect 343974 399786 344002 400044
rect 344066 399906 344094 400044
rect 344158 399906 344186 400044
rect 344054 399900 344106 399906
rect 344054 399842 344106 399848
rect 344146 399900 344198 399906
rect 344146 399842 344198 399848
rect 344098 399800 344154 399809
rect 343974 399758 344048 399786
rect 343836 399724 343910 399752
rect 343836 399566 343864 399724
rect 344020 399650 344048 399758
rect 344098 399735 344154 399744
rect 344250 399752 344278 400044
rect 344342 399945 344370 400044
rect 344328 399936 344384 399945
rect 344328 399871 344384 399880
rect 344434 399838 344462 400044
rect 344526 399906 344554 400044
rect 344618 399906 344646 400044
rect 344710 399945 344738 400044
rect 344696 399936 344752 399945
rect 344514 399900 344566 399906
rect 344514 399842 344566 399848
rect 344606 399900 344658 399906
rect 344802 399906 344830 400044
rect 344696 399871 344752 399880
rect 344790 399900 344842 399906
rect 344606 399842 344658 399848
rect 344790 399842 344842 399848
rect 344422 399832 344474 399838
rect 344422 399774 344474 399780
rect 344744 399764 344796 399770
rect 343928 399622 344048 399650
rect 343824 399560 343876 399566
rect 343824 399502 343876 399508
rect 343824 398744 343876 398750
rect 343824 398686 343876 398692
rect 343640 396636 343692 396642
rect 343640 396578 343692 396584
rect 343640 395276 343692 395282
rect 343640 395218 343692 395224
rect 343548 395208 343600 395214
rect 343548 395150 343600 395156
rect 343272 393916 343324 393922
rect 343272 393858 343324 393864
rect 343546 393544 343602 393553
rect 343546 393479 343602 393488
rect 343456 392964 343508 392970
rect 343456 392906 343508 392912
rect 343364 391332 343416 391338
rect 343364 391274 343416 391280
rect 343180 388612 343232 388618
rect 343180 388554 343232 388560
rect 343180 384668 343232 384674
rect 343180 384610 343232 384616
rect 343088 305652 343140 305658
rect 343088 305594 343140 305600
rect 343192 302802 343220 384610
rect 343272 381676 343324 381682
rect 343272 381618 343324 381624
rect 343180 302796 343232 302802
rect 343180 302738 343232 302744
rect 343284 302734 343312 381618
rect 343376 312798 343404 391274
rect 343468 321065 343496 392906
rect 343560 392562 343588 393479
rect 343548 392556 343600 392562
rect 343548 392498 343600 392504
rect 343548 388680 343600 388686
rect 343548 388622 343600 388628
rect 343454 321056 343510 321065
rect 343454 320991 343510 321000
rect 343364 312792 343416 312798
rect 343364 312734 343416 312740
rect 343560 312497 343588 388622
rect 343652 319462 343680 395218
rect 343836 381721 343864 398686
rect 343928 398478 343956 399622
rect 344008 399560 344060 399566
rect 344008 399502 344060 399508
rect 343916 398472 343968 398478
rect 343916 398414 343968 398420
rect 343822 381712 343878 381721
rect 343822 381647 343878 381656
rect 344020 319705 344048 399502
rect 344112 398410 344140 399735
rect 344250 399724 344324 399752
rect 344192 399628 344244 399634
rect 344192 399570 344244 399576
rect 344100 398404 344152 398410
rect 344100 398346 344152 398352
rect 344098 393408 344154 393417
rect 344098 393343 344154 393352
rect 344006 319696 344062 319705
rect 344006 319631 344062 319640
rect 343640 319456 343692 319462
rect 343640 319398 343692 319404
rect 344112 319190 344140 393343
rect 344204 387297 344232 399570
rect 344296 393530 344324 399724
rect 344744 399706 344796 399712
rect 344376 399696 344428 399702
rect 344376 399638 344428 399644
rect 344652 399696 344704 399702
rect 344652 399638 344704 399644
rect 344388 393854 344416 399638
rect 344560 399492 344612 399498
rect 344560 399434 344612 399440
rect 344376 393848 344428 393854
rect 344376 393790 344428 393796
rect 344296 393502 344416 393530
rect 344388 393310 344416 393502
rect 344376 393304 344428 393310
rect 344376 393246 344428 393252
rect 344284 392420 344336 392426
rect 344284 392362 344336 392368
rect 344190 387288 344246 387297
rect 344190 387223 344246 387232
rect 344100 319184 344152 319190
rect 344100 319126 344152 319132
rect 343546 312488 343602 312497
rect 343546 312423 343602 312432
rect 344296 305930 344324 392362
rect 344572 389881 344600 399434
rect 344664 398585 344692 399638
rect 344756 398721 344784 399706
rect 344894 399684 344922 400044
rect 344848 399656 344922 399684
rect 344848 398750 344876 399656
rect 344986 399616 345014 400044
rect 345078 399945 345106 400044
rect 345064 399936 345120 399945
rect 345064 399871 345120 399880
rect 345170 399752 345198 400044
rect 344940 399588 345014 399616
rect 345124 399724 345198 399752
rect 344836 398744 344888 398750
rect 344742 398712 344798 398721
rect 344836 398686 344888 398692
rect 344742 398647 344798 398656
rect 344650 398576 344706 398585
rect 344940 398528 344968 399588
rect 344650 398511 344706 398520
rect 344756 398500 344968 398528
rect 345020 398540 345072 398546
rect 344650 398168 344706 398177
rect 344650 398103 344706 398112
rect 344664 391406 344692 398103
rect 344652 391400 344704 391406
rect 344756 391377 344784 398500
rect 345020 398482 345072 398488
rect 344928 398404 344980 398410
rect 344928 398346 344980 398352
rect 344836 397928 344888 397934
rect 344836 397870 344888 397876
rect 344652 391342 344704 391348
rect 344742 391368 344798 391377
rect 344742 391303 344798 391312
rect 344558 389872 344614 389881
rect 344558 389807 344614 389816
rect 344560 387184 344612 387190
rect 344560 387126 344612 387132
rect 344468 385008 344520 385014
rect 344468 384950 344520 384956
rect 344374 381984 344430 381993
rect 344374 381919 344430 381928
rect 344284 305924 344336 305930
rect 344284 305866 344336 305872
rect 343272 302728 343324 302734
rect 343272 302670 343324 302676
rect 343638 301744 343694 301753
rect 343638 301679 343694 301688
rect 342996 296608 343048 296614
rect 342996 296550 343048 296556
rect 343652 232665 343680 301679
rect 344388 301442 344416 381919
rect 344480 304434 344508 384950
rect 344572 307358 344600 387126
rect 344848 386414 344876 397870
rect 344756 386386 344876 386414
rect 344756 321162 344784 386386
rect 344836 384736 344888 384742
rect 344836 384678 344888 384684
rect 344744 321156 344796 321162
rect 344744 321098 344796 321104
rect 344848 309874 344876 384678
rect 344940 378593 344968 398346
rect 345032 395146 345060 398482
rect 345124 398342 345152 399724
rect 345262 399684 345290 400044
rect 345354 399906 345382 400044
rect 345342 399900 345394 399906
rect 345342 399842 345394 399848
rect 345446 399786 345474 400044
rect 345216 399656 345290 399684
rect 345400 399758 345474 399786
rect 345112 398336 345164 398342
rect 345112 398278 345164 398284
rect 345020 395140 345072 395146
rect 345020 395082 345072 395088
rect 345020 395004 345072 395010
rect 345020 394946 345072 394952
rect 345032 389065 345060 394946
rect 345216 392902 345244 399656
rect 345296 399560 345348 399566
rect 345296 399502 345348 399508
rect 345308 393666 345336 399502
rect 345400 398041 345428 399758
rect 345538 399684 345566 400044
rect 345630 399945 345658 400044
rect 345616 399936 345672 399945
rect 345616 399871 345672 399880
rect 345722 399820 345750 400044
rect 345492 399656 345566 399684
rect 345676 399792 345750 399820
rect 345386 398032 345442 398041
rect 345386 397967 345442 397976
rect 345308 393638 345428 393666
rect 345296 393508 345348 393514
rect 345296 393450 345348 393456
rect 345204 392896 345256 392902
rect 345204 392838 345256 392844
rect 345018 389056 345074 389065
rect 345018 388991 345074 389000
rect 345308 378894 345336 393450
rect 345296 378888 345348 378894
rect 345296 378830 345348 378836
rect 344926 378584 344982 378593
rect 344926 378519 344982 378528
rect 345400 356726 345428 393638
rect 345492 392970 345520 399656
rect 345572 399560 345624 399566
rect 345572 399502 345624 399508
rect 345480 392964 345532 392970
rect 345480 392906 345532 392912
rect 345584 390250 345612 399502
rect 345676 398857 345704 399792
rect 345814 399752 345842 400044
rect 345906 399809 345934 400044
rect 345998 399838 346026 400044
rect 346090 399945 346118 400044
rect 346076 399936 346132 399945
rect 346182 399906 346210 400044
rect 346076 399871 346132 399880
rect 346170 399900 346222 399906
rect 346170 399842 346222 399848
rect 345986 399832 346038 399838
rect 345768 399724 345842 399752
rect 345892 399800 345948 399809
rect 345986 399774 346038 399780
rect 346274 399752 346302 400044
rect 346366 399906 346394 400044
rect 346458 399945 346486 400044
rect 346444 399936 346500 399945
rect 346354 399900 346406 399906
rect 346444 399871 346500 399880
rect 346354 399842 346406 399848
rect 346550 399820 346578 400044
rect 345892 399735 345948 399744
rect 346228 399724 346302 399752
rect 346504 399792 346578 399820
rect 345662 398848 345718 398857
rect 345662 398783 345718 398792
rect 345664 398472 345716 398478
rect 345664 398414 345716 398420
rect 345676 397730 345704 398414
rect 345664 397724 345716 397730
rect 345664 397666 345716 397672
rect 345664 397384 345716 397390
rect 345664 397326 345716 397332
rect 345676 396778 345704 397326
rect 345664 396772 345716 396778
rect 345664 396714 345716 396720
rect 345768 394330 345796 399724
rect 345940 399628 345992 399634
rect 345940 399570 345992 399576
rect 345952 398546 345980 399570
rect 346032 398744 346084 398750
rect 346032 398686 346084 398692
rect 345940 398540 345992 398546
rect 345940 398482 345992 398488
rect 346044 398002 346072 398686
rect 346124 398540 346176 398546
rect 346124 398482 346176 398488
rect 346136 398342 346164 398482
rect 346124 398336 346176 398342
rect 346124 398278 346176 398284
rect 346032 397996 346084 398002
rect 346032 397938 346084 397944
rect 345848 397724 345900 397730
rect 345848 397666 345900 397672
rect 345756 394324 345808 394330
rect 345756 394266 345808 394272
rect 345664 393576 345716 393582
rect 345664 393518 345716 393524
rect 345572 390244 345624 390250
rect 345572 390186 345624 390192
rect 345570 388376 345626 388385
rect 345570 388311 345626 388320
rect 345584 371958 345612 388311
rect 345572 371952 345624 371958
rect 345572 371894 345624 371900
rect 345388 356720 345440 356726
rect 345388 356662 345440 356668
rect 345018 325816 345074 325825
rect 345018 325751 345074 325760
rect 344926 325408 344982 325417
rect 344926 325343 344982 325352
rect 344836 309868 344888 309874
rect 344836 309810 344888 309816
rect 344560 307352 344612 307358
rect 344560 307294 344612 307300
rect 344468 304428 344520 304434
rect 344468 304370 344520 304376
rect 344940 301753 344968 325343
rect 344926 301744 344982 301753
rect 344926 301679 344982 301688
rect 344376 301436 344428 301442
rect 344376 301378 344428 301384
rect 343638 232656 343694 232665
rect 343638 232591 343694 232600
rect 345032 226302 345060 325751
rect 345676 301578 345704 393518
rect 345860 390017 345888 397666
rect 346032 396704 346084 396710
rect 346032 396646 346084 396652
rect 345940 390516 345992 390522
rect 345940 390458 345992 390464
rect 345846 390008 345902 390017
rect 345846 389943 345902 389952
rect 345952 389881 345980 390458
rect 345938 389872 345994 389881
rect 345938 389807 345994 389816
rect 345940 384940 345992 384946
rect 345940 384882 345992 384888
rect 345848 384600 345900 384606
rect 345848 384542 345900 384548
rect 345756 381608 345808 381614
rect 345756 381550 345808 381556
rect 345664 301572 345716 301578
rect 345664 301514 345716 301520
rect 345768 297634 345796 381550
rect 345860 300150 345888 384542
rect 345952 304502 345980 384882
rect 346044 317966 346072 396646
rect 346124 392964 346176 392970
rect 346124 392906 346176 392912
rect 346136 321201 346164 392906
rect 346228 388249 346256 399724
rect 346504 399650 346532 399792
rect 346642 399752 346670 400044
rect 346734 399906 346762 400044
rect 346722 399900 346774 399906
rect 346722 399842 346774 399848
rect 346826 399786 346854 400044
rect 346412 399622 346532 399650
rect 346596 399724 346670 399752
rect 346780 399758 346854 399786
rect 346308 399492 346360 399498
rect 346308 399434 346360 399440
rect 346320 391241 346348 399434
rect 346306 391232 346362 391241
rect 346306 391167 346362 391176
rect 346214 388240 346270 388249
rect 346214 388175 346270 388184
rect 346412 387569 346440 399622
rect 346492 396092 346544 396098
rect 346492 396034 346544 396040
rect 346398 387560 346454 387569
rect 346398 387495 346454 387504
rect 346504 386414 346532 396034
rect 346596 393446 346624 399724
rect 346780 399650 346808 399758
rect 346918 399684 346946 400044
rect 347010 399906 347038 400044
rect 346998 399900 347050 399906
rect 346998 399842 347050 399848
rect 347102 399752 347130 400044
rect 347194 399906 347222 400044
rect 347286 399945 347314 400044
rect 347272 399936 347328 399945
rect 347182 399900 347234 399906
rect 347378 399906 347406 400044
rect 347470 399945 347498 400044
rect 347456 399936 347512 399945
rect 347272 399871 347328 399880
rect 347366 399900 347418 399906
rect 347182 399842 347234 399848
rect 347456 399871 347512 399880
rect 347366 399842 347418 399848
rect 347562 399838 347590 400044
rect 347654 399838 347682 400044
rect 347746 399911 347774 400044
rect 347732 399902 347788 399911
rect 347838 399906 347866 400044
rect 347930 399906 347958 400044
rect 348022 399945 348050 400044
rect 348008 399936 348064 399945
rect 347550 399832 347602 399838
rect 347410 399800 347466 399809
rect 346688 399622 346808 399650
rect 346872 399656 346946 399684
rect 347056 399724 347130 399752
rect 347228 399764 347280 399770
rect 346688 393514 346716 399622
rect 346768 399424 346820 399430
rect 346768 399366 346820 399372
rect 346780 399129 346808 399366
rect 346766 399120 346822 399129
rect 346766 399055 346822 399064
rect 346872 396098 346900 399656
rect 346952 399424 347004 399430
rect 346952 399366 347004 399372
rect 346964 397526 346992 399366
rect 346952 397520 347004 397526
rect 346952 397462 347004 397468
rect 346860 396092 346912 396098
rect 346860 396034 346912 396040
rect 346860 395412 346912 395418
rect 346860 395354 346912 395360
rect 346676 393508 346728 393514
rect 346676 393450 346728 393456
rect 346584 393440 346636 393446
rect 346584 393382 346636 393388
rect 346768 393304 346820 393310
rect 346768 393246 346820 393252
rect 346504 386386 346624 386414
rect 346216 384804 346268 384810
rect 346216 384746 346268 384752
rect 346122 321192 346178 321201
rect 346122 321127 346178 321136
rect 346032 317960 346084 317966
rect 346032 317902 346084 317908
rect 346228 311438 346256 384746
rect 346306 326632 346362 326641
rect 346306 326567 346362 326576
rect 346320 325825 346348 326567
rect 346306 325816 346362 325825
rect 346306 325751 346362 325760
rect 346596 319802 346624 386386
rect 346780 319841 346808 393246
rect 346872 386414 346900 395354
rect 347056 394058 347084 399724
rect 347228 399706 347280 399712
rect 347320 399764 347372 399770
rect 347550 399774 347602 399780
rect 347642 399832 347694 399838
rect 347732 399837 347788 399846
rect 347826 399900 347878 399906
rect 347826 399842 347878 399848
rect 347918 399900 347970 399906
rect 348008 399871 348064 399880
rect 347918 399842 347970 399848
rect 348114 399820 348142 400044
rect 348206 399906 348234 400044
rect 348298 399906 348326 400044
rect 348390 399945 348418 400044
rect 348376 399936 348432 399945
rect 348194 399900 348246 399906
rect 348194 399842 348246 399848
rect 348286 399900 348338 399906
rect 348376 399871 348432 399880
rect 348286 399842 348338 399848
rect 348482 399820 348510 400044
rect 347642 399774 347694 399780
rect 347962 399800 348018 399809
rect 347410 399735 347466 399744
rect 347780 399764 347832 399770
rect 347320 399706 347372 399712
rect 347136 399560 347188 399566
rect 347136 399502 347188 399508
rect 347044 394052 347096 394058
rect 347044 393994 347096 394000
rect 347044 392760 347096 392766
rect 347044 392702 347096 392708
rect 346872 386386 346992 386414
rect 346766 319832 346822 319841
rect 346584 319796 346636 319802
rect 346766 319767 346822 319776
rect 346584 319738 346636 319744
rect 346964 319161 346992 386386
rect 346950 319152 347006 319161
rect 346950 319087 347006 319096
rect 346216 311432 346268 311438
rect 346216 311374 346268 311380
rect 345940 304496 345992 304502
rect 345940 304438 345992 304444
rect 345848 300144 345900 300150
rect 345848 300086 345900 300092
rect 345756 297628 345808 297634
rect 345756 297570 345808 297576
rect 347056 295254 347084 392702
rect 347148 389842 347176 399502
rect 347240 398392 347268 399706
rect 347332 399265 347360 399706
rect 347318 399256 347374 399265
rect 347318 399191 347374 399200
rect 347240 398364 347360 398392
rect 347332 393310 347360 398364
rect 347424 395418 347452 399735
rect 347962 399735 348018 399744
rect 348068 399792 348142 399820
rect 348436 399792 348510 399820
rect 347780 399706 347832 399712
rect 347504 399696 347556 399702
rect 347504 399638 347556 399644
rect 347412 395412 347464 395418
rect 347412 395354 347464 395360
rect 347516 393582 347544 399638
rect 347596 399628 347648 399634
rect 347596 399570 347648 399576
rect 347504 393576 347556 393582
rect 347504 393518 347556 393524
rect 347320 393304 347372 393310
rect 347320 393246 347372 393252
rect 347136 389836 347188 389842
rect 347136 389778 347188 389784
rect 347136 389564 347188 389570
rect 347136 389506 347188 389512
rect 347148 307426 347176 389506
rect 347502 388512 347558 388521
rect 347608 388482 347636 399570
rect 347792 399265 347820 399706
rect 347872 399696 347924 399702
rect 347872 399638 347924 399644
rect 347778 399256 347834 399265
rect 347778 399191 347834 399200
rect 347778 398848 347834 398857
rect 347778 398783 347834 398792
rect 347792 398750 347820 398783
rect 347780 398744 347832 398750
rect 347780 398686 347832 398692
rect 347884 388929 347912 399638
rect 347976 395554 348004 399735
rect 348068 399498 348096 399792
rect 348240 399764 348292 399770
rect 348240 399706 348292 399712
rect 348148 399696 348200 399702
rect 348148 399638 348200 399644
rect 348056 399492 348108 399498
rect 348056 399434 348108 399440
rect 348160 398936 348188 399638
rect 348068 398908 348188 398936
rect 347964 395548 348016 395554
rect 347964 395490 348016 395496
rect 347964 393440 348016 393446
rect 347964 393382 348016 393388
rect 347870 388920 347926 388929
rect 347870 388855 347926 388864
rect 347502 388447 347558 388456
rect 347596 388476 347648 388482
rect 347320 387252 347372 387258
rect 347320 387194 347372 387200
rect 347226 381712 347282 381721
rect 347226 381647 347282 381656
rect 347136 307420 347188 307426
rect 347136 307362 347188 307368
rect 347240 297702 347268 381647
rect 347332 304638 347360 387194
rect 347412 384532 347464 384538
rect 347412 384474 347464 384480
rect 347424 311098 347452 384474
rect 347516 372026 347544 388447
rect 347596 388418 347648 388424
rect 347976 374785 348004 393382
rect 348068 388550 348096 398908
rect 348148 398812 348200 398818
rect 348148 398754 348200 398760
rect 348160 398342 348188 398754
rect 348148 398336 348200 398342
rect 348148 398278 348200 398284
rect 348252 391270 348280 399706
rect 348332 399696 348384 399702
rect 348332 399638 348384 399644
rect 348344 398410 348372 399638
rect 348436 399566 348464 399792
rect 348574 399752 348602 400044
rect 348528 399724 348602 399752
rect 348528 399566 348556 399724
rect 348666 399684 348694 400044
rect 348758 399838 348786 400044
rect 348850 399906 348878 400044
rect 348838 399900 348890 399906
rect 348838 399842 348890 399848
rect 348746 399832 348798 399838
rect 348746 399774 348798 399780
rect 348942 399752 348970 400044
rect 349034 399838 349062 400044
rect 349022 399832 349074 399838
rect 349126 399809 349154 400044
rect 349218 399945 349246 400044
rect 349204 399936 349260 399945
rect 349204 399871 349260 399880
rect 349310 399820 349338 400044
rect 349022 399774 349074 399780
rect 349112 399800 349168 399809
rect 348896 399724 348970 399752
rect 349112 399735 349168 399744
rect 349264 399792 349338 399820
rect 348620 399656 348694 399684
rect 348792 399696 348844 399702
rect 348424 399560 348476 399566
rect 348424 399502 348476 399508
rect 348516 399560 348568 399566
rect 348516 399502 348568 399508
rect 348424 399288 348476 399294
rect 348424 399230 348476 399236
rect 348436 399129 348464 399230
rect 348422 399120 348478 399129
rect 348422 399055 348478 399064
rect 348516 399016 348568 399022
rect 348516 398958 348568 398964
rect 348528 398750 348556 398958
rect 348516 398744 348568 398750
rect 348516 398686 348568 398692
rect 348332 398404 348384 398410
rect 348332 398346 348384 398352
rect 348424 397792 348476 397798
rect 348424 397734 348476 397740
rect 348240 391264 348292 391270
rect 348240 391206 348292 391212
rect 348056 388544 348108 388550
rect 348056 388486 348108 388492
rect 347962 374776 348018 374785
rect 347962 374711 348018 374720
rect 347504 372020 347556 372026
rect 347504 371962 347556 371968
rect 347504 316872 347556 316878
rect 347504 316814 347556 316820
rect 347516 316742 347544 316814
rect 347504 316736 347556 316742
rect 347504 316678 347556 316684
rect 347412 311092 347464 311098
rect 347412 311034 347464 311040
rect 347320 304632 347372 304638
rect 347320 304574 347372 304580
rect 347228 297696 347280 297702
rect 347228 297638 347280 297644
rect 347044 295248 347096 295254
rect 347044 295190 347096 295196
rect 347516 262886 347544 316678
rect 348436 307562 348464 397734
rect 348620 394694 348648 399656
rect 348792 399638 348844 399644
rect 348700 399220 348752 399226
rect 348700 399162 348752 399168
rect 348712 399129 348740 399162
rect 348698 399120 348754 399129
rect 348698 399055 348754 399064
rect 348700 398812 348752 398818
rect 348700 398754 348752 398760
rect 348712 398313 348740 398754
rect 348698 398304 348754 398313
rect 348698 398239 348754 398248
rect 348528 394666 348648 394694
rect 348528 393417 348556 394666
rect 348700 393576 348752 393582
rect 348700 393518 348752 393524
rect 348514 393408 348570 393417
rect 348514 393343 348570 393352
rect 348516 387796 348568 387802
rect 348516 387738 348568 387744
rect 348424 307556 348476 307562
rect 348424 307498 348476 307504
rect 348528 304570 348556 387738
rect 348608 387660 348660 387666
rect 348608 387602 348660 387608
rect 348516 304564 348568 304570
rect 348516 304506 348568 304512
rect 348620 304298 348648 387602
rect 348712 386414 348740 393518
rect 348804 393310 348832 399638
rect 348792 393304 348844 393310
rect 348792 393246 348844 393252
rect 348896 392766 348924 399724
rect 349068 399696 349120 399702
rect 349068 399638 349120 399644
rect 349160 399696 349212 399702
rect 349160 399638 349212 399644
rect 348976 399628 349028 399634
rect 348976 399570 349028 399576
rect 348884 392760 348936 392766
rect 348884 392702 348936 392708
rect 348712 386386 348832 386414
rect 348700 384872 348752 384878
rect 348700 384814 348752 384820
rect 348712 305862 348740 384814
rect 348804 318986 348832 386386
rect 348882 377904 348938 377913
rect 348882 377839 348938 377848
rect 348792 318980 348844 318986
rect 348792 318922 348844 318928
rect 348792 316736 348844 316742
rect 348792 316678 348844 316684
rect 348700 305856 348752 305862
rect 348700 305798 348752 305804
rect 348608 304292 348660 304298
rect 348608 304234 348660 304240
rect 347504 262880 347556 262886
rect 347504 262822 347556 262828
rect 348804 239426 348832 316678
rect 348896 308718 348924 377839
rect 348884 308712 348936 308718
rect 348884 308654 348936 308660
rect 348988 296682 349016 399570
rect 349080 393446 349108 399638
rect 349172 397372 349200 399638
rect 349264 398614 349292 399792
rect 349402 399752 349430 400044
rect 349494 399838 349522 400044
rect 349586 399838 349614 400044
rect 349678 399838 349706 400044
rect 349482 399832 349534 399838
rect 349482 399774 349534 399780
rect 349574 399832 349626 399838
rect 349574 399774 349626 399780
rect 349666 399832 349718 399838
rect 349666 399774 349718 399780
rect 349356 399724 349430 399752
rect 349252 398608 349304 398614
rect 349252 398550 349304 398556
rect 349172 397344 349292 397372
rect 349160 396976 349212 396982
rect 349160 396918 349212 396924
rect 349068 393440 349120 393446
rect 349068 393382 349120 393388
rect 349068 393304 349120 393310
rect 349068 393246 349120 393252
rect 349080 298110 349108 393246
rect 349172 392902 349200 396918
rect 349264 393582 349292 397344
rect 349252 393576 349304 393582
rect 349252 393518 349304 393524
rect 349356 393417 349384 399724
rect 349528 399696 349580 399702
rect 349770 399684 349798 400044
rect 349862 399838 349890 400044
rect 349954 399838 349982 400044
rect 349850 399832 349902 399838
rect 349850 399774 349902 399780
rect 349942 399832 349994 399838
rect 350046 399809 350074 400044
rect 350138 399838 350166 400044
rect 350126 399832 350178 399838
rect 349942 399774 349994 399780
rect 350032 399800 350088 399809
rect 350126 399774 350178 399780
rect 350032 399735 350088 399744
rect 349528 399638 349580 399644
rect 349724 399656 349798 399684
rect 350080 399696 350132 399702
rect 349436 399628 349488 399634
rect 349436 399570 349488 399576
rect 349448 397730 349476 399570
rect 349436 397724 349488 397730
rect 349436 397666 349488 397672
rect 349436 397520 349488 397526
rect 349436 397462 349488 397468
rect 349342 393408 349398 393417
rect 349342 393343 349398 393352
rect 349252 393304 349304 393310
rect 349252 393246 349304 393252
rect 349160 392896 349212 392902
rect 349160 392838 349212 392844
rect 349264 348430 349292 393246
rect 349344 392896 349396 392902
rect 349344 392838 349396 392844
rect 349356 358057 349384 392838
rect 349448 378729 349476 397462
rect 349540 396982 349568 399638
rect 349620 399424 349672 399430
rect 349620 399366 349672 399372
rect 349632 399226 349660 399366
rect 349620 399220 349672 399226
rect 349620 399162 349672 399168
rect 349620 397860 349672 397866
rect 349620 397802 349672 397808
rect 349528 396976 349580 396982
rect 349528 396918 349580 396924
rect 349528 393440 349580 393446
rect 349528 393382 349580 393388
rect 349540 379273 349568 393382
rect 349526 379264 349582 379273
rect 349526 379199 349582 379208
rect 349434 378720 349490 378729
rect 349434 378655 349490 378664
rect 349342 358048 349398 358057
rect 349342 357983 349398 357992
rect 349252 348424 349304 348430
rect 349252 348366 349304 348372
rect 349632 342922 349660 397802
rect 349724 397526 349752 399656
rect 350080 399638 350132 399644
rect 349804 399560 349856 399566
rect 349804 399502 349856 399508
rect 349712 397520 349764 397526
rect 349712 397462 349764 397468
rect 349816 393446 349844 399502
rect 349896 399492 349948 399498
rect 349896 399434 349948 399440
rect 349804 393440 349856 393446
rect 349804 393382 349856 393388
rect 349908 392748 349936 399434
rect 349988 399016 350040 399022
rect 349988 398958 350040 398964
rect 350000 398886 350028 398958
rect 349988 398880 350040 398886
rect 349988 398822 350040 398828
rect 350092 397866 350120 399638
rect 350230 399616 350258 400044
rect 350322 399838 350350 400044
rect 350414 399945 350442 400044
rect 350400 399936 350456 399945
rect 350400 399871 350456 399880
rect 350506 399838 350534 400044
rect 350598 399906 350626 400044
rect 350690 399906 350718 400044
rect 350782 399945 350810 400044
rect 350768 399936 350824 399945
rect 350586 399900 350638 399906
rect 350586 399842 350638 399848
rect 350678 399900 350730 399906
rect 350768 399871 350824 399880
rect 350678 399842 350730 399848
rect 350310 399832 350362 399838
rect 350310 399774 350362 399780
rect 350494 399832 350546 399838
rect 350494 399774 350546 399780
rect 350632 399764 350684 399770
rect 350632 399706 350684 399712
rect 350724 399764 350776 399770
rect 350874 399752 350902 400044
rect 350966 399906 350994 400044
rect 351058 399945 351086 400044
rect 351044 399936 351100 399945
rect 350954 399900 351006 399906
rect 351044 399871 351100 399880
rect 350954 399842 351006 399848
rect 350724 399706 350776 399712
rect 350828 399724 350902 399752
rect 350184 399588 350258 399616
rect 350448 399628 350500 399634
rect 350080 397860 350132 397866
rect 350080 397802 350132 397808
rect 350080 397724 350132 397730
rect 350080 397666 350132 397672
rect 350092 392834 350120 397666
rect 350080 392828 350132 392834
rect 350080 392770 350132 392776
rect 349908 392720 350028 392748
rect 349804 389360 349856 389366
rect 349804 389302 349856 389308
rect 349620 342916 349672 342922
rect 349620 342858 349672 342864
rect 349816 304706 349844 389302
rect 349896 388544 349948 388550
rect 349896 388486 349948 388492
rect 349908 305522 349936 388486
rect 350000 386034 350028 392720
rect 350184 390153 350212 399588
rect 350448 399570 350500 399576
rect 350264 399492 350316 399498
rect 350264 399434 350316 399440
rect 350276 392970 350304 399434
rect 350460 396914 350488 399570
rect 350538 397488 350594 397497
rect 350538 397423 350594 397432
rect 350448 396908 350500 396914
rect 350448 396850 350500 396856
rect 350552 393310 350580 397423
rect 350644 395010 350672 399706
rect 350632 395004 350684 395010
rect 350632 394946 350684 394952
rect 350632 393848 350684 393854
rect 350632 393790 350684 393796
rect 350540 393304 350592 393310
rect 350540 393246 350592 393252
rect 350264 392964 350316 392970
rect 350264 392906 350316 392912
rect 350170 390144 350226 390153
rect 350170 390079 350226 390088
rect 349988 386028 350040 386034
rect 349988 385970 350040 385976
rect 349986 382120 350042 382129
rect 349986 382055 350042 382064
rect 349896 305516 349948 305522
rect 349896 305458 349948 305464
rect 349804 304700 349856 304706
rect 349804 304642 349856 304648
rect 350000 300218 350028 382055
rect 350172 381540 350224 381546
rect 350172 381482 350224 381488
rect 350078 378040 350134 378049
rect 350078 377975 350134 377984
rect 350092 308786 350120 377975
rect 350184 312866 350212 381482
rect 350644 355366 350672 393790
rect 350736 393530 350764 399706
rect 350828 395282 350856 399724
rect 351150 399684 351178 400044
rect 351242 399838 351270 400044
rect 351230 399832 351282 399838
rect 351230 399774 351282 399780
rect 351104 399656 351178 399684
rect 351334 399684 351362 400044
rect 351426 399906 351454 400044
rect 351414 399900 351466 399906
rect 351414 399842 351466 399848
rect 351518 399684 351546 400044
rect 351610 399945 351638 400044
rect 351596 399936 351652 399945
rect 351702 399906 351730 400044
rect 351794 399945 351822 400044
rect 351780 399936 351836 399945
rect 351596 399871 351652 399880
rect 351690 399900 351742 399906
rect 351886 399906 351914 400044
rect 351978 399906 352006 400044
rect 351780 399871 351836 399880
rect 351874 399900 351926 399906
rect 351690 399842 351742 399848
rect 351874 399842 351926 399848
rect 351966 399900 352018 399906
rect 351966 399842 352018 399848
rect 351826 399800 351882 399809
rect 351644 399764 351696 399770
rect 352070 399786 352098 400044
rect 352162 399838 352190 400044
rect 352254 399906 352282 400044
rect 352242 399900 352294 399906
rect 352242 399842 352294 399848
rect 351826 399735 351882 399744
rect 352024 399758 352098 399786
rect 352150 399832 352202 399838
rect 352150 399774 352202 399780
rect 351644 399706 351696 399712
rect 351334 399656 351408 399684
rect 351518 399656 351592 399684
rect 351000 399628 351052 399634
rect 351000 399570 351052 399576
rect 350908 399424 350960 399430
rect 350908 399366 350960 399372
rect 350920 396001 350948 399366
rect 350906 395992 350962 396001
rect 350906 395927 350962 395936
rect 350908 395548 350960 395554
rect 350908 395490 350960 395496
rect 350816 395276 350868 395282
rect 350816 395218 350868 395224
rect 350736 393502 350856 393530
rect 350724 393304 350776 393310
rect 350724 393246 350776 393252
rect 350736 359417 350764 393246
rect 350828 378865 350856 393502
rect 350920 379409 350948 395490
rect 351012 393310 351040 399570
rect 351104 397934 351132 399656
rect 351184 399560 351236 399566
rect 351184 399502 351236 399508
rect 351092 397928 351144 397934
rect 351092 397870 351144 397876
rect 351092 397520 351144 397526
rect 351092 397462 351144 397468
rect 351000 393304 351052 393310
rect 351000 393246 351052 393252
rect 351104 390289 351132 397462
rect 351196 396710 351224 399502
rect 351380 397526 351408 399656
rect 351564 398698 351592 399656
rect 351472 398670 351592 398698
rect 351368 397520 351420 397526
rect 351368 397462 351420 397468
rect 351472 397372 351500 398670
rect 351552 398608 351604 398614
rect 351550 398576 351552 398585
rect 351604 398576 351606 398585
rect 351550 398511 351606 398520
rect 351380 397344 351500 397372
rect 351184 396704 351236 396710
rect 351184 396646 351236 396652
rect 351184 396228 351236 396234
rect 351184 396170 351236 396176
rect 351090 390280 351146 390289
rect 351090 390215 351146 390224
rect 351000 389020 351052 389026
rect 351000 388962 351052 388968
rect 350906 379400 350962 379409
rect 350906 379335 350962 379344
rect 351012 379137 351040 388962
rect 350998 379128 351054 379137
rect 350998 379063 351054 379072
rect 350814 378856 350870 378865
rect 350814 378791 350870 378800
rect 350722 359408 350778 359417
rect 350722 359343 350778 359352
rect 350632 355360 350684 355366
rect 350632 355302 350684 355308
rect 350172 312860 350224 312866
rect 350172 312802 350224 312808
rect 350080 308780 350132 308786
rect 350080 308722 350132 308728
rect 351196 303142 351224 396170
rect 351380 393854 351408 397344
rect 351656 394694 351684 399706
rect 351736 399696 351788 399702
rect 351736 399638 351788 399644
rect 351748 395554 351776 399638
rect 351736 395548 351788 395554
rect 351736 395490 351788 395496
rect 351472 394666 351684 394694
rect 351368 393848 351420 393854
rect 351368 393790 351420 393796
rect 351368 393508 351420 393514
rect 351368 393450 351420 393456
rect 351276 389768 351328 389774
rect 351276 389710 351328 389716
rect 351288 304774 351316 389710
rect 351380 307630 351408 393450
rect 351472 389026 351500 394666
rect 351460 389020 351512 389026
rect 351460 388962 351512 388968
rect 351840 386414 351868 399735
rect 352024 399684 352052 399758
rect 352346 399752 352374 400044
rect 352438 399906 352466 400044
rect 352530 399906 352558 400044
rect 352426 399900 352478 399906
rect 352426 399842 352478 399848
rect 352518 399900 352570 399906
rect 352518 399842 352570 399848
rect 352300 399724 352374 399752
rect 352470 399800 352526 399809
rect 352622 399752 352650 400044
rect 352470 399735 352526 399744
rect 351932 399656 352052 399684
rect 352104 399696 352156 399702
rect 351932 393938 351960 399656
rect 352104 399638 352156 399644
rect 352012 399560 352064 399566
rect 352012 399502 352064 399508
rect 352024 396574 352052 399502
rect 352116 398818 352144 399638
rect 352196 399628 352248 399634
rect 352196 399570 352248 399576
rect 352104 398812 352156 398818
rect 352104 398754 352156 398760
rect 352104 398336 352156 398342
rect 352104 398278 352156 398284
rect 352116 397934 352144 398278
rect 352104 397928 352156 397934
rect 352104 397870 352156 397876
rect 352012 396568 352064 396574
rect 352012 396510 352064 396516
rect 352208 394694 352236 399570
rect 352300 395457 352328 399724
rect 352380 399628 352432 399634
rect 352380 399570 352432 399576
rect 352392 397798 352420 399570
rect 352484 399498 352512 399735
rect 352576 399724 352650 399752
rect 352472 399492 352524 399498
rect 352472 399434 352524 399440
rect 352472 397996 352524 398002
rect 352472 397938 352524 397944
rect 352380 397792 352432 397798
rect 352380 397734 352432 397740
rect 352378 396808 352434 396817
rect 352378 396743 352434 396752
rect 352392 396409 352420 396743
rect 352378 396400 352434 396409
rect 352378 396335 352434 396344
rect 352286 395448 352342 395457
rect 352286 395383 352342 395392
rect 352208 394666 352328 394694
rect 351932 393910 352236 393938
rect 352104 393848 352156 393854
rect 352104 393790 352156 393796
rect 351656 386386 351868 386414
rect 351550 381848 351606 381857
rect 351550 381783 351606 381792
rect 351460 377460 351512 377466
rect 351460 377402 351512 377408
rect 351368 307624 351420 307630
rect 351368 307566 351420 307572
rect 351276 304768 351328 304774
rect 351276 304710 351328 304716
rect 351184 303136 351236 303142
rect 351184 303078 351236 303084
rect 351472 301510 351500 377402
rect 351564 311166 351592 381783
rect 351656 349858 351684 386386
rect 351644 349852 351696 349858
rect 351644 349794 351696 349800
rect 352116 319122 352144 393790
rect 352208 358086 352236 393910
rect 352300 379001 352328 394666
rect 352380 394052 352432 394058
rect 352380 393994 352432 394000
rect 352286 378992 352342 379001
rect 352286 378927 352342 378936
rect 352196 358080 352248 358086
rect 352196 358022 352248 358028
rect 352104 319116 352156 319122
rect 352104 319058 352156 319064
rect 352392 311710 352420 393994
rect 352484 319394 352512 397938
rect 352576 393854 352604 399724
rect 352714 399684 352742 400044
rect 352668 399656 352742 399684
rect 352806 399684 352834 400044
rect 352898 399809 352926 400044
rect 352884 399800 352940 399809
rect 352884 399735 352940 399744
rect 352990 399684 353018 400044
rect 352806 399656 352880 399684
rect 352668 394058 352696 399656
rect 352748 399560 352800 399566
rect 352748 399502 352800 399508
rect 352760 395350 352788 399502
rect 352852 398002 352880 399656
rect 352944 399656 353018 399684
rect 353082 399684 353110 400044
rect 353174 399786 353202 400044
rect 353266 399906 353294 400044
rect 353254 399900 353306 399906
rect 353254 399842 353306 399848
rect 353358 399820 353386 400044
rect 353450 399945 353478 400044
rect 353436 399936 353492 399945
rect 353436 399871 353492 399880
rect 353358 399792 353432 399820
rect 353174 399758 353248 399786
rect 353082 399656 353156 399684
rect 352840 397996 352892 398002
rect 352840 397938 352892 397944
rect 352944 397576 352972 399656
rect 352852 397548 352972 397576
rect 352748 395344 352800 395350
rect 352748 395286 352800 395292
rect 352748 394256 352800 394262
rect 352748 394198 352800 394204
rect 352656 394052 352708 394058
rect 352656 393994 352708 394000
rect 352564 393848 352616 393854
rect 352564 393790 352616 393796
rect 352760 392850 352788 394198
rect 352668 392822 352788 392850
rect 352564 387932 352616 387938
rect 352564 387874 352616 387880
rect 352472 319388 352524 319394
rect 352472 319330 352524 319336
rect 352380 311704 352432 311710
rect 352380 311646 352432 311652
rect 351552 311160 351604 311166
rect 351552 311102 351604 311108
rect 352576 303074 352604 387874
rect 352668 314838 352696 392822
rect 352748 392760 352800 392766
rect 352748 392702 352800 392708
rect 352760 317257 352788 392702
rect 352852 384334 352880 397548
rect 352930 397488 352986 397497
rect 352930 397423 352986 397432
rect 352944 389174 352972 397423
rect 353128 396846 353156 399656
rect 353116 396840 353168 396846
rect 353116 396782 353168 396788
rect 353024 395004 353076 395010
rect 353024 394946 353076 394952
rect 353036 391105 353064 394946
rect 353220 392698 353248 399758
rect 353300 399696 353352 399702
rect 353300 399638 353352 399644
rect 353312 399401 353340 399638
rect 353298 399392 353354 399401
rect 353298 399327 353354 399336
rect 353404 393310 353432 399792
rect 353542 399752 353570 400044
rect 353634 399906 353662 400044
rect 353622 399900 353674 399906
rect 353622 399842 353674 399848
rect 353726 399752 353754 400044
rect 353818 399906 353846 400044
rect 353806 399900 353858 399906
rect 353806 399842 353858 399848
rect 353910 399838 353938 400044
rect 354002 399945 354030 400044
rect 353988 399936 354044 399945
rect 353988 399871 354044 399880
rect 354094 399838 354122 400044
rect 354186 399945 354214 400044
rect 354172 399936 354228 399945
rect 354278 399906 354306 400044
rect 354172 399871 354228 399880
rect 354266 399900 354318 399906
rect 354266 399842 354318 399848
rect 353898 399832 353950 399838
rect 353898 399774 353950 399780
rect 354082 399832 354134 399838
rect 354082 399774 354134 399780
rect 353542 399724 353616 399752
rect 353726 399724 353800 399752
rect 353482 399392 353538 399401
rect 353482 399327 353538 399336
rect 353496 399226 353524 399327
rect 353484 399220 353536 399226
rect 353484 399162 353536 399168
rect 353484 398132 353536 398138
rect 353484 398074 353536 398080
rect 353496 397594 353524 398074
rect 353484 397588 353536 397594
rect 353484 397530 353536 397536
rect 353482 397216 353538 397225
rect 353482 397151 353538 397160
rect 353496 396817 353524 397151
rect 353482 396808 353538 396817
rect 353482 396743 353538 396752
rect 353484 395276 353536 395282
rect 353484 395218 353536 395224
rect 353392 393304 353444 393310
rect 353392 393246 353444 393252
rect 353208 392692 353260 392698
rect 353208 392634 353260 392640
rect 353022 391096 353078 391105
rect 353022 391031 353078 391040
rect 352944 389146 353064 389174
rect 353036 385830 353064 389146
rect 353496 386414 353524 395218
rect 353588 392426 353616 399724
rect 353668 399628 353720 399634
rect 353668 399570 353720 399576
rect 353680 395486 353708 399570
rect 353668 395480 353720 395486
rect 353668 395422 353720 395428
rect 353576 392420 353628 392426
rect 353576 392362 353628 392368
rect 353772 386414 353800 399724
rect 354220 399628 354272 399634
rect 354370 399616 354398 400044
rect 354462 399838 354490 400044
rect 354450 399832 354502 399838
rect 354450 399774 354502 399780
rect 354554 399684 354582 400044
rect 354646 399838 354674 400044
rect 354738 399906 354766 400044
rect 354726 399900 354778 399906
rect 354726 399842 354778 399848
rect 354634 399832 354686 399838
rect 354634 399774 354686 399780
rect 354830 399752 354858 400044
rect 354922 399906 354950 400044
rect 354910 399900 354962 399906
rect 354910 399842 354962 399848
rect 354784 399724 354858 399752
rect 354220 399570 354272 399576
rect 354324 399588 354398 399616
rect 354508 399656 354582 399684
rect 354680 399696 354732 399702
rect 353852 399560 353904 399566
rect 353852 399502 353904 399508
rect 354128 399560 354180 399566
rect 354128 399502 354180 399508
rect 353864 393514 353892 399502
rect 353944 399492 353996 399498
rect 353944 399434 353996 399440
rect 353852 393508 353904 393514
rect 353852 393450 353904 393456
rect 353404 386386 353524 386414
rect 353588 386386 353800 386414
rect 353024 385824 353076 385830
rect 353024 385766 353076 385772
rect 352840 384328 352892 384334
rect 352840 384270 352892 384276
rect 353404 319258 353432 386386
rect 353588 381585 353616 386386
rect 353574 381576 353630 381585
rect 353574 381511 353630 381520
rect 353392 319252 353444 319258
rect 353392 319194 353444 319200
rect 352746 317248 352802 317257
rect 352746 317183 352802 317192
rect 352656 314832 352708 314838
rect 352656 314774 352708 314780
rect 352564 303068 352616 303074
rect 352564 303010 352616 303016
rect 351460 301504 351512 301510
rect 351460 301446 351512 301452
rect 349988 300212 350040 300218
rect 349988 300154 350040 300160
rect 353956 299334 353984 399434
rect 354036 399220 354088 399226
rect 354036 399162 354088 399168
rect 354048 399129 354076 399162
rect 354034 399120 354090 399129
rect 354034 399055 354090 399064
rect 354036 398812 354088 398818
rect 354036 398754 354088 398760
rect 354048 303210 354076 398754
rect 354140 394312 354168 399502
rect 354232 395010 354260 399570
rect 354324 395282 354352 399588
rect 354404 399424 354456 399430
rect 354404 399366 354456 399372
rect 354416 399265 354444 399366
rect 354402 399256 354458 399265
rect 354402 399191 354458 399200
rect 354404 398880 354456 398886
rect 354404 398822 354456 398828
rect 354416 398478 354444 398822
rect 354404 398472 354456 398478
rect 354404 398414 354456 398420
rect 354508 398206 354536 399656
rect 354680 399638 354732 399644
rect 354588 399356 354640 399362
rect 354588 399298 354640 399304
rect 354600 399265 354628 399298
rect 354586 399256 354642 399265
rect 354586 399191 354642 399200
rect 354588 398336 354640 398342
rect 354588 398278 354640 398284
rect 354496 398200 354548 398206
rect 354496 398142 354548 398148
rect 354600 397934 354628 398278
rect 354588 397928 354640 397934
rect 354588 397870 354640 397876
rect 354496 396840 354548 396846
rect 354496 396782 354548 396788
rect 354312 395276 354364 395282
rect 354312 395218 354364 395224
rect 354220 395004 354272 395010
rect 354220 394946 354272 394952
rect 354140 394284 354444 394312
rect 354128 394188 354180 394194
rect 354128 394130 354180 394136
rect 354140 309738 354168 394130
rect 354312 393304 354364 393310
rect 354312 393246 354364 393252
rect 354220 388476 354272 388482
rect 354220 388418 354272 388424
rect 354232 318034 354260 388418
rect 354324 320890 354352 393246
rect 354312 320884 354364 320890
rect 354312 320826 354364 320832
rect 354416 319326 354444 394284
rect 354508 389570 354536 396782
rect 354692 396001 354720 399638
rect 354784 399634 354812 399724
rect 355014 399684 355042 400044
rect 355106 399838 355134 400044
rect 355094 399832 355146 399838
rect 355094 399774 355146 399780
rect 355198 399684 355226 400044
rect 355290 399786 355318 400044
rect 355382 399945 355410 400044
rect 355368 399936 355424 399945
rect 355368 399871 355424 399880
rect 355474 399786 355502 400044
rect 355566 399906 355594 400044
rect 355554 399900 355606 399906
rect 355554 399842 355606 399848
rect 355290 399758 355364 399786
rect 354968 399656 355042 399684
rect 355152 399656 355226 399684
rect 354772 399628 354824 399634
rect 354772 399570 354824 399576
rect 354864 399628 354916 399634
rect 354864 399570 354916 399576
rect 354772 399424 354824 399430
rect 354772 399366 354824 399372
rect 354784 396166 354812 399366
rect 354772 396160 354824 396166
rect 354772 396102 354824 396108
rect 354678 395992 354734 396001
rect 354876 395978 354904 399570
rect 354968 396846 354996 399656
rect 355152 399480 355180 399656
rect 355060 399452 355180 399480
rect 355232 399492 355284 399498
rect 355060 397662 355088 399452
rect 355232 399434 355284 399440
rect 355140 399356 355192 399362
rect 355140 399298 355192 399304
rect 355048 397656 355100 397662
rect 355048 397598 355100 397604
rect 355152 397372 355180 399298
rect 355060 397344 355180 397372
rect 354956 396840 355008 396846
rect 354956 396782 355008 396788
rect 354876 395950 354996 395978
rect 354678 395927 354734 395936
rect 354864 395412 354916 395418
rect 354864 395354 354916 395360
rect 354496 389564 354548 389570
rect 354496 389506 354548 389512
rect 354876 387938 354904 395354
rect 354968 391066 354996 395950
rect 354956 391060 355008 391066
rect 354956 391002 355008 391008
rect 354864 387932 354916 387938
rect 354864 387874 354916 387880
rect 354404 319320 354456 319326
rect 354404 319262 354456 319268
rect 354220 318028 354272 318034
rect 354220 317970 354272 317976
rect 355060 316538 355088 397344
rect 355140 396772 355192 396778
rect 355140 396714 355192 396720
rect 355152 389366 355180 396714
rect 355244 394058 355272 399434
rect 355336 396234 355364 399758
rect 355428 399758 355502 399786
rect 355428 399673 355456 399758
rect 355658 399752 355686 400044
rect 355612 399724 355686 399752
rect 355508 399696 355560 399702
rect 355414 399664 355470 399673
rect 355508 399638 355560 399644
rect 355414 399599 355470 399608
rect 355416 399560 355468 399566
rect 355416 399502 355468 399508
rect 355428 398818 355456 399502
rect 355416 398812 355468 398818
rect 355416 398754 355468 398760
rect 355520 398698 355548 399638
rect 355428 398670 355548 398698
rect 355324 396228 355376 396234
rect 355324 396170 355376 396176
rect 355232 394052 355284 394058
rect 355232 393994 355284 394000
rect 355428 393224 355456 398670
rect 355508 398540 355560 398546
rect 355508 398482 355560 398488
rect 355244 393196 355456 393224
rect 355140 389360 355192 389366
rect 355140 389302 355192 389308
rect 355244 387598 355272 393196
rect 355520 393122 355548 398482
rect 355612 397594 355640 399724
rect 355750 399684 355778 400044
rect 355842 399752 355870 400044
rect 355934 399906 355962 400044
rect 355922 399900 355974 399906
rect 355922 399842 355974 399848
rect 356026 399752 356054 400044
rect 355842 399724 355916 399752
rect 355750 399656 355824 399684
rect 355692 399356 355744 399362
rect 355692 399298 355744 399304
rect 355600 397588 355652 397594
rect 355600 397530 355652 397536
rect 355704 397372 355732 399298
rect 355796 398721 355824 399656
rect 355888 399566 355916 399724
rect 355980 399724 356054 399752
rect 355876 399560 355928 399566
rect 355876 399502 355928 399508
rect 355876 399424 355928 399430
rect 355876 399366 355928 399372
rect 355888 398886 355916 399366
rect 355980 398954 356008 399724
rect 356118 399684 356146 400044
rect 356210 399752 356238 400044
rect 356302 399906 356330 400044
rect 356290 399900 356342 399906
rect 356290 399842 356342 399848
rect 356394 399786 356422 400044
rect 356348 399758 356422 399786
rect 356210 399724 356284 399752
rect 356072 399656 356146 399684
rect 355968 398948 356020 398954
rect 355968 398890 356020 398896
rect 355876 398880 355928 398886
rect 355876 398822 355928 398828
rect 355782 398712 355838 398721
rect 355782 398647 355838 398656
rect 355612 397344 355732 397372
rect 355612 394369 355640 397344
rect 355692 396908 355744 396914
rect 355692 396850 355744 396856
rect 355598 394360 355654 394369
rect 355598 394295 355654 394304
rect 355598 393816 355654 393825
rect 355598 393751 355654 393760
rect 355336 393094 355548 393122
rect 355232 387592 355284 387598
rect 355232 387534 355284 387540
rect 355048 316532 355100 316538
rect 355048 316474 355100 316480
rect 355336 310010 355364 393094
rect 355612 392170 355640 393751
rect 355428 392142 355640 392170
rect 355324 310004 355376 310010
rect 355324 309946 355376 309952
rect 354128 309732 354180 309738
rect 354128 309674 354180 309680
rect 355428 307154 355456 392142
rect 355508 392080 355560 392086
rect 355704 392034 355732 396850
rect 355876 396500 355928 396506
rect 355876 396442 355928 396448
rect 355508 392022 355560 392028
rect 355520 308650 355548 392022
rect 355612 392006 355732 392034
rect 355612 311574 355640 392006
rect 355888 389174 355916 396442
rect 356072 395418 356100 399656
rect 356152 399560 356204 399566
rect 356152 399502 356204 399508
rect 356164 399401 356192 399502
rect 356150 399392 356206 399401
rect 356256 399362 356284 399724
rect 356348 399616 356376 399758
rect 356486 399752 356514 400044
rect 356578 399906 356606 400044
rect 356566 399900 356618 399906
rect 356566 399842 356618 399848
rect 356670 399786 356698 400044
rect 356624 399770 356698 399786
rect 356612 399764 356698 399770
rect 356486 399724 356560 399752
rect 356532 399650 356560 399724
rect 356664 399758 356698 399764
rect 356612 399706 356664 399712
rect 356762 399684 356790 400044
rect 356854 399906 356882 400044
rect 356842 399900 356894 399906
rect 356842 399842 356894 399848
rect 356946 399752 356974 400044
rect 356716 399656 356790 399684
rect 356900 399724 356974 399752
rect 356900 399673 356928 399724
rect 357038 399684 357066 400044
rect 357130 399906 357158 400044
rect 357118 399900 357170 399906
rect 357118 399842 357170 399848
rect 357222 399752 357250 400044
rect 356886 399664 356942 399673
rect 356532 399622 356652 399650
rect 356348 399588 356468 399616
rect 356440 399498 356468 399588
rect 356520 399560 356572 399566
rect 356520 399502 356572 399508
rect 356336 399492 356388 399498
rect 356336 399434 356388 399440
rect 356428 399492 356480 399498
rect 356428 399434 356480 399440
rect 356150 399327 356206 399336
rect 356244 399356 356296 399362
rect 356244 399298 356296 399304
rect 356152 398948 356204 398954
rect 356152 398890 356204 398896
rect 356060 395412 356112 395418
rect 356060 395354 356112 395360
rect 355968 395344 356020 395350
rect 355968 395286 356020 395292
rect 355704 389146 355916 389174
rect 355704 387802 355732 389146
rect 355692 387796 355744 387802
rect 355692 387738 355744 387744
rect 355600 311568 355652 311574
rect 355600 311510 355652 311516
rect 355508 308644 355560 308650
rect 355508 308586 355560 308592
rect 355416 307148 355468 307154
rect 355416 307090 355468 307096
rect 354036 303204 354088 303210
rect 354036 303146 354088 303152
rect 353944 299328 353996 299334
rect 353944 299270 353996 299276
rect 349068 298104 349120 298110
rect 349068 298046 349120 298052
rect 348976 296676 349028 296682
rect 348976 296618 349028 296624
rect 355980 291922 356008 395286
rect 356164 314430 356192 398890
rect 356348 398857 356376 399434
rect 356428 399356 356480 399362
rect 356428 399298 356480 399304
rect 356334 398848 356390 398857
rect 356334 398783 356390 398792
rect 356440 398750 356468 399298
rect 356532 398954 356560 399502
rect 356520 398948 356572 398954
rect 356520 398890 356572 398896
rect 356520 398812 356572 398818
rect 356520 398754 356572 398760
rect 356428 398744 356480 398750
rect 356428 398686 356480 398692
rect 356428 397724 356480 397730
rect 356428 397666 356480 397672
rect 356440 394641 356468 397666
rect 356532 397497 356560 398754
rect 356518 397488 356574 397497
rect 356518 397423 356574 397432
rect 356426 394632 356482 394641
rect 356426 394567 356482 394576
rect 356244 394052 356296 394058
rect 356244 393994 356296 394000
rect 356256 374649 356284 393994
rect 356624 386414 356652 399622
rect 356716 390386 356744 399656
rect 356886 399599 356942 399608
rect 356992 399656 357066 399684
rect 357176 399724 357250 399752
rect 356796 399492 356848 399498
rect 356992 399480 357020 399656
rect 357176 399616 357204 399724
rect 357314 399684 357342 400044
rect 356796 399434 356848 399440
rect 356900 399452 357020 399480
rect 357084 399588 357204 399616
rect 357268 399656 357342 399684
rect 356808 397610 356836 399434
rect 356900 397730 356928 399452
rect 356888 397724 356940 397730
rect 356888 397666 356940 397672
rect 356808 397582 356928 397610
rect 356796 397520 356848 397526
rect 356796 397462 356848 397468
rect 356704 390380 356756 390386
rect 356704 390322 356756 390328
rect 356704 388068 356756 388074
rect 356704 388010 356756 388016
rect 356348 386386 356652 386414
rect 356348 376009 356376 386386
rect 356334 376000 356390 376009
rect 356334 375935 356390 375944
rect 356242 374640 356298 374649
rect 356242 374575 356298 374584
rect 356152 314424 356204 314430
rect 356152 314366 356204 314372
rect 356716 307494 356744 388010
rect 356808 310146 356836 397462
rect 356900 386414 356928 397582
rect 357084 397066 357112 399588
rect 357164 399288 357216 399294
rect 357164 399230 357216 399236
rect 357176 398857 357204 399230
rect 357162 398848 357218 398857
rect 357162 398783 357218 398792
rect 356992 397038 357112 397066
rect 356992 396953 357020 397038
rect 356978 396944 357034 396953
rect 356978 396879 357034 396888
rect 356980 395548 357032 395554
rect 356980 395490 357032 395496
rect 356992 388074 357020 395490
rect 357268 394058 357296 399656
rect 357406 399650 357434 400044
rect 357498 399752 357526 400044
rect 357590 399906 357618 400044
rect 357578 399900 357630 399906
rect 357578 399842 357630 399848
rect 357682 399752 357710 400044
rect 357774 399906 357802 400044
rect 357866 399906 357894 400044
rect 357958 399906 357986 400044
rect 357762 399900 357814 399906
rect 357762 399842 357814 399848
rect 357854 399900 357906 399906
rect 357854 399842 357906 399848
rect 357946 399900 357998 399906
rect 357946 399842 357998 399848
rect 358050 399786 358078 400044
rect 357498 399724 357572 399752
rect 357406 399622 357480 399650
rect 357348 399560 357400 399566
rect 357348 399502 357400 399508
rect 357360 399401 357388 399502
rect 357346 399392 357402 399401
rect 357346 399327 357402 399336
rect 357452 398970 357480 399622
rect 357360 398942 357480 398970
rect 357360 398546 357388 398942
rect 357348 398540 357400 398546
rect 357348 398482 357400 398488
rect 357544 398041 357572 399724
rect 357636 399724 357710 399752
rect 357820 399758 358078 399786
rect 357636 399673 357664 399724
rect 357622 399664 357678 399673
rect 357622 399599 357678 399608
rect 357624 399560 357676 399566
rect 357624 399502 357676 399508
rect 357530 398032 357586 398041
rect 357530 397967 357586 397976
rect 357438 397488 357494 397497
rect 357438 397423 357494 397432
rect 357256 394052 357308 394058
rect 357256 393994 357308 394000
rect 357164 393984 357216 393990
rect 357164 393926 357216 393932
rect 356980 388068 357032 388074
rect 356980 388010 357032 388016
rect 357176 387666 357204 393926
rect 357452 389174 357480 397423
rect 357452 389146 357572 389174
rect 357164 387660 357216 387666
rect 357164 387602 357216 387608
rect 356900 386386 357112 386414
rect 356796 310140 356848 310146
rect 356796 310082 356848 310088
rect 356704 307488 356756 307494
rect 356704 307430 356756 307436
rect 357084 304910 357112 386386
rect 357544 384441 357572 389146
rect 357636 387433 357664 399502
rect 357820 399412 357848 399758
rect 357992 399696 358044 399702
rect 357898 399664 357954 399673
rect 358142 399684 358170 400044
rect 358234 399906 358262 400044
rect 358222 399900 358274 399906
rect 358222 399842 358274 399848
rect 358326 399786 358354 400044
rect 358418 399906 358446 400044
rect 358406 399900 358458 399906
rect 358406 399842 358458 399848
rect 358510 399838 358538 400044
rect 358498 399832 358550 399838
rect 358326 399758 358400 399786
rect 358498 399774 358550 399780
rect 358602 399786 358630 400044
rect 358694 399906 358722 400044
rect 358682 399900 358734 399906
rect 358682 399842 358734 399848
rect 358786 399786 358814 400044
rect 358878 399906 358906 400044
rect 358866 399900 358918 399906
rect 358866 399842 358918 399848
rect 358602 399758 358676 399786
rect 358786 399758 358906 399786
rect 357992 399638 358044 399644
rect 358096 399656 358170 399684
rect 358268 399696 358320 399702
rect 357898 399599 357954 399608
rect 357728 399384 357848 399412
rect 357622 387424 357678 387433
rect 357622 387359 357678 387368
rect 357728 387190 357756 399384
rect 357912 399344 357940 399599
rect 357820 399316 357940 399344
rect 357820 398070 357848 399316
rect 357898 399256 357954 399265
rect 357898 399191 357954 399200
rect 357808 398064 357860 398070
rect 357808 398006 357860 398012
rect 357808 397588 357860 397594
rect 357808 397530 357860 397536
rect 357716 387184 357768 387190
rect 357716 387126 357768 387132
rect 357530 384432 357586 384441
rect 357530 384367 357586 384376
rect 357072 304904 357124 304910
rect 357072 304846 357124 304852
rect 357820 302122 357848 397530
rect 357912 393281 357940 399191
rect 358004 397526 358032 399638
rect 358096 399401 358124 399656
rect 358268 399638 358320 399644
rect 358176 399560 358228 399566
rect 358176 399502 358228 399508
rect 358082 399392 358138 399401
rect 358082 399327 358138 399336
rect 358084 399288 358136 399294
rect 358084 399230 358136 399236
rect 357992 397520 358044 397526
rect 357992 397462 358044 397468
rect 358096 397361 358124 399230
rect 358082 397352 358138 397361
rect 358082 397287 358138 397296
rect 358188 393314 358216 399502
rect 358280 399265 358308 399638
rect 358266 399256 358322 399265
rect 358266 399191 358322 399200
rect 358372 397905 358400 399758
rect 358544 399696 358596 399702
rect 358544 399638 358596 399644
rect 358452 399628 358504 399634
rect 358452 399570 358504 399576
rect 358464 398177 358492 399570
rect 358450 398168 358506 398177
rect 358556 398138 358584 399638
rect 358450 398103 358506 398112
rect 358544 398132 358596 398138
rect 358544 398074 358596 398080
rect 358358 397896 358414 397905
rect 358358 397831 358414 397840
rect 358360 397520 358412 397526
rect 358360 397462 358412 397468
rect 358268 396704 358320 396710
rect 358268 396646 358320 396652
rect 358004 393286 358216 393314
rect 357898 393272 357954 393281
rect 357898 393207 357954 393216
rect 358004 321094 358032 393286
rect 358280 393122 358308 396646
rect 358188 393094 358308 393122
rect 358082 392592 358138 392601
rect 358082 392527 358138 392536
rect 357992 321088 358044 321094
rect 357992 321030 358044 321036
rect 358096 311778 358124 392527
rect 358188 321026 358216 393094
rect 358268 392964 358320 392970
rect 358268 392906 358320 392912
rect 358280 385014 358308 392906
rect 358372 385966 358400 397462
rect 358648 397254 358676 399758
rect 358878 399684 358906 399758
rect 358832 399656 358906 399684
rect 358728 399356 358780 399362
rect 358728 399298 358780 399304
rect 358636 397248 358688 397254
rect 358636 397190 358688 397196
rect 358740 392970 358768 399298
rect 358832 396710 358860 399656
rect 358970 399616 358998 400044
rect 358924 399588 358998 399616
rect 358924 396953 358952 399588
rect 359062 399548 359090 400044
rect 359154 399838 359182 400044
rect 359246 399906 359274 400044
rect 359234 399900 359286 399906
rect 359234 399842 359286 399848
rect 359142 399832 359194 399838
rect 359142 399774 359194 399780
rect 359338 399752 359366 400044
rect 359430 399906 359458 400044
rect 359418 399900 359470 399906
rect 359418 399842 359470 399848
rect 359522 399752 359550 400044
rect 359614 399906 359642 400044
rect 359602 399900 359654 399906
rect 359602 399842 359654 399848
rect 359706 399838 359734 400044
rect 359798 399838 359826 400044
rect 359890 399838 359918 400044
rect 359694 399832 359746 399838
rect 359694 399774 359746 399780
rect 359786 399832 359838 399838
rect 359786 399774 359838 399780
rect 359878 399832 359930 399838
rect 359878 399774 359930 399780
rect 359338 399724 359458 399752
rect 359522 399724 359596 399752
rect 359430 399684 359458 399724
rect 359430 399673 359504 399684
rect 359430 399664 359518 399673
rect 359430 399656 359462 399664
rect 359280 399628 359332 399634
rect 359462 399599 359518 399608
rect 359280 399570 359332 399576
rect 359016 399520 359090 399548
rect 358910 396944 358966 396953
rect 358910 396879 358966 396888
rect 358820 396704 358872 396710
rect 358820 396646 358872 396652
rect 359016 394482 359044 399520
rect 359096 399424 359148 399430
rect 359096 399366 359148 399372
rect 359108 397458 359136 399366
rect 359188 398744 359240 398750
rect 359188 398686 359240 398692
rect 359096 397452 359148 397458
rect 359096 397394 359148 397400
rect 359200 394602 359228 398686
rect 359188 394596 359240 394602
rect 359188 394538 359240 394544
rect 358924 394454 359044 394482
rect 358924 394330 358952 394454
rect 358912 394324 358964 394330
rect 358912 394266 358964 394272
rect 359004 394324 359056 394330
rect 359004 394266 359056 394272
rect 358728 392964 358780 392970
rect 358728 392906 358780 392912
rect 358360 385960 358412 385966
rect 358360 385902 358412 385908
rect 358268 385008 358320 385014
rect 358268 384950 358320 384956
rect 359016 381682 359044 394266
rect 359188 391264 359240 391270
rect 359188 391206 359240 391212
rect 359004 381676 359056 381682
rect 359004 381618 359056 381624
rect 358176 321020 358228 321026
rect 358176 320962 358228 320968
rect 359200 319666 359228 391206
rect 359292 377466 359320 399570
rect 359372 399560 359424 399566
rect 359372 399502 359424 399508
rect 359464 399560 359516 399566
rect 359464 399502 359516 399508
rect 359384 387258 359412 399502
rect 359476 393990 359504 399502
rect 359568 398750 359596 399724
rect 359648 399696 359700 399702
rect 359982 399684 360010 400044
rect 360074 399906 360102 400044
rect 360062 399900 360114 399906
rect 360062 399842 360114 399848
rect 359648 399638 359700 399644
rect 359936 399656 360010 399684
rect 359556 398744 359608 398750
rect 359556 398686 359608 398692
rect 359556 398540 359608 398546
rect 359556 398482 359608 398488
rect 359568 396114 359596 398482
rect 359660 397322 359688 399638
rect 359740 399628 359792 399634
rect 359740 399570 359792 399576
rect 359832 399628 359884 399634
rect 359832 399570 359884 399576
rect 359648 397316 359700 397322
rect 359648 397258 359700 397264
rect 359568 396086 359688 396114
rect 359464 393984 359516 393990
rect 359464 393926 359516 393932
rect 359464 392964 359516 392970
rect 359464 392906 359516 392912
rect 359372 387252 359424 387258
rect 359372 387194 359424 387200
rect 359280 377460 359332 377466
rect 359280 377402 359332 377408
rect 359188 319660 359240 319666
rect 359188 319602 359240 319608
rect 358084 311772 358136 311778
rect 358084 311714 358136 311720
rect 357808 302116 357860 302122
rect 357808 302058 357860 302064
rect 359476 300286 359504 392906
rect 359556 392556 359608 392562
rect 359556 392498 359608 392504
rect 359568 304978 359596 392498
rect 359660 308854 359688 396086
rect 359752 394330 359780 399570
rect 359740 394324 359792 394330
rect 359740 394266 359792 394272
rect 359740 393304 359792 393310
rect 359740 393246 359792 393252
rect 359752 319054 359780 393246
rect 359844 391270 359872 399570
rect 359936 396409 359964 399656
rect 360166 399650 360194 400044
rect 360258 399906 360286 400044
rect 360350 399906 360378 400044
rect 360246 399900 360298 399906
rect 360246 399842 360298 399848
rect 360338 399900 360390 399906
rect 360338 399842 360390 399848
rect 360442 399752 360470 400044
rect 360396 399724 360470 399752
rect 360166 399622 360240 399650
rect 360016 399560 360068 399566
rect 360016 399502 360068 399508
rect 359922 396400 359978 396409
rect 359922 396335 359978 396344
rect 360028 396250 360056 399502
rect 360108 399492 360160 399498
rect 360108 399434 360160 399440
rect 359936 396222 360056 396250
rect 359936 394097 359964 396222
rect 360120 396114 360148 399434
rect 360028 396086 360148 396114
rect 360028 394670 360056 396086
rect 360108 396024 360160 396030
rect 360108 395966 360160 395972
rect 360016 394664 360068 394670
rect 360016 394606 360068 394612
rect 359922 394088 359978 394097
rect 359922 394023 359978 394032
rect 360120 392562 360148 395966
rect 360212 393310 360240 399622
rect 360292 399628 360344 399634
rect 360292 399570 360344 399576
rect 360304 396545 360332 399570
rect 360396 398342 360424 399724
rect 360534 399684 360562 400044
rect 360488 399656 360562 399684
rect 360384 398336 360436 398342
rect 360384 398278 360436 398284
rect 360290 396536 360346 396545
rect 360290 396471 360346 396480
rect 360488 393446 360516 399656
rect 360626 399616 360654 400044
rect 360718 399906 360746 400044
rect 360810 399906 360838 400044
rect 360706 399900 360758 399906
rect 360706 399842 360758 399848
rect 360798 399900 360850 399906
rect 360798 399842 360850 399848
rect 360750 399800 360806 399809
rect 360902 399786 360930 400044
rect 360806 399758 360930 399786
rect 360750 399735 360806 399744
rect 360994 399684 361022 400044
rect 361086 399906 361114 400044
rect 361178 399906 361206 400044
rect 361270 399906 361298 400044
rect 361074 399900 361126 399906
rect 361074 399842 361126 399848
rect 361166 399900 361218 399906
rect 361166 399842 361218 399848
rect 361258 399900 361310 399906
rect 361258 399842 361310 399848
rect 361362 399684 361390 400044
rect 361454 399838 361482 400044
rect 361546 399906 361574 400044
rect 361534 399900 361586 399906
rect 361534 399842 361586 399848
rect 361638 399838 361666 400044
rect 361442 399832 361494 399838
rect 361442 399774 361494 399780
rect 361626 399832 361678 399838
rect 361730 399809 361758 400044
rect 361626 399774 361678 399780
rect 361716 399800 361772 399809
rect 361716 399735 361772 399744
rect 360994 399656 361068 399684
rect 360580 399588 360654 399616
rect 360476 393440 360528 393446
rect 360476 393382 360528 393388
rect 360200 393304 360252 393310
rect 360200 393246 360252 393252
rect 360474 393272 360530 393281
rect 360474 393207 360530 393216
rect 360108 392556 360160 392562
rect 360108 392498 360160 392504
rect 359832 391264 359884 391270
rect 359832 391206 359884 391212
rect 360488 385937 360516 393207
rect 360580 392873 360608 399588
rect 360936 399560 360988 399566
rect 360936 399502 360988 399508
rect 360660 399492 360712 399498
rect 360660 399434 360712 399440
rect 360844 399492 360896 399498
rect 360844 399434 360896 399440
rect 360672 398478 360700 399434
rect 360752 399288 360804 399294
rect 360752 399230 360804 399236
rect 360660 398472 360712 398478
rect 360660 398414 360712 398420
rect 360764 397882 360792 399230
rect 360672 397854 360792 397882
rect 360566 392864 360622 392873
rect 360566 392799 360622 392808
rect 360568 390380 360620 390386
rect 360568 390322 360620 390328
rect 360474 385928 360530 385937
rect 360474 385863 360530 385872
rect 359740 319048 359792 319054
rect 359740 318990 359792 318996
rect 359648 308848 359700 308854
rect 359648 308790 359700 308796
rect 359556 304972 359608 304978
rect 359556 304914 359608 304920
rect 360580 302190 360608 390322
rect 360672 314362 360700 397854
rect 360856 397780 360884 399434
rect 360764 397752 360884 397780
rect 360764 396778 360792 397752
rect 360948 397712 360976 399502
rect 360856 397684 360976 397712
rect 360856 396914 360884 397684
rect 360936 397588 360988 397594
rect 360936 397530 360988 397536
rect 360844 396908 360896 396914
rect 360844 396850 360896 396856
rect 360752 396772 360804 396778
rect 360752 396714 360804 396720
rect 360844 396364 360896 396370
rect 360844 396306 360896 396312
rect 360752 391876 360804 391882
rect 360752 391818 360804 391824
rect 360764 385898 360792 391818
rect 360752 385892 360804 385898
rect 360752 385834 360804 385840
rect 360660 314356 360712 314362
rect 360660 314298 360712 314304
rect 360856 304842 360884 396306
rect 360948 308922 360976 397530
rect 361040 395554 361068 399656
rect 361316 399656 361390 399684
rect 361822 399684 361850 400044
rect 361914 399906 361942 400044
rect 361902 399900 361954 399906
rect 361902 399842 361954 399848
rect 362006 399838 362034 400044
rect 361994 399832 362046 399838
rect 361994 399774 362046 399780
rect 362098 399684 362126 400044
rect 361822 399656 361896 399684
rect 361316 399480 361344 399656
rect 361396 399560 361448 399566
rect 361396 399502 361448 399508
rect 361580 399560 361632 399566
rect 361580 399502 361632 399508
rect 361764 399560 361816 399566
rect 361764 399502 361816 399508
rect 361224 399452 361344 399480
rect 361120 397724 361172 397730
rect 361120 397666 361172 397672
rect 361028 395548 361080 395554
rect 361028 395490 361080 395496
rect 361028 395412 361080 395418
rect 361028 395354 361080 395360
rect 361040 321230 361068 395354
rect 361132 391882 361160 397666
rect 361120 391876 361172 391882
rect 361120 391818 361172 391824
rect 361224 384946 361252 399452
rect 361304 399356 361356 399362
rect 361304 399298 361356 399304
rect 361316 393009 361344 399298
rect 361408 397769 361436 399502
rect 361488 399492 361540 399498
rect 361488 399434 361540 399440
rect 361394 397760 361450 397769
rect 361500 397730 361528 399434
rect 361394 397695 361450 397704
rect 361488 397724 361540 397730
rect 361488 397666 361540 397672
rect 361592 396506 361620 399502
rect 361672 399424 361724 399430
rect 361672 399366 361724 399372
rect 361580 396500 361632 396506
rect 361580 396442 361632 396448
rect 361488 393440 361540 393446
rect 361488 393382 361540 393388
rect 361302 393000 361358 393009
rect 361302 392935 361358 392944
rect 361212 384940 361264 384946
rect 361212 384882 361264 384888
rect 361028 321224 361080 321230
rect 361028 321166 361080 321172
rect 361500 318918 361528 393382
rect 361684 392494 361712 399366
rect 361776 396409 361804 399502
rect 361762 396400 361818 396409
rect 361762 396335 361818 396344
rect 361868 396098 361896 399656
rect 362052 399656 362126 399684
rect 362052 396681 362080 399656
rect 362190 399650 362218 400044
rect 362282 399838 362310 400044
rect 362374 399838 362402 400044
rect 362466 399838 362494 400044
rect 362270 399832 362322 399838
rect 362270 399774 362322 399780
rect 362362 399832 362414 399838
rect 362362 399774 362414 399780
rect 362454 399832 362506 399838
rect 362558 399809 362586 400044
rect 362454 399774 362506 399780
rect 362544 399800 362600 399809
rect 362650 399786 362678 400044
rect 362742 399906 362770 400044
rect 362730 399900 362782 399906
rect 362730 399842 362782 399848
rect 362650 399758 362724 399786
rect 362544 399735 362600 399744
rect 362316 399696 362368 399702
rect 362190 399622 362264 399650
rect 362316 399638 362368 399644
rect 362592 399696 362644 399702
rect 362592 399638 362644 399644
rect 362132 399560 362184 399566
rect 362132 399502 362184 399508
rect 362038 396672 362094 396681
rect 362038 396607 362094 396616
rect 361946 396128 362002 396137
rect 361856 396092 361908 396098
rect 361946 396063 362002 396072
rect 361856 396034 361908 396040
rect 361764 395072 361816 395078
rect 361764 395014 361816 395020
rect 361672 392488 361724 392494
rect 361672 392430 361724 392436
rect 361776 389774 361804 395014
rect 361856 394732 361908 394738
rect 361856 394674 361908 394680
rect 361764 389768 361816 389774
rect 361764 389710 361816 389716
rect 361868 384810 361896 394674
rect 361856 384804 361908 384810
rect 361856 384746 361908 384752
rect 361488 318912 361540 318918
rect 361488 318854 361540 318860
rect 360936 308916 360988 308922
rect 360936 308858 360988 308864
rect 360844 304836 360896 304842
rect 360844 304778 360896 304784
rect 360568 302184 360620 302190
rect 360568 302126 360620 302132
rect 361960 301850 361988 396063
rect 362144 303482 362172 399502
rect 362236 395078 362264 399622
rect 362328 397526 362356 399638
rect 362408 399628 362460 399634
rect 362408 399570 362460 399576
rect 362316 397520 362368 397526
rect 362316 397462 362368 397468
rect 362316 396908 362368 396914
rect 362316 396850 362368 396856
rect 362224 395072 362276 395078
rect 362224 395014 362276 395020
rect 362224 393440 362276 393446
rect 362224 393382 362276 393388
rect 362236 305998 362264 393382
rect 362328 316878 362356 396850
rect 362420 384742 362448 399570
rect 362500 399560 362552 399566
rect 362500 399502 362552 399508
rect 362512 397390 362540 399502
rect 362500 397384 362552 397390
rect 362500 397326 362552 397332
rect 362604 394738 362632 399638
rect 362696 398410 362724 399758
rect 362834 399684 362862 400044
rect 362926 399906 362954 400044
rect 362914 399900 362966 399906
rect 362914 399842 362966 399848
rect 363018 399786 363046 400044
rect 363110 399906 363138 400044
rect 363098 399900 363150 399906
rect 363098 399842 363150 399848
rect 363018 399758 363092 399786
rect 362788 399656 362862 399684
rect 362684 398404 362736 398410
rect 362684 398346 362736 398352
rect 362592 394732 362644 394738
rect 362592 394674 362644 394680
rect 362788 392465 362816 399656
rect 363064 399650 363092 399758
rect 363202 399684 363230 400044
rect 362972 399622 363092 399650
rect 363156 399656 363230 399684
rect 362868 399084 362920 399090
rect 362868 399026 362920 399032
rect 362880 392737 362908 399026
rect 362972 396370 363000 399622
rect 363052 399560 363104 399566
rect 363052 399502 363104 399508
rect 363064 396953 363092 399502
rect 363156 398546 363184 399656
rect 363294 399548 363322 400044
rect 363386 399684 363414 400044
rect 363478 399752 363506 400044
rect 363570 399906 363598 400044
rect 363662 399906 363690 400044
rect 363558 399900 363610 399906
rect 363558 399842 363610 399848
rect 363650 399900 363702 399906
rect 363650 399842 363702 399848
rect 363754 399752 363782 400044
rect 363478 399724 363644 399752
rect 363386 399656 363552 399684
rect 363294 399520 363460 399548
rect 363236 399424 363288 399430
rect 363236 399366 363288 399372
rect 363328 399424 363380 399430
rect 363328 399366 363380 399372
rect 363144 398540 363196 398546
rect 363144 398482 363196 398488
rect 363050 396944 363106 396953
rect 363050 396879 363106 396888
rect 362960 396364 363012 396370
rect 362960 396306 363012 396312
rect 363144 393508 363196 393514
rect 363144 393450 363196 393456
rect 362866 392728 362922 392737
rect 362866 392663 362922 392672
rect 362774 392456 362830 392465
rect 362774 392391 362830 392400
rect 362408 384736 362460 384742
rect 362408 384678 362460 384684
rect 363156 384674 363184 393450
rect 363248 384878 363276 399366
rect 363340 392630 363368 399366
rect 363432 396642 363460 399520
rect 363524 398274 363552 399656
rect 363512 398268 363564 398274
rect 363512 398210 363564 398216
rect 363616 397594 363644 399724
rect 363708 399724 363782 399752
rect 363708 398818 363736 399724
rect 363846 399684 363874 400044
rect 363938 399809 363966 400044
rect 364030 399906 364058 400044
rect 364018 399900 364070 399906
rect 364018 399842 364070 399848
rect 363924 399800 363980 399809
rect 363924 399735 363980 399744
rect 363800 399656 363874 399684
rect 363972 399696 364024 399702
rect 363696 398812 363748 398818
rect 363696 398754 363748 398760
rect 363800 398698 363828 399656
rect 364122 399684 364150 400044
rect 364214 399752 364242 400044
rect 364306 399906 364334 400044
rect 364398 399906 364426 400044
rect 364294 399900 364346 399906
rect 364294 399842 364346 399848
rect 364386 399900 364438 399906
rect 364386 399842 364438 399848
rect 364490 399786 364518 400044
rect 364582 399906 364610 400044
rect 364570 399900 364622 399906
rect 364570 399842 364622 399848
rect 364490 399758 364564 399786
rect 364214 399724 364288 399752
rect 364122 399656 364196 399684
rect 363972 399638 364024 399644
rect 363708 398670 363828 398698
rect 363604 397588 363656 397594
rect 363604 397530 363656 397536
rect 363512 396704 363564 396710
rect 363512 396646 363564 396652
rect 363420 396636 363472 396642
rect 363420 396578 363472 396584
rect 363420 393576 363472 393582
rect 363420 393518 363472 393524
rect 363328 392624 363380 392630
rect 363328 392566 363380 392572
rect 363236 384872 363288 384878
rect 363236 384814 363288 384820
rect 363144 384668 363196 384674
rect 363144 384610 363196 384616
rect 362316 316872 362368 316878
rect 362316 316814 362368 316820
rect 362224 305992 362276 305998
rect 362224 305934 362276 305940
rect 362132 303476 362184 303482
rect 362132 303418 362184 303424
rect 361948 301844 362000 301850
rect 361948 301786 362000 301792
rect 359464 300280 359516 300286
rect 359464 300222 359516 300228
rect 363432 297906 363460 393518
rect 363524 387122 363552 396646
rect 363708 396030 363736 398670
rect 363984 396710 364012 399638
rect 364064 399560 364116 399566
rect 364064 399502 364116 399508
rect 364076 399401 364104 399502
rect 364062 399392 364118 399401
rect 364062 399327 364118 399336
rect 364064 399288 364116 399294
rect 364064 399230 364116 399236
rect 364076 398993 364104 399230
rect 364062 398984 364118 398993
rect 364062 398919 364118 398928
rect 364064 398812 364116 398818
rect 364064 398754 364116 398760
rect 363972 396704 364024 396710
rect 363972 396646 364024 396652
rect 363880 396636 363932 396642
rect 363880 396578 363932 396584
rect 363696 396024 363748 396030
rect 363696 395966 363748 395972
rect 363604 392896 363656 392902
rect 363604 392838 363656 392844
rect 363512 387116 363564 387122
rect 363512 387058 363564 387064
rect 363616 300354 363644 392838
rect 363696 391264 363748 391270
rect 363696 391206 363748 391212
rect 363708 312633 363736 391206
rect 363694 312624 363750 312633
rect 363694 312559 363750 312568
rect 363892 300558 363920 396578
rect 364076 393314 364104 398754
rect 364168 393514 364196 399656
rect 364260 393582 364288 399724
rect 364432 399696 364484 399702
rect 364432 399638 364484 399644
rect 364340 399628 364392 399634
rect 364340 399570 364392 399576
rect 364248 393576 364300 393582
rect 364248 393518 364300 393524
rect 364156 393508 364208 393514
rect 364156 393450 364208 393456
rect 364076 393286 364288 393314
rect 364260 393106 364288 393286
rect 364248 393100 364300 393106
rect 364248 393042 364300 393048
rect 364352 392086 364380 399570
rect 364444 393106 364472 399638
rect 364536 399090 364564 399758
rect 364674 399752 364702 400044
rect 364766 399838 364794 400044
rect 364754 399832 364806 399838
rect 364754 399774 364806 399780
rect 364628 399724 364702 399752
rect 364628 399514 364656 399724
rect 364858 399684 364886 400044
rect 364950 399752 364978 400044
rect 365042 399906 365070 400044
rect 365030 399900 365082 399906
rect 365030 399842 365082 399848
rect 365134 399786 365162 400044
rect 365226 399906 365254 400044
rect 365318 399906 365346 400044
rect 365214 399900 365266 399906
rect 365214 399842 365266 399848
rect 365306 399900 365358 399906
rect 365306 399842 365358 399848
rect 365410 399786 365438 400044
rect 365502 399906 365530 400044
rect 365490 399900 365542 399906
rect 365490 399842 365542 399848
rect 365088 399758 365162 399786
rect 365260 399764 365312 399770
rect 364950 399724 365024 399752
rect 364812 399656 364886 399684
rect 364628 399486 364702 399514
rect 364674 399480 364702 399486
rect 364674 399452 364748 399480
rect 364614 399392 364670 399401
rect 364614 399327 364670 399336
rect 364524 399084 364576 399090
rect 364524 399026 364576 399032
rect 364524 397384 364576 397390
rect 364524 397326 364576 397332
rect 364536 393514 364564 397326
rect 364524 393508 364576 393514
rect 364524 393450 364576 393456
rect 364524 393304 364576 393310
rect 364524 393246 364576 393252
rect 364432 393100 364484 393106
rect 364432 393042 364484 393048
rect 364340 392080 364392 392086
rect 364340 392022 364392 392028
rect 364536 308990 364564 393246
rect 364628 309126 364656 399327
rect 364720 397390 364748 399452
rect 364708 397384 364760 397390
rect 364708 397326 364760 397332
rect 364812 393310 364840 399656
rect 364892 399560 364944 399566
rect 364892 399502 364944 399508
rect 364904 399265 364932 399502
rect 364890 399256 364946 399265
rect 364890 399191 364946 399200
rect 364892 395140 364944 395146
rect 364892 395082 364944 395088
rect 364904 393786 364932 395082
rect 364892 393780 364944 393786
rect 364892 393722 364944 393728
rect 364892 393508 364944 393514
rect 364892 393450 364944 393456
rect 364800 393304 364852 393310
rect 364800 393246 364852 393252
rect 364708 393100 364760 393106
rect 364708 393042 364760 393048
rect 364800 393100 364852 393106
rect 364800 393042 364852 393048
rect 364720 384470 364748 393042
rect 364708 384464 364760 384470
rect 364708 384406 364760 384412
rect 364616 309120 364668 309126
rect 364616 309062 364668 309068
rect 364524 308984 364576 308990
rect 364524 308926 364576 308932
rect 363880 300552 363932 300558
rect 363880 300494 363932 300500
rect 363604 300348 363656 300354
rect 363604 300290 363656 300296
rect 363420 297900 363472 297906
rect 363420 297842 363472 297848
rect 364812 297838 364840 393042
rect 364904 300626 364932 393450
rect 364996 392970 365024 399724
rect 365088 395146 365116 399758
rect 365260 399706 365312 399712
rect 365364 399758 365438 399786
rect 365168 399696 365220 399702
rect 365168 399638 365220 399644
rect 365076 395140 365128 395146
rect 365076 395082 365128 395088
rect 364984 392964 365036 392970
rect 364984 392906 365036 392912
rect 365076 392352 365128 392358
rect 365076 392294 365128 392300
rect 364984 392012 365036 392018
rect 364984 391954 365036 391960
rect 364892 300620 364944 300626
rect 364892 300562 364944 300568
rect 364996 299062 365024 391954
rect 365088 306134 365116 392294
rect 365180 388754 365208 399638
rect 365272 397361 365300 399706
rect 365258 397352 365314 397361
rect 365258 397287 365314 397296
rect 365168 388748 365220 388754
rect 365168 388690 365220 388696
rect 365364 387530 365392 399758
rect 365594 399752 365622 400044
rect 365548 399724 365622 399752
rect 365444 399696 365496 399702
rect 365444 399638 365496 399644
rect 365456 395758 365484 399638
rect 365548 399634 365576 399724
rect 365686 399684 365714 400044
rect 365778 399752 365806 400044
rect 365870 399945 365898 400044
rect 365856 399936 365912 399945
rect 365856 399871 365912 399880
rect 365962 399820 365990 400044
rect 366054 399906 366082 400044
rect 366146 399906 366174 400044
rect 366238 399906 366266 400044
rect 366330 399945 366358 400044
rect 366316 399936 366372 399945
rect 366042 399900 366094 399906
rect 366042 399842 366094 399848
rect 366134 399900 366186 399906
rect 366134 399842 366186 399848
rect 366226 399900 366278 399906
rect 366316 399871 366372 399880
rect 366226 399842 366278 399848
rect 365916 399792 365990 399820
rect 366422 399809 366450 400044
rect 366408 399800 366464 399809
rect 365778 399724 365852 399752
rect 365640 399656 365714 399684
rect 365824 399673 365852 399724
rect 365810 399664 365866 399673
rect 365536 399628 365588 399634
rect 365536 399570 365588 399576
rect 365640 398936 365668 399656
rect 365810 399599 365866 399608
rect 365720 399560 365772 399566
rect 365720 399502 365772 399508
rect 365812 399560 365864 399566
rect 365812 399502 365864 399508
rect 365548 398908 365668 398936
rect 365548 398682 365576 398908
rect 365628 398812 365680 398818
rect 365628 398754 365680 398760
rect 365536 398676 365588 398682
rect 365536 398618 365588 398624
rect 365640 397633 365668 398754
rect 365626 397624 365682 397633
rect 365626 397559 365682 397568
rect 365444 395752 365496 395758
rect 365444 395694 365496 395700
rect 365732 393106 365760 399502
rect 365720 393100 365772 393106
rect 365720 393042 365772 393048
rect 365352 387524 365404 387530
rect 365352 387466 365404 387472
rect 365824 306338 365852 399502
rect 365916 398954 365944 399792
rect 366514 399786 366542 400044
rect 366606 399906 366634 400044
rect 366594 399900 366646 399906
rect 366594 399842 366646 399848
rect 366698 399786 366726 400044
rect 366790 399945 366818 400044
rect 366776 399936 366832 399945
rect 366882 399906 366910 400044
rect 366776 399871 366832 399880
rect 366870 399900 366922 399906
rect 366870 399842 366922 399848
rect 366974 399786 367002 400044
rect 366514 399770 366588 399786
rect 366698 399770 366772 399786
rect 366514 399764 366600 399770
rect 366514 399758 366548 399764
rect 366408 399735 366464 399744
rect 366698 399764 366784 399770
rect 366698 399758 366732 399764
rect 366548 399706 366600 399712
rect 366732 399706 366784 399712
rect 366824 399764 366876 399770
rect 366824 399706 366876 399712
rect 366928 399758 367002 399786
rect 366364 399696 366416 399702
rect 366836 399673 366864 399706
rect 366364 399638 366416 399644
rect 366822 399664 366878 399673
rect 366088 399628 366140 399634
rect 366088 399570 366140 399576
rect 365904 398948 365956 398954
rect 365904 398890 365956 398896
rect 365996 398268 366048 398274
rect 365996 398210 366048 398216
rect 366008 397390 366036 398210
rect 365996 397384 366048 397390
rect 365996 397326 366048 397332
rect 365996 393304 366048 393310
rect 365996 393246 366048 393252
rect 365902 393136 365958 393145
rect 365902 393071 365958 393080
rect 365916 318306 365944 393071
rect 366008 318374 366036 393246
rect 366100 384606 366128 399570
rect 366180 399152 366232 399158
rect 366180 399094 366232 399100
rect 366192 399022 366220 399094
rect 366180 399016 366232 399022
rect 366180 398958 366232 398964
rect 366180 397384 366232 397390
rect 366180 397326 366232 397332
rect 366088 384600 366140 384606
rect 366088 384542 366140 384548
rect 365996 318368 366048 318374
rect 365996 318310 366048 318316
rect 365904 318300 365956 318306
rect 365904 318242 365956 318248
rect 365812 306332 365864 306338
rect 365812 306274 365864 306280
rect 365076 306128 365128 306134
rect 365076 306070 365128 306076
rect 364984 299056 365036 299062
rect 364984 298998 365036 299004
rect 366192 298042 366220 397326
rect 366376 397050 366404 399638
rect 366640 399628 366692 399634
rect 366822 399599 366878 399608
rect 366640 399570 366692 399576
rect 366456 399560 366508 399566
rect 366456 399502 366508 399508
rect 366364 397044 366416 397050
rect 366364 396986 366416 396992
rect 366364 395548 366416 395554
rect 366364 395490 366416 395496
rect 366376 385694 366404 395490
rect 366468 393174 366496 399502
rect 366548 399492 366600 399498
rect 366548 399434 366600 399440
rect 366456 393168 366508 393174
rect 366456 393110 366508 393116
rect 366364 385688 366416 385694
rect 366364 385630 366416 385636
rect 366560 300490 366588 399434
rect 366652 393961 366680 399570
rect 366732 399560 366784 399566
rect 366732 399502 366784 399508
rect 366638 393952 366694 393961
rect 366638 393887 366694 393896
rect 366744 392902 366772 399502
rect 366928 393310 366956 399758
rect 367066 399684 367094 400044
rect 367020 399656 367094 399684
rect 366916 393304 366968 393310
rect 366916 393246 366968 393252
rect 366732 392896 366784 392902
rect 366732 392838 366784 392844
rect 367020 389978 367048 399656
rect 367158 399616 367186 400044
rect 367250 399809 367278 400044
rect 367236 399800 367292 399809
rect 367236 399735 367292 399744
rect 367342 399684 367370 400044
rect 367434 399838 367462 400044
rect 367422 399832 367474 399838
rect 367422 399774 367474 399780
rect 367526 399786 367554 400044
rect 367618 399906 367646 400044
rect 367710 399945 367738 400044
rect 367696 399936 367752 399945
rect 367606 399900 367658 399906
rect 367696 399871 367752 399880
rect 367606 399842 367658 399848
rect 367802 399820 367830 400044
rect 367650 399800 367706 399809
rect 367526 399758 367600 399786
rect 367296 399656 367370 399684
rect 367468 399696 367520 399702
rect 367158 399588 367232 399616
rect 367204 391814 367232 399588
rect 367296 393281 367324 399656
rect 367468 399638 367520 399644
rect 367376 399424 367428 399430
rect 367376 399366 367428 399372
rect 367282 393272 367338 393281
rect 367282 393207 367338 393216
rect 367282 392864 367338 392873
rect 367282 392799 367338 392808
rect 367192 391808 367244 391814
rect 367192 391750 367244 391756
rect 367008 389972 367060 389978
rect 367008 389914 367060 389920
rect 367296 377505 367324 392799
rect 367388 378826 367416 399366
rect 367480 393514 367508 399638
rect 367572 399430 367600 399758
rect 367650 399735 367706 399744
rect 367756 399792 367830 399820
rect 367560 399424 367612 399430
rect 367560 399366 367612 399372
rect 367560 399288 367612 399294
rect 367558 399256 367560 399265
rect 367612 399256 367614 399265
rect 367558 399191 367614 399200
rect 367664 395865 367692 399735
rect 367756 397372 367784 399792
rect 367894 399752 367922 400044
rect 367848 399724 367922 399752
rect 367986 399752 368014 400044
rect 368078 399945 368106 400044
rect 368064 399936 368120 399945
rect 368064 399871 368120 399880
rect 368170 399752 368198 400044
rect 368262 399838 368290 400044
rect 368354 399838 368382 400044
rect 368250 399832 368302 399838
rect 368250 399774 368302 399780
rect 368342 399832 368394 399838
rect 368342 399774 368394 399780
rect 367986 399724 368060 399752
rect 367848 398002 367876 399724
rect 367928 399628 367980 399634
rect 367928 399570 367980 399576
rect 367836 397996 367888 398002
rect 367836 397938 367888 397944
rect 367756 397344 367876 397372
rect 367940 397361 367968 399570
rect 367650 395856 367706 395865
rect 367650 395791 367706 395800
rect 367744 395276 367796 395282
rect 367744 395218 367796 395224
rect 367468 393508 367520 393514
rect 367468 393450 367520 393456
rect 367650 393000 367706 393009
rect 367650 392935 367706 392944
rect 367376 378820 367428 378826
rect 367376 378762 367428 378768
rect 367282 377496 367338 377505
rect 367282 377431 367338 377440
rect 367098 315616 367154 315625
rect 367098 315551 367154 315560
rect 366548 300484 366600 300490
rect 366548 300426 366600 300432
rect 366180 298036 366232 298042
rect 366180 297978 366232 297984
rect 364800 297832 364852 297838
rect 364800 297774 364852 297780
rect 355968 291916 356020 291922
rect 355968 291858 356020 291864
rect 357440 291916 357492 291922
rect 357440 291858 357492 291864
rect 349252 252748 349304 252754
rect 349252 252690 349304 252696
rect 348792 239420 348844 239426
rect 348792 239362 348844 239368
rect 345020 226296 345072 226302
rect 345020 226238 345072 226244
rect 342260 199504 342312 199510
rect 342260 199446 342312 199452
rect 342904 199504 342956 199510
rect 342904 199446 342956 199452
rect 338764 193180 338816 193186
rect 338764 193122 338816 193128
rect 341524 144356 341576 144362
rect 341524 144298 341576 144304
rect 338120 137420 338172 137426
rect 338120 137362 338172 137368
rect 337384 100700 337436 100706
rect 337384 100642 337436 100648
rect 336738 66872 336794 66881
rect 336738 66807 336794 66816
rect 336752 16574 336780 66807
rect 338132 16574 338160 137362
rect 340970 65512 341026 65521
rect 340970 65447 341026 65456
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 332692 3392 332744 3398
rect 332692 3334 332744 3340
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 332612 734 332732 762
rect 332704 480 332732 734
rect 333900 480 333928 3334
rect 335084 3188 335136 3194
rect 335084 3130 335136 3136
rect 335096 480 335124 3130
rect 336292 480 336320 16546
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339868 3664 339920 3670
rect 339868 3606 339920 3612
rect 339880 480 339908 3606
rect 340984 480 341012 65447
rect 341536 3670 341564 144298
rect 342272 16574 342300 199446
rect 345020 148368 345072 148374
rect 345020 148310 345072 148316
rect 343638 115288 343694 115297
rect 343638 115223 343694 115232
rect 343652 16574 343680 115223
rect 345032 16574 345060 148310
rect 347780 104168 347832 104174
rect 347780 104110 347832 104116
rect 347792 16574 347820 104110
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 347792 16546 348096 16574
rect 342168 3868 342220 3874
rect 342168 3810 342220 3816
rect 341524 3664 341576 3670
rect 341524 3606 341576 3612
rect 342180 480 342208 3810
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346952 3596 347004 3602
rect 346952 3538 347004 3544
rect 346964 480 346992 3538
rect 348068 480 348096 16546
rect 349160 3664 349212 3670
rect 349160 3606 349212 3612
rect 349172 1850 349200 3606
rect 349264 3602 349292 252690
rect 353300 245744 353352 245750
rect 353300 245686 353352 245692
rect 351920 135992 351972 135998
rect 351920 135934 351972 135940
rect 351184 134700 351236 134706
rect 351184 134642 351236 134648
rect 350538 64152 350594 64161
rect 350538 64087 350594 64096
rect 350552 6914 350580 64087
rect 351196 16574 351224 134642
rect 351932 16574 351960 135934
rect 353312 16574 353340 245686
rect 355324 155372 355376 155378
rect 355324 155314 355376 155320
rect 354678 62792 354734 62801
rect 354678 62727 354734 62736
rect 354692 16574 354720 62727
rect 351196 16546 351316 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 350552 6886 351224 6914
rect 349252 3596 349304 3602
rect 349252 3538 349304 3544
rect 350448 3596 350500 3602
rect 350448 3538 350500 3544
rect 349172 1822 349292 1850
rect 349264 480 349292 1822
rect 350460 480 350488 3538
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 6886
rect 351288 3602 351316 16546
rect 351276 3596 351328 3602
rect 351276 3538 351328 3544
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 355336 3670 355364 155314
rect 356060 145716 356112 145722
rect 356060 145658 356112 145664
rect 356072 16574 356100 145658
rect 356072 16546 356376 16574
rect 355324 3664 355376 3670
rect 355324 3606 355376 3612
rect 356348 480 356376 16546
rect 357452 3346 357480 291858
rect 360200 259480 360252 259486
rect 360200 259422 360252 259428
rect 358820 127696 358872 127702
rect 358820 127638 358872 127644
rect 357530 40624 357586 40633
rect 357530 40559 357586 40568
rect 357544 3466 357572 40559
rect 358832 16574 358860 127638
rect 360212 16574 360240 259422
rect 364340 254040 364392 254046
rect 364340 253982 364392 253988
rect 361580 184204 361632 184210
rect 361580 184146 361632 184152
rect 361592 16574 361620 184146
rect 363604 140072 363656 140078
rect 363604 140014 363656 140020
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 357532 3460 357584 3466
rect 357532 3402 357584 3408
rect 358728 3460 358780 3466
rect 358728 3402 358780 3408
rect 357452 3318 357572 3346
rect 357544 480 357572 3318
rect 358740 480 358768 3402
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361132 480 361160 16546
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363616 3942 363644 140014
rect 364352 16574 364380 253982
rect 367112 16574 367140 315551
rect 367664 300694 367692 392935
rect 367652 300688 367704 300694
rect 367652 300630 367704 300636
rect 367756 291174 367784 395218
rect 367848 393310 367876 397344
rect 367926 397352 367982 397361
rect 367926 397287 367982 397296
rect 367928 396772 367980 396778
rect 367928 396714 367980 396720
rect 367836 393304 367888 393310
rect 367836 393246 367888 393252
rect 367836 392284 367888 392290
rect 367836 392226 367888 392232
rect 367848 306202 367876 392226
rect 367940 306270 367968 396714
rect 368032 395894 368060 399724
rect 368124 399724 368198 399752
rect 368020 395888 368072 395894
rect 368020 395830 368072 395836
rect 368018 393272 368074 393281
rect 368018 393207 368074 393216
rect 368032 320958 368060 393207
rect 368124 385762 368152 399724
rect 368204 399628 368256 399634
rect 368446 399616 368474 400044
rect 368538 399684 368566 400044
rect 368630 399786 368658 400044
rect 368722 399906 368750 400044
rect 368814 399906 368842 400044
rect 368710 399900 368762 399906
rect 368710 399842 368762 399848
rect 368802 399900 368854 399906
rect 368802 399842 368854 399848
rect 368630 399758 368796 399786
rect 368664 399696 368716 399702
rect 368538 399656 368612 399684
rect 368446 399588 368520 399616
rect 368204 399570 368256 399576
rect 368216 395690 368244 399570
rect 368296 399560 368348 399566
rect 368296 399502 368348 399508
rect 368204 395684 368256 395690
rect 368204 395626 368256 395632
rect 368308 390554 368336 399502
rect 368388 399288 368440 399294
rect 368388 399230 368440 399236
rect 368400 395185 368428 399230
rect 368386 395176 368442 395185
rect 368386 395111 368442 395120
rect 368492 392290 368520 399588
rect 368584 395282 368612 399656
rect 368664 399638 368716 399644
rect 368676 396778 368704 399638
rect 368664 396772 368716 396778
rect 368664 396714 368716 396720
rect 368572 395276 368624 395282
rect 368572 395218 368624 395224
rect 368480 392284 368532 392290
rect 368480 392226 368532 392232
rect 368664 391332 368716 391338
rect 368664 391274 368716 391280
rect 368216 390526 368336 390554
rect 368112 385756 368164 385762
rect 368112 385698 368164 385704
rect 368020 320952 368072 320958
rect 368020 320894 368072 320900
rect 367928 306264 367980 306270
rect 367928 306206 367980 306212
rect 367836 306196 367888 306202
rect 367836 306138 367888 306144
rect 368216 297770 368244 390526
rect 368676 318238 368704 391274
rect 368768 381614 368796 399758
rect 368906 399752 368934 400044
rect 368860 399724 368934 399752
rect 368860 395593 368888 399724
rect 368998 399684 369026 400044
rect 369090 399752 369118 400044
rect 369182 399906 369210 400044
rect 369170 399900 369222 399906
rect 369170 399842 369222 399848
rect 369090 399724 369164 399752
rect 368998 399656 369072 399684
rect 368940 399560 368992 399566
rect 368940 399502 368992 399508
rect 368952 395962 368980 399502
rect 369044 397225 369072 399656
rect 369136 399514 369164 399724
rect 369274 399616 369302 400044
rect 369366 399684 369394 400044
rect 369458 399945 369486 400044
rect 369444 399936 369500 399945
rect 369444 399871 369500 399880
rect 369550 399752 369578 400044
rect 369504 399724 369578 399752
rect 369642 399752 369670 400044
rect 369734 399945 369762 400044
rect 369720 399936 369776 399945
rect 369720 399871 369776 399880
rect 369826 399752 369854 400044
rect 369918 399906 369946 400044
rect 369906 399900 369958 399906
rect 369906 399842 369958 399848
rect 370010 399838 370038 400044
rect 370102 399906 370130 400044
rect 370090 399900 370142 399906
rect 370090 399842 370142 399848
rect 369998 399832 370050 399838
rect 369998 399774 370050 399780
rect 370194 399752 370222 400044
rect 370286 399786 370314 400044
rect 370378 399906 370406 400044
rect 370366 399900 370418 399906
rect 370366 399842 370418 399848
rect 370286 399758 370360 399786
rect 369642 399724 369716 399752
rect 369826 399724 369900 399752
rect 369366 399656 369440 399684
rect 369274 399588 369348 399616
rect 369136 399486 369256 399514
rect 369030 397216 369086 397225
rect 369030 397151 369086 397160
rect 368940 395956 368992 395962
rect 368940 395898 368992 395904
rect 369032 395684 369084 395690
rect 369032 395626 369084 395632
rect 368846 395584 368902 395593
rect 368846 395519 368902 395528
rect 368938 394632 368994 394641
rect 368938 394567 368994 394576
rect 368952 394534 368980 394567
rect 368940 394528 368992 394534
rect 368940 394470 368992 394476
rect 368848 393508 368900 393514
rect 368848 393450 368900 393456
rect 368756 381608 368808 381614
rect 368756 381550 368808 381556
rect 368664 318232 368716 318238
rect 368664 318174 368716 318180
rect 368860 301918 368888 393450
rect 368848 301912 368900 301918
rect 368848 301854 368900 301860
rect 369044 301646 369072 395626
rect 369228 309942 369256 399486
rect 369320 391338 369348 399588
rect 369412 391338 369440 399656
rect 369504 398313 369532 399724
rect 369688 399514 369716 399724
rect 369688 399486 369808 399514
rect 369676 399424 369728 399430
rect 369676 399366 369728 399372
rect 369584 399356 369636 399362
rect 369584 399298 369636 399304
rect 369490 398304 369546 398313
rect 369490 398239 369546 398248
rect 369596 393553 369624 399298
rect 369688 395826 369716 399366
rect 369676 395820 369728 395826
rect 369676 395762 369728 395768
rect 369780 395690 369808 399486
rect 369768 395684 369820 395690
rect 369768 395626 369820 395632
rect 369768 395344 369820 395350
rect 369768 395286 369820 395292
rect 369582 393544 369638 393553
rect 369582 393479 369638 393488
rect 369308 391332 369360 391338
rect 369308 391274 369360 391280
rect 369400 391332 369452 391338
rect 369400 391274 369452 391280
rect 369780 311642 369808 395286
rect 369872 392358 369900 399724
rect 370148 399724 370222 399752
rect 370148 399684 370176 399724
rect 369964 399656 370176 399684
rect 369964 395282 369992 399656
rect 370332 399616 370360 399758
rect 370470 399752 370498 400044
rect 370562 399838 370590 400044
rect 370550 399832 370602 399838
rect 370550 399774 370602 399780
rect 370148 399588 370360 399616
rect 370424 399724 370498 399752
rect 370654 399752 370682 400044
rect 370746 399906 370774 400044
rect 370734 399900 370786 399906
rect 370734 399842 370786 399848
rect 370838 399809 370866 400044
rect 370930 399906 370958 400044
rect 371022 399945 371050 400044
rect 371008 399936 371064 399945
rect 370918 399900 370970 399906
rect 371008 399871 371064 399880
rect 370918 399842 370970 399848
rect 371114 399809 371142 400044
rect 370824 399800 370880 399809
rect 370654 399724 370728 399752
rect 370824 399735 370880 399744
rect 371100 399800 371156 399809
rect 371100 399735 371156 399744
rect 371206 399752 371234 400044
rect 371298 399906 371326 400044
rect 371390 399911 371418 400044
rect 371286 399900 371338 399906
rect 371286 399842 371338 399848
rect 371376 399902 371432 399911
rect 371376 399837 371432 399846
rect 371332 399764 371384 399770
rect 371206 399724 371280 399752
rect 370044 399560 370096 399566
rect 370044 399502 370096 399508
rect 369952 395276 370004 395282
rect 369952 395218 370004 395224
rect 370056 395146 370084 399502
rect 370044 395140 370096 395146
rect 370044 395082 370096 395088
rect 370148 393145 370176 399588
rect 370228 399492 370280 399498
rect 370424 399480 370452 399724
rect 370700 399634 370728 399724
rect 370504 399628 370556 399634
rect 370504 399570 370556 399576
rect 370688 399628 370740 399634
rect 370688 399570 370740 399576
rect 370228 399434 370280 399440
rect 370332 399452 370452 399480
rect 370240 393446 370268 399434
rect 370228 393440 370280 393446
rect 370228 393382 370280 393388
rect 370228 393304 370280 393310
rect 370228 393246 370280 393252
rect 370134 393136 370190 393145
rect 370134 393071 370190 393080
rect 369860 392352 369912 392358
rect 369860 392294 369912 392300
rect 369860 391808 369912 391814
rect 369860 391750 369912 391756
rect 369768 311636 369820 311642
rect 369768 311578 369820 311584
rect 369216 309936 369268 309942
rect 369216 309878 369268 309884
rect 369032 301640 369084 301646
rect 369032 301582 369084 301588
rect 369872 300830 369900 391750
rect 369860 300824 369912 300830
rect 369860 300766 369912 300772
rect 370240 297974 370268 393246
rect 370332 301782 370360 399452
rect 370516 399378 370544 399570
rect 370964 399560 371016 399566
rect 370964 399502 371016 399508
rect 370596 399492 370648 399498
rect 370596 399434 370648 399440
rect 370424 399350 370544 399378
rect 370424 392018 370452 399350
rect 370502 399120 370558 399129
rect 370502 399055 370558 399064
rect 370412 392012 370464 392018
rect 370412 391954 370464 391960
rect 370516 307018 370544 399055
rect 370608 395554 370636 399434
rect 370688 399424 370740 399430
rect 370688 399366 370740 399372
rect 370596 395548 370648 395554
rect 370596 395490 370648 395496
rect 370596 392828 370648 392834
rect 370596 392770 370648 392776
rect 370608 321298 370636 392770
rect 370700 384538 370728 399366
rect 370976 392834 371004 399502
rect 371056 399424 371108 399430
rect 371056 399366 371108 399372
rect 371068 396545 371096 399366
rect 371252 398449 371280 399724
rect 371482 399752 371510 400044
rect 371332 399706 371384 399712
rect 371436 399724 371510 399752
rect 371574 399752 371602 400044
rect 371666 399906 371694 400044
rect 371758 399945 371786 400044
rect 371744 399936 371800 399945
rect 371654 399900 371706 399906
rect 371744 399871 371800 399880
rect 371654 399842 371706 399848
rect 371850 399786 371878 400044
rect 371942 399945 371970 400044
rect 371928 399936 371984 399945
rect 372034 399906 372062 400044
rect 372126 399906 372154 400044
rect 372218 399945 372246 400044
rect 372204 399936 372260 399945
rect 371928 399871 371984 399880
rect 372022 399900 372074 399906
rect 372022 399842 372074 399848
rect 372114 399900 372166 399906
rect 372310 399906 372338 400044
rect 372204 399871 372260 399880
rect 372298 399900 372350 399906
rect 372114 399842 372166 399848
rect 372298 399842 372350 399848
rect 372402 399809 372430 400044
rect 372494 399838 372522 400044
rect 372586 399945 372614 400044
rect 372572 399936 372628 399945
rect 372678 399906 372706 400044
rect 372572 399871 372628 399880
rect 372666 399900 372718 399906
rect 372666 399842 372718 399848
rect 372482 399832 372534 399838
rect 371700 399764 371752 399770
rect 371574 399724 371648 399752
rect 371238 398440 371294 398449
rect 371238 398375 371294 398384
rect 371054 396536 371110 396545
rect 371054 396471 371110 396480
rect 370964 392828 371016 392834
rect 370964 392770 371016 392776
rect 371344 390554 371372 399706
rect 371436 398614 371464 399724
rect 371516 399356 371568 399362
rect 371516 399298 371568 399304
rect 371424 398608 371476 398614
rect 371424 398550 371476 398556
rect 371424 398336 371476 398342
rect 371424 398278 371476 398284
rect 371160 390526 371372 390554
rect 370688 384532 370740 384538
rect 370688 384474 370740 384480
rect 370596 321292 370648 321298
rect 370596 321234 370648 321240
rect 371160 311114 371188 390526
rect 371436 311506 371464 398278
rect 371528 318170 371556 399298
rect 371620 395350 371648 399724
rect 371700 399706 371752 399712
rect 371804 399758 371878 399786
rect 372158 399800 372214 399809
rect 371608 395344 371660 395350
rect 371608 395286 371660 395292
rect 371608 395140 371660 395146
rect 371608 395082 371660 395088
rect 371516 318164 371568 318170
rect 371516 318106 371568 318112
rect 371424 311500 371476 311506
rect 371424 311442 371476 311448
rect 371160 311086 371280 311114
rect 371252 310962 371280 311086
rect 371240 310956 371292 310962
rect 371240 310898 371292 310904
rect 370504 307012 370556 307018
rect 370504 306954 370556 306960
rect 370320 301776 370372 301782
rect 370320 301718 370372 301724
rect 370228 297968 370280 297974
rect 370228 297910 370280 297916
rect 368204 297764 368256 297770
rect 368204 297706 368256 297712
rect 367744 291168 367796 291174
rect 367744 291110 367796 291116
rect 369860 145648 369912 145654
rect 369860 145590 369912 145596
rect 369872 16574 369900 145590
rect 364352 16546 364656 16574
rect 367112 16546 367784 16574
rect 369872 16546 370176 16574
rect 363604 3936 363656 3942
rect 363604 3878 363656 3884
rect 363512 3392 363564 3398
rect 363512 3334 363564 3340
rect 363524 480 363552 3334
rect 364628 480 364656 16546
rect 365810 6488 365866 6497
rect 365810 6423 365866 6432
rect 365824 480 365852 6423
rect 367008 3936 367060 3942
rect 367008 3878 367060 3884
rect 367020 480 367048 3878
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369400 6316 369452 6322
rect 369400 6258 369452 6264
rect 369412 480 369440 6258
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 310898
rect 371332 309052 371384 309058
rect 371332 308994 371384 309000
rect 371344 308446 371372 308994
rect 371332 308440 371384 308446
rect 371332 308382 371384 308388
rect 371620 299470 371648 395082
rect 371712 391474 371740 399706
rect 371804 395350 371832 399758
rect 372158 399735 372214 399744
rect 372388 399800 372444 399809
rect 372770 399786 372798 400044
rect 372862 399906 372890 400044
rect 372954 399945 372982 400044
rect 372940 399936 372996 399945
rect 372850 399900 372902 399906
rect 373046 399906 373074 400044
rect 372940 399871 372996 399880
rect 373034 399900 373086 399906
rect 372850 399842 372902 399848
rect 373034 399842 373086 399848
rect 372482 399774 372534 399780
rect 372388 399735 372444 399744
rect 372724 399758 372798 399786
rect 372172 399684 372200 399735
rect 372344 399696 372396 399702
rect 372172 399656 372292 399684
rect 371976 399560 372028 399566
rect 371976 399502 372028 399508
rect 371988 396914 372016 399502
rect 372264 397798 372292 399656
rect 372344 399638 372396 399644
rect 372436 399696 372488 399702
rect 372436 399638 372488 399644
rect 372252 397792 372304 397798
rect 372252 397734 372304 397740
rect 372250 397624 372306 397633
rect 372250 397559 372306 397568
rect 372068 397452 372120 397458
rect 372068 397394 372120 397400
rect 371976 396908 372028 396914
rect 371976 396850 372028 396856
rect 371792 395344 371844 395350
rect 371792 395286 371844 395292
rect 371884 392624 371936 392630
rect 371884 392566 371936 392572
rect 371700 391468 371752 391474
rect 371700 391410 371752 391416
rect 371700 391332 371752 391338
rect 371700 391274 371752 391280
rect 371712 301986 371740 391274
rect 371896 312390 371924 392566
rect 372080 389174 372108 397394
rect 372160 395344 372212 395350
rect 372160 395286 372212 395292
rect 371988 389146 372108 389174
rect 371988 387326 372016 389146
rect 371976 387320 372028 387326
rect 371976 387262 372028 387268
rect 371884 312384 371936 312390
rect 371884 312326 371936 312332
rect 372172 308446 372200 395286
rect 372160 308440 372212 308446
rect 372160 308382 372212 308388
rect 371700 301980 371752 301986
rect 371700 301922 371752 301928
rect 372264 301714 372292 397559
rect 372356 397225 372384 399638
rect 372448 398342 372476 399638
rect 372528 399628 372580 399634
rect 372528 399570 372580 399576
rect 372436 398336 372488 398342
rect 372436 398278 372488 398284
rect 372436 398200 372488 398206
rect 372436 398142 372488 398148
rect 372342 397216 372398 397225
rect 372342 397151 372398 397160
rect 372448 389745 372476 398142
rect 372540 395690 372568 399570
rect 372724 397372 372752 399758
rect 373138 399752 373166 400044
rect 373230 399906 373258 400044
rect 373218 399900 373270 399906
rect 373218 399842 373270 399848
rect 373322 399786 373350 400044
rect 373414 399809 373442 400044
rect 373506 399838 373534 400044
rect 373598 399838 373626 400044
rect 373690 399838 373718 400044
rect 373782 399838 373810 400044
rect 373874 399838 373902 400044
rect 373966 399911 373994 400044
rect 373952 399902 374008 399911
rect 373494 399832 373546 399838
rect 373092 399724 373166 399752
rect 373276 399758 373350 399786
rect 373400 399800 373456 399809
rect 372804 399696 372856 399702
rect 372986 399664 373042 399673
rect 372804 399638 372856 399644
rect 372632 397344 372752 397372
rect 372528 395684 372580 395690
rect 372528 395626 372580 395632
rect 372632 390658 372660 397344
rect 372712 396228 372764 396234
rect 372712 396170 372764 396176
rect 372620 390652 372672 390658
rect 372620 390594 372672 390600
rect 372434 389736 372490 389745
rect 372434 389671 372490 389680
rect 372620 324964 372672 324970
rect 372620 324906 372672 324912
rect 372632 323746 372660 324906
rect 372620 323740 372672 323746
rect 372620 323682 372672 323688
rect 372252 301708 372304 301714
rect 372252 301650 372304 301656
rect 371608 299464 371660 299470
rect 371608 299406 371660 299412
rect 372724 299266 372752 396170
rect 372816 313138 372844 399638
rect 372908 399622 372986 399650
rect 372908 314974 372936 399622
rect 372986 399599 373042 399608
rect 372986 399528 373042 399537
rect 372986 399463 373042 399472
rect 373000 326398 373028 399463
rect 373092 397361 373120 399724
rect 373078 397352 373134 397361
rect 373078 397287 373134 397296
rect 373276 396234 373304 399758
rect 373494 399774 373546 399780
rect 373586 399832 373638 399838
rect 373586 399774 373638 399780
rect 373678 399832 373730 399838
rect 373678 399774 373730 399780
rect 373770 399832 373822 399838
rect 373770 399774 373822 399780
rect 373862 399832 373914 399838
rect 373952 399837 374008 399846
rect 373862 399774 373914 399780
rect 374058 399786 374086 400044
rect 374150 399911 374178 400044
rect 374136 399902 374192 399911
rect 374242 399906 374270 400044
rect 374136 399837 374192 399846
rect 374230 399900 374282 399906
rect 374230 399842 374282 399848
rect 374058 399758 374224 399786
rect 373400 399735 373456 399744
rect 373908 399696 373960 399702
rect 373354 399664 373410 399673
rect 374090 399664 374146 399673
rect 373908 399638 373960 399644
rect 373354 399599 373410 399608
rect 373540 399628 373592 399634
rect 373264 396228 373316 396234
rect 373264 396170 373316 396176
rect 373172 393168 373224 393174
rect 373172 393110 373224 393116
rect 372988 326392 373040 326398
rect 372988 326334 373040 326340
rect 372896 314968 372948 314974
rect 372896 314910 372948 314916
rect 372804 313132 372856 313138
rect 372804 313074 372856 313080
rect 372712 299260 372764 299266
rect 372712 299202 372764 299208
rect 373184 292534 373212 393110
rect 373368 390554 373396 399599
rect 373540 399570 373592 399576
rect 373724 399628 373776 399634
rect 373724 399570 373776 399576
rect 373448 399560 373500 399566
rect 373448 399502 373500 399508
rect 373460 395457 373488 399502
rect 373446 395448 373502 395457
rect 373446 395383 373502 395392
rect 373552 393961 373580 399570
rect 373632 399492 373684 399498
rect 373632 399434 373684 399440
rect 373538 393952 373594 393961
rect 373538 393887 373594 393896
rect 373644 390554 373672 399434
rect 373736 393174 373764 399570
rect 373816 399560 373868 399566
rect 373816 399502 373868 399508
rect 373828 398410 373856 399502
rect 373816 398404 373868 398410
rect 373816 398346 373868 398352
rect 373724 393168 373776 393174
rect 373724 393110 373776 393116
rect 373920 390969 373948 399638
rect 374012 399622 374090 399650
rect 373906 390960 373962 390969
rect 373906 390895 373962 390904
rect 374012 390590 374040 399622
rect 374090 399599 374146 399608
rect 374092 399492 374144 399498
rect 374092 399434 374144 399440
rect 374104 393825 374132 399434
rect 374196 398002 374224 399758
rect 374334 399752 374362 400044
rect 374426 399906 374454 400044
rect 374414 399900 374466 399906
rect 374414 399842 374466 399848
rect 374518 399752 374546 400044
rect 374610 399838 374638 400044
rect 374702 399906 374730 400044
rect 374690 399900 374742 399906
rect 374690 399842 374742 399848
rect 374794 399838 374822 400044
rect 374598 399832 374650 399838
rect 374598 399774 374650 399780
rect 374782 399832 374834 399838
rect 374886 399809 374914 400044
rect 374782 399774 374834 399780
rect 374872 399800 374928 399809
rect 374334 399724 374408 399752
rect 374276 399628 374328 399634
rect 374276 399570 374328 399576
rect 374288 398886 374316 399570
rect 374380 399072 374408 399724
rect 374472 399724 374546 399752
rect 374872 399735 374928 399744
rect 374472 399566 374500 399724
rect 374828 399628 374880 399634
rect 374656 399588 374828 399616
rect 374460 399560 374512 399566
rect 374460 399502 374512 399508
rect 374460 399424 374512 399430
rect 374460 399366 374512 399372
rect 374472 399265 374500 399366
rect 374458 399256 374514 399265
rect 374458 399191 374514 399200
rect 374380 399044 374500 399072
rect 374276 398880 374328 398886
rect 374276 398822 374328 398828
rect 374184 397996 374236 398002
rect 374184 397938 374236 397944
rect 374368 397792 374420 397798
rect 374368 397734 374420 397740
rect 374276 395344 374328 395350
rect 374276 395286 374328 395292
rect 374184 395208 374236 395214
rect 374184 395150 374236 395156
rect 374090 393816 374146 393825
rect 374090 393751 374146 393760
rect 373276 390526 373396 390554
rect 373460 390526 373672 390554
rect 374000 390584 374052 390590
rect 374000 390526 374052 390532
rect 373276 310078 373304 390526
rect 373460 387462 373488 390526
rect 373906 389192 373962 389201
rect 373906 389127 373962 389136
rect 373448 387456 373500 387462
rect 373448 387398 373500 387404
rect 373920 383761 373948 389127
rect 373906 383752 373962 383761
rect 373906 383687 373962 383696
rect 373906 383616 373962 383625
rect 373906 383551 373962 383560
rect 373920 374105 373948 383551
rect 373906 374096 373962 374105
rect 373906 374031 373962 374040
rect 373906 373960 373962 373969
rect 373906 373895 373962 373904
rect 373920 364449 373948 373895
rect 373906 364440 373962 364449
rect 373906 364375 373962 364384
rect 373906 364304 373962 364313
rect 373906 364239 373962 364248
rect 373920 354793 373948 364239
rect 373906 354784 373962 354793
rect 373906 354719 373962 354728
rect 373906 354648 373962 354657
rect 373906 354583 373962 354592
rect 373920 345137 373948 354583
rect 374196 351121 374224 395150
rect 374288 381546 374316 395286
rect 374276 381540 374328 381546
rect 374276 381482 374328 381488
rect 374182 351112 374238 351121
rect 374182 351047 374238 351056
rect 373906 345128 373962 345137
rect 373906 345063 373962 345072
rect 373906 344992 373962 345001
rect 373906 344927 373962 344936
rect 373920 340785 373948 344927
rect 373906 340776 373962 340785
rect 373906 340711 373962 340720
rect 373906 331256 373962 331265
rect 373906 331191 373962 331200
rect 373920 325825 373948 331191
rect 373906 325816 373962 325825
rect 373906 325751 373962 325760
rect 374092 311636 374144 311642
rect 374092 311578 374144 311584
rect 373264 310072 373316 310078
rect 373264 310014 373316 310020
rect 372620 292528 372672 292534
rect 372620 292470 372672 292476
rect 373172 292528 373224 292534
rect 373172 292470 373224 292476
rect 372632 291854 372660 292470
rect 372620 291848 372672 291854
rect 372620 291790 372672 291796
rect 372896 6248 372948 6254
rect 372896 6190 372948 6196
rect 372908 480 372936 6190
rect 374104 3738 374132 311578
rect 374380 300762 374408 397734
rect 374472 391134 374500 399044
rect 374552 395684 374604 395690
rect 374552 395626 374604 395632
rect 374460 391128 374512 391134
rect 374460 391070 374512 391076
rect 374564 389174 374592 395626
rect 374656 395418 374684 399588
rect 374978 399616 375006 400044
rect 375070 399838 375098 400044
rect 375162 399838 375190 400044
rect 375254 399906 375282 400044
rect 375346 399945 375374 400044
rect 375332 399936 375388 399945
rect 375242 399900 375294 399906
rect 375332 399871 375388 399880
rect 375242 399842 375294 399848
rect 375058 399832 375110 399838
rect 375058 399774 375110 399780
rect 375150 399832 375202 399838
rect 375150 399774 375202 399780
rect 375196 399696 375248 399702
rect 375248 399656 375328 399684
rect 375196 399638 375248 399644
rect 375104 399628 375156 399634
rect 374978 399588 375052 399616
rect 374828 399570 374880 399576
rect 374826 399528 374882 399537
rect 374736 399492 374788 399498
rect 374826 399463 374882 399472
rect 374920 399492 374972 399498
rect 374736 399434 374788 399440
rect 374644 395412 374696 395418
rect 374644 395354 374696 395360
rect 374644 395276 374696 395282
rect 374644 395218 374696 395224
rect 374656 390554 374684 395218
rect 374748 393972 374776 399434
rect 374840 394262 374868 399463
rect 374920 399434 374972 399440
rect 374932 397361 374960 399434
rect 374918 397352 374974 397361
rect 374918 397287 374974 397296
rect 374828 394256 374880 394262
rect 374828 394198 374880 394204
rect 375024 394040 375052 399588
rect 375104 399570 375156 399576
rect 375116 395214 375144 399570
rect 375196 399560 375248 399566
rect 375196 399502 375248 399508
rect 375208 395457 375236 399502
rect 375194 395448 375250 395457
rect 375194 395383 375250 395392
rect 375300 395350 375328 399656
rect 375438 399616 375466 400044
rect 375530 399684 375558 400044
rect 375622 399838 375650 400044
rect 375610 399832 375662 399838
rect 375610 399774 375662 399780
rect 375714 399684 375742 400044
rect 375806 399752 375834 400044
rect 375898 399906 375926 400044
rect 375886 399900 375938 399906
rect 375886 399842 375938 399848
rect 375990 399752 376018 400044
rect 376082 399906 376110 400044
rect 376070 399900 376122 399906
rect 376070 399842 376122 399848
rect 376174 399752 376202 400044
rect 376266 399945 376294 400044
rect 376252 399936 376308 399945
rect 376358 399906 376386 400044
rect 376450 399906 376478 400044
rect 376252 399871 376308 399880
rect 376346 399900 376398 399906
rect 376346 399842 376398 399848
rect 376438 399900 376490 399906
rect 376438 399842 376490 399848
rect 376542 399752 376570 400044
rect 375806 399724 375880 399752
rect 375990 399724 376064 399752
rect 375530 399656 375604 399684
rect 375438 399588 375512 399616
rect 375380 399492 375432 399498
rect 375380 399434 375432 399440
rect 375392 396953 375420 399434
rect 375484 398993 375512 399588
rect 375470 398984 375526 398993
rect 375470 398919 375526 398928
rect 375472 398880 375524 398886
rect 375472 398822 375524 398828
rect 375378 396944 375434 396953
rect 375378 396879 375434 396888
rect 375288 395344 375340 395350
rect 375288 395286 375340 395292
rect 375104 395208 375156 395214
rect 375104 395150 375156 395156
rect 375024 394012 375144 394040
rect 374748 393944 375052 393972
rect 374828 393780 374880 393786
rect 374828 393722 374880 393728
rect 374656 390526 374776 390554
rect 374472 389146 374592 389174
rect 374472 302054 374500 389146
rect 374748 377369 374776 390526
rect 374840 387394 374868 393722
rect 374920 391128 374972 391134
rect 374920 391070 374972 391076
rect 374828 387388 374880 387394
rect 374828 387330 374880 387336
rect 374734 377360 374790 377369
rect 374734 377295 374790 377304
rect 374932 310282 374960 391070
rect 375024 315722 375052 393944
rect 375116 393038 375144 394012
rect 375104 393032 375156 393038
rect 375104 392974 375156 392980
rect 375484 390522 375512 398822
rect 375576 395282 375604 399656
rect 375668 399656 375742 399684
rect 375564 395276 375616 395282
rect 375564 395218 375616 395224
rect 375564 394256 375616 394262
rect 375564 394198 375616 394204
rect 375472 390516 375524 390522
rect 375472 390458 375524 390464
rect 375012 315716 375064 315722
rect 375012 315658 375064 315664
rect 375576 311409 375604 394198
rect 375668 315790 375696 399656
rect 375748 399560 375800 399566
rect 375748 399502 375800 399508
rect 375760 398954 375788 399502
rect 375852 399378 375880 399724
rect 375852 399350 375972 399378
rect 375748 398948 375800 398954
rect 375748 398890 375800 398896
rect 375840 395276 375892 395282
rect 375840 395218 375892 395224
rect 375748 392420 375800 392426
rect 375748 392362 375800 392368
rect 375760 354006 375788 392362
rect 375852 359514 375880 395218
rect 375944 369073 375972 399350
rect 376036 393990 376064 399724
rect 376128 399724 376202 399752
rect 376496 399724 376570 399752
rect 376024 393984 376076 393990
rect 376024 393926 376076 393932
rect 376024 393848 376076 393854
rect 376024 393790 376076 393796
rect 376036 370569 376064 393790
rect 376128 392426 376156 399724
rect 376208 399628 376260 399634
rect 376208 399570 376260 399576
rect 376116 392420 376168 392426
rect 376116 392362 376168 392368
rect 376022 370560 376078 370569
rect 376022 370495 376078 370504
rect 375930 369064 375986 369073
rect 375930 368999 375986 369008
rect 375840 359508 375892 359514
rect 375840 359450 375892 359456
rect 375748 354000 375800 354006
rect 375748 353942 375800 353948
rect 375656 315784 375708 315790
rect 375656 315726 375708 315732
rect 375562 311400 375618 311409
rect 375562 311335 375618 311344
rect 374920 310276 374972 310282
rect 374920 310218 374972 310224
rect 374460 302048 374512 302054
rect 374460 301990 374512 301996
rect 374368 300756 374420 300762
rect 374368 300698 374420 300704
rect 376220 299130 376248 399570
rect 376392 399560 376444 399566
rect 376392 399502 376444 399508
rect 376300 399288 376352 399294
rect 376300 399230 376352 399236
rect 376312 398041 376340 399230
rect 376298 398032 376354 398041
rect 376298 397967 376354 397976
rect 376404 395282 376432 399502
rect 376392 395276 376444 395282
rect 376392 395218 376444 395224
rect 376496 394262 376524 399724
rect 376634 399684 376662 400044
rect 376588 399656 376662 399684
rect 376726 399684 376754 400044
rect 376818 399906 376846 400044
rect 376806 399900 376858 399906
rect 376806 399842 376858 399848
rect 376910 399786 376938 400044
rect 377002 399945 377030 400044
rect 376988 399936 377044 399945
rect 376988 399871 377044 399880
rect 377094 399838 377122 400044
rect 377186 399838 377214 400044
rect 377278 399945 377306 400044
rect 377264 399936 377320 399945
rect 377264 399871 377320 399880
rect 377370 399838 377398 400044
rect 377462 399838 377490 400044
rect 376864 399758 376938 399786
rect 377082 399832 377134 399838
rect 377082 399774 377134 399780
rect 377174 399832 377226 399838
rect 377174 399774 377226 399780
rect 377358 399832 377410 399838
rect 377358 399774 377410 399780
rect 377450 399832 377502 399838
rect 377450 399774 377502 399780
rect 377554 399786 377582 400044
rect 377646 399945 377674 400044
rect 377632 399936 377688 399945
rect 377738 399906 377766 400044
rect 377830 399906 377858 400044
rect 377922 399945 377950 400044
rect 377908 399936 377964 399945
rect 377632 399871 377688 399880
rect 377726 399900 377778 399906
rect 377726 399842 377778 399848
rect 377818 399900 377870 399906
rect 377908 399871 377964 399880
rect 377818 399842 377870 399848
rect 377554 399758 377628 399786
rect 376726 399656 376800 399684
rect 376484 394256 376536 394262
rect 376484 394198 376536 394204
rect 376300 393984 376352 393990
rect 376300 393926 376352 393932
rect 376312 307086 376340 393926
rect 376588 393854 376616 399656
rect 376666 399528 376722 399537
rect 376666 399463 376722 399472
rect 376576 393848 376628 393854
rect 376576 393790 376628 393796
rect 376680 390554 376708 399463
rect 376772 397730 376800 399656
rect 376864 398206 376892 399758
rect 376944 399696 376996 399702
rect 376944 399638 376996 399644
rect 377036 399696 377088 399702
rect 377312 399696 377364 399702
rect 377036 399638 377088 399644
rect 377232 399656 377312 399684
rect 376956 399129 376984 399638
rect 376942 399120 376998 399129
rect 376942 399055 376998 399064
rect 376944 398812 376996 398818
rect 376944 398754 376996 398760
rect 376852 398200 376904 398206
rect 376852 398142 376904 398148
rect 376852 398064 376904 398070
rect 376852 398006 376904 398012
rect 376760 397724 376812 397730
rect 376760 397666 376812 397672
rect 376864 394126 376892 398006
rect 376956 395321 376984 398754
rect 376942 395312 376998 395321
rect 376942 395247 376998 395256
rect 376852 394120 376904 394126
rect 376852 394062 376904 394068
rect 376680 390526 376984 390554
rect 376956 314294 376984 390526
rect 377048 316033 377076 399638
rect 377232 394694 377260 399656
rect 377312 399638 377364 399644
rect 377404 399560 377456 399566
rect 377404 399502 377456 399508
rect 377310 399120 377366 399129
rect 377310 399055 377366 399064
rect 377324 398070 377352 399055
rect 377312 398064 377364 398070
rect 377312 398006 377364 398012
rect 377312 396772 377364 396778
rect 377312 396714 377364 396720
rect 377140 394666 377260 394694
rect 377034 316024 377090 316033
rect 377034 315959 377090 315968
rect 377140 315042 377168 394666
rect 377220 393848 377272 393854
rect 377220 393790 377272 393796
rect 377232 325038 377260 393790
rect 377220 325032 377272 325038
rect 377220 324974 377272 324980
rect 377128 315036 377180 315042
rect 377128 314978 377180 314984
rect 376944 314288 376996 314294
rect 376944 314230 376996 314236
rect 376300 307080 376352 307086
rect 376300 307022 376352 307028
rect 377324 304745 377352 396714
rect 377416 396710 377444 399502
rect 377600 399480 377628 399758
rect 377680 399764 377732 399770
rect 377680 399706 377732 399712
rect 377772 399764 377824 399770
rect 377772 399706 377824 399712
rect 377508 399452 377628 399480
rect 377404 396704 377456 396710
rect 377404 396646 377456 396652
rect 377508 393786 377536 399452
rect 377692 399378 377720 399706
rect 377600 399350 377720 399378
rect 377600 398070 377628 399350
rect 377680 399288 377732 399294
rect 377680 399230 377732 399236
rect 377588 398064 377640 398070
rect 377588 398006 377640 398012
rect 377692 396794 377720 399230
rect 377600 396766 377720 396794
rect 377496 393780 377548 393786
rect 377496 393722 377548 393728
rect 377600 390425 377628 396766
rect 377680 396704 377732 396710
rect 377680 396646 377732 396652
rect 377586 390416 377642 390425
rect 377586 390351 377642 390360
rect 377310 304736 377366 304745
rect 377310 304671 377366 304680
rect 377692 299198 377720 396646
rect 377784 393854 377812 399706
rect 378014 399684 378042 400044
rect 377862 399664 377918 399673
rect 377862 399599 377918 399608
rect 377968 399656 378042 399684
rect 378106 399684 378134 400044
rect 378198 399906 378226 400044
rect 378290 399906 378318 400044
rect 378382 399945 378410 400044
rect 378368 399936 378424 399945
rect 378186 399900 378238 399906
rect 378186 399842 378238 399848
rect 378278 399900 378330 399906
rect 378368 399871 378424 399880
rect 378278 399842 378330 399848
rect 378474 399752 378502 400044
rect 378428 399724 378502 399752
rect 378106 399656 378180 399684
rect 377876 396982 377904 399599
rect 377864 396976 377916 396982
rect 377864 396918 377916 396924
rect 377864 396840 377916 396846
rect 377864 396782 377916 396788
rect 377772 393848 377824 393854
rect 377772 393790 377824 393796
rect 377876 389174 377904 396782
rect 377784 389146 377904 389174
rect 377784 323649 377812 389146
rect 377770 323640 377826 323649
rect 377770 323575 377826 323584
rect 377968 300422 377996 399656
rect 378046 396808 378102 396817
rect 378046 396743 378102 396752
rect 378060 393258 378088 396743
rect 378152 395486 378180 399656
rect 378230 399528 378286 399537
rect 378230 399463 378286 399472
rect 378140 395480 378192 395486
rect 378140 395422 378192 395428
rect 378244 395146 378272 399463
rect 378322 395176 378378 395185
rect 378232 395140 378284 395146
rect 378322 395111 378378 395120
rect 378232 395082 378284 395088
rect 378138 393544 378194 393553
rect 378138 393479 378194 393488
rect 378152 393378 378180 393479
rect 378140 393372 378192 393378
rect 378140 393314 378192 393320
rect 378060 393230 378180 393258
rect 378152 390114 378180 393230
rect 378140 390108 378192 390114
rect 378140 390050 378192 390056
rect 378138 389328 378194 389337
rect 378138 389263 378194 389272
rect 378152 389230 378180 389263
rect 378140 389224 378192 389230
rect 378140 389166 378192 389172
rect 378046 321736 378102 321745
rect 378046 321671 378102 321680
rect 378060 321638 378088 321671
rect 378048 321632 378100 321638
rect 378048 321574 378100 321580
rect 377956 300416 378008 300422
rect 377956 300358 378008 300364
rect 377680 299192 377732 299198
rect 377680 299134 377732 299140
rect 376208 299124 376260 299130
rect 376208 299066 376260 299072
rect 376022 151192 376078 151201
rect 376022 151127 376078 151136
rect 376036 3738 376064 151127
rect 376760 124908 376812 124914
rect 376760 124850 376812 124856
rect 376772 16574 376800 124850
rect 376772 16546 377720 16574
rect 376482 6352 376538 6361
rect 376482 6287 376538 6296
rect 374092 3732 374144 3738
rect 374092 3674 374144 3680
rect 375288 3732 375340 3738
rect 375288 3674 375340 3680
rect 376024 3732 376076 3738
rect 376024 3674 376076 3680
rect 374092 3596 374144 3602
rect 374092 3538 374144 3544
rect 374104 480 374132 3538
rect 375300 480 375328 3674
rect 376496 480 376524 6287
rect 377692 480 377720 16546
rect 378060 3602 378088 321574
rect 378336 316606 378364 395111
rect 378428 321638 378456 399724
rect 378566 399684 378594 400044
rect 378520 399656 378594 399684
rect 378658 399684 378686 400044
rect 378750 399752 378778 400044
rect 378842 399945 378870 400044
rect 378828 399936 378884 399945
rect 378934 399906 378962 400044
rect 378828 399871 378884 399880
rect 378922 399900 378974 399906
rect 378922 399842 378974 399848
rect 379026 399752 379054 400044
rect 379118 399906 379146 400044
rect 379106 399900 379158 399906
rect 379106 399842 379158 399848
rect 378750 399724 378916 399752
rect 379026 399724 379100 399752
rect 378658 399656 378824 399684
rect 378520 396914 378548 399656
rect 378600 399560 378652 399566
rect 378598 399528 378600 399537
rect 378652 399528 378654 399537
rect 378598 399463 378654 399472
rect 378600 399424 378652 399430
rect 378600 399366 378652 399372
rect 378508 396908 378560 396914
rect 378508 396850 378560 396856
rect 378612 396692 378640 399366
rect 378692 399356 378744 399362
rect 378692 399298 378744 399304
rect 378520 396664 378640 396692
rect 378520 325106 378548 396664
rect 378704 393836 378732 399298
rect 378796 398274 378824 399656
rect 378784 398268 378836 398274
rect 378784 398210 378836 398216
rect 378784 398064 378836 398070
rect 378784 398006 378836 398012
rect 378612 393808 378732 393836
rect 378612 326466 378640 393808
rect 378796 393314 378824 398006
rect 378888 393650 378916 399724
rect 378966 399664 379022 399673
rect 378966 399599 379022 399608
rect 378980 394466 379008 399599
rect 379072 398818 379100 399724
rect 379210 399684 379238 400044
rect 379302 399945 379330 400044
rect 379288 399936 379344 399945
rect 379394 399906 379422 400044
rect 379486 399945 379514 400044
rect 379472 399936 379528 399945
rect 379288 399871 379344 399880
rect 379382 399900 379434 399906
rect 379472 399871 379528 399880
rect 379382 399842 379434 399848
rect 379578 399786 379606 400044
rect 379670 399911 379698 400044
rect 379656 399902 379712 399911
rect 379762 399906 379790 400044
rect 379656 399837 379712 399846
rect 379750 399900 379802 399906
rect 379750 399842 379802 399848
rect 379336 399764 379388 399770
rect 379336 399706 379388 399712
rect 379532 399758 379606 399786
rect 379704 399764 379756 399770
rect 379210 399656 379284 399684
rect 379152 399560 379204 399566
rect 379152 399502 379204 399508
rect 379060 398812 379112 398818
rect 379060 398754 379112 398760
rect 378968 394460 379020 394466
rect 378968 394402 379020 394408
rect 378876 393644 378928 393650
rect 378876 393586 378928 393592
rect 378704 393286 378824 393314
rect 378600 326460 378652 326466
rect 378600 326402 378652 326408
rect 378508 325100 378560 325106
rect 378508 325042 378560 325048
rect 378416 321632 378468 321638
rect 378416 321574 378468 321580
rect 378324 316600 378376 316606
rect 378324 316542 378376 316548
rect 378140 308440 378192 308446
rect 378140 308382 378192 308388
rect 378152 16574 378180 308382
rect 378704 299402 378732 393286
rect 379164 314498 379192 399502
rect 379256 399362 379284 399656
rect 379244 399356 379296 399362
rect 379244 399298 379296 399304
rect 379242 399256 379298 399265
rect 379242 399191 379298 399200
rect 379256 399158 379284 399191
rect 379244 399152 379296 399158
rect 379244 399094 379296 399100
rect 379348 396681 379376 399706
rect 379428 399696 379480 399702
rect 379428 399638 379480 399644
rect 379334 396672 379390 396681
rect 379334 396607 379390 396616
rect 379244 393644 379296 393650
rect 379244 393586 379296 393592
rect 379152 314492 379204 314498
rect 379152 314434 379204 314440
rect 379256 313954 379284 393586
rect 379440 393314 379468 399638
rect 379532 396030 379560 399758
rect 379854 399752 379882 400044
rect 379946 399945 379974 400044
rect 379932 399936 379988 399945
rect 379932 399871 379988 399880
rect 380038 399786 380066 400044
rect 380130 399809 380158 400044
rect 380222 399945 380250 400044
rect 380208 399936 380264 399945
rect 380314 399906 380342 400044
rect 380208 399871 380264 399880
rect 380302 399900 380354 399906
rect 380302 399842 380354 399848
rect 379992 399770 380066 399786
rect 379704 399706 379756 399712
rect 379808 399724 379882 399752
rect 379980 399764 380066 399770
rect 379612 399696 379664 399702
rect 379612 399638 379664 399644
rect 379624 399226 379652 399638
rect 379612 399220 379664 399226
rect 379612 399162 379664 399168
rect 379716 396846 379744 399706
rect 379808 399566 379836 399724
rect 380032 399758 380066 399764
rect 380116 399800 380172 399809
rect 380406 399752 380434 400044
rect 380498 399838 380526 400044
rect 380486 399832 380538 399838
rect 380486 399774 380538 399780
rect 380590 399786 380618 400044
rect 380682 399906 380710 400044
rect 380670 399900 380722 399906
rect 380670 399842 380722 399848
rect 380774 399786 380802 400044
rect 380590 399758 380664 399786
rect 380116 399735 380172 399744
rect 379980 399706 380032 399712
rect 380360 399724 380434 399752
rect 379978 399664 380034 399673
rect 379978 399599 380034 399608
rect 379796 399560 379848 399566
rect 379796 399502 379848 399508
rect 379992 399242 380020 399599
rect 380162 399528 380218 399537
rect 380162 399463 380218 399472
rect 380256 399492 380308 399498
rect 379900 399214 380020 399242
rect 379704 396840 379756 396846
rect 379704 396782 379756 396788
rect 379702 396672 379758 396681
rect 379702 396607 379758 396616
rect 379520 396024 379572 396030
rect 379520 395966 379572 395972
rect 379348 393286 379468 393314
rect 379348 390182 379376 393286
rect 379336 390176 379388 390182
rect 379336 390118 379388 390124
rect 379244 313948 379296 313954
rect 379244 313890 379296 313896
rect 379256 313818 379284 313890
rect 379244 313812 379296 313818
rect 379244 313754 379296 313760
rect 379716 313750 379744 396607
rect 379796 396024 379848 396030
rect 379796 395966 379848 395972
rect 379808 314129 379836 395966
rect 379900 332654 379928 399214
rect 379980 395480 380032 395486
rect 379980 395422 380032 395428
rect 379992 384402 380020 395422
rect 380072 394256 380124 394262
rect 380072 394198 380124 394204
rect 379980 384396 380032 384402
rect 379980 384338 380032 384344
rect 379888 332648 379940 332654
rect 379888 332590 379940 332596
rect 379900 331906 379928 332590
rect 379888 331900 379940 331906
rect 379888 331842 379940 331848
rect 379794 314120 379850 314129
rect 379794 314055 379850 314064
rect 379704 313744 379756 313750
rect 379704 313686 379756 313692
rect 380084 303346 380112 394198
rect 380176 390046 380204 399463
rect 380256 399434 380308 399440
rect 380268 395729 380296 399434
rect 380254 395720 380310 395729
rect 380254 395655 380310 395664
rect 380360 394262 380388 399724
rect 380532 399696 380584 399702
rect 380532 399638 380584 399644
rect 380440 399628 380492 399634
rect 380440 399570 380492 399576
rect 380348 394256 380400 394262
rect 380348 394198 380400 394204
rect 380452 393314 380480 399570
rect 380544 395321 380572 399638
rect 380636 397186 380664 399758
rect 380728 399758 380802 399786
rect 380728 397905 380756 399758
rect 380866 399684 380894 400044
rect 380958 399786 380986 400044
rect 381050 399945 381078 400044
rect 381036 399936 381092 399945
rect 381036 399871 381092 399880
rect 380958 399758 381032 399786
rect 380820 399656 380894 399684
rect 380820 399265 380848 399656
rect 380900 399560 380952 399566
rect 380900 399502 380952 399508
rect 380806 399256 380862 399265
rect 380806 399191 380862 399200
rect 380714 397896 380770 397905
rect 380714 397831 380770 397840
rect 380624 397180 380676 397186
rect 380624 397122 380676 397128
rect 380530 395312 380586 395321
rect 380530 395247 380586 395256
rect 380912 394694 380940 399502
rect 381004 398546 381032 399758
rect 381142 399752 381170 400044
rect 381234 399906 381262 400044
rect 381222 399900 381274 399906
rect 381222 399842 381274 399848
rect 381326 399752 381354 400044
rect 381096 399724 381170 399752
rect 381280 399724 381354 399752
rect 381418 399752 381446 400044
rect 381510 399906 381538 400044
rect 381602 399906 381630 400044
rect 381694 399945 381722 400044
rect 381680 399936 381736 399945
rect 381498 399900 381550 399906
rect 381498 399842 381550 399848
rect 381590 399900 381642 399906
rect 381680 399871 381736 399880
rect 381590 399842 381642 399848
rect 381786 399786 381814 400044
rect 381740 399758 381814 399786
rect 381418 399724 381492 399752
rect 381096 398750 381124 399724
rect 381174 399664 381230 399673
rect 381174 399599 381230 399608
rect 381188 398954 381216 399599
rect 381176 398948 381228 398954
rect 381176 398890 381228 398896
rect 381084 398744 381136 398750
rect 381084 398686 381136 398692
rect 380992 398540 381044 398546
rect 380992 398482 381044 398488
rect 381280 397798 381308 399724
rect 381360 399628 381412 399634
rect 381360 399570 381412 399576
rect 381268 397792 381320 397798
rect 381268 397734 381320 397740
rect 380992 397180 381044 397186
rect 380992 397122 381044 397128
rect 380360 393286 380480 393314
rect 380820 394666 380940 394694
rect 380164 390040 380216 390046
rect 380164 389982 380216 389988
rect 380164 334008 380216 334014
rect 380164 333950 380216 333956
rect 380176 303414 380204 333950
rect 380164 303408 380216 303414
rect 380164 303350 380216 303356
rect 380072 303340 380124 303346
rect 380072 303282 380124 303288
rect 380360 303278 380388 393286
rect 380820 334014 380848 394666
rect 381004 393314 381032 397122
rect 381084 396976 381136 396982
rect 381084 396918 381136 396924
rect 380912 393286 381032 393314
rect 380808 334008 380860 334014
rect 380808 333950 380860 333956
rect 380912 310321 380940 393286
rect 381096 391406 381124 396918
rect 381268 396908 381320 396914
rect 381268 396850 381320 396856
rect 381174 396536 381230 396545
rect 381174 396471 381230 396480
rect 381084 391400 381136 391406
rect 381084 391342 381136 391348
rect 381188 310350 381216 396471
rect 381280 318102 381308 396850
rect 381268 318096 381320 318102
rect 381268 318038 381320 318044
rect 381372 312458 381400 399570
rect 381464 396778 381492 399724
rect 381544 399560 381596 399566
rect 381544 399502 381596 399508
rect 381556 397934 381584 399502
rect 381636 399152 381688 399158
rect 381636 399094 381688 399100
rect 381544 397928 381596 397934
rect 381544 397870 381596 397876
rect 381544 397792 381596 397798
rect 381544 397734 381596 397740
rect 381452 396772 381504 396778
rect 381452 396714 381504 396720
rect 381452 395956 381504 395962
rect 381452 395898 381504 395904
rect 381464 388550 381492 395898
rect 381556 394233 381584 397734
rect 381648 395622 381676 399094
rect 381636 395616 381688 395622
rect 381636 395558 381688 395564
rect 381542 394224 381598 394233
rect 381542 394159 381598 394168
rect 381740 392766 381768 399758
rect 381878 399684 381906 400044
rect 381970 399906 381998 400044
rect 381958 399900 382010 399906
rect 381958 399842 382010 399848
rect 382062 399786 382090 400044
rect 381832 399656 381906 399684
rect 382016 399758 382090 399786
rect 381832 397769 381860 399656
rect 381912 399560 381964 399566
rect 381912 399502 381964 399508
rect 381924 399158 381952 399502
rect 381912 399152 381964 399158
rect 381912 399094 381964 399100
rect 381912 397928 381964 397934
rect 381912 397870 381964 397876
rect 381818 397760 381874 397769
rect 381818 397695 381874 397704
rect 381728 392760 381780 392766
rect 381728 392702 381780 392708
rect 381452 388544 381504 388550
rect 381452 388486 381504 388492
rect 381924 315761 381952 397870
rect 382016 395962 382044 399758
rect 382154 399684 382182 400044
rect 382246 399906 382274 400044
rect 382234 399900 382286 399906
rect 382234 399842 382286 399848
rect 382338 399786 382366 400044
rect 382108 399656 382182 399684
rect 382292 399758 382366 399786
rect 382108 397633 382136 399656
rect 382188 398948 382240 398954
rect 382188 398890 382240 398896
rect 382094 397624 382150 397633
rect 382094 397559 382150 397568
rect 382200 397338 382228 398890
rect 382292 397497 382320 399758
rect 382430 399684 382458 400044
rect 382522 399786 382550 400044
rect 382614 399906 382642 400044
rect 382706 399945 382734 400044
rect 382692 399936 382748 399945
rect 382602 399900 382654 399906
rect 382798 399906 382826 400044
rect 382692 399871 382748 399880
rect 382786 399900 382838 399906
rect 382602 399842 382654 399848
rect 382786 399842 382838 399848
rect 382522 399758 382596 399786
rect 382430 399656 382504 399684
rect 382372 399560 382424 399566
rect 382372 399502 382424 399508
rect 382384 398614 382412 399502
rect 382476 398954 382504 399656
rect 382464 398948 382516 398954
rect 382464 398890 382516 398896
rect 382568 398682 382596 399758
rect 382648 399764 382700 399770
rect 382890 399752 382918 400044
rect 382982 399809 383010 400044
rect 382648 399706 382700 399712
rect 382752 399724 382918 399752
rect 382968 399800 383024 399809
rect 382968 399735 383024 399744
rect 382556 398676 382608 398682
rect 382556 398618 382608 398624
rect 382372 398608 382424 398614
rect 382372 398550 382424 398556
rect 382278 397488 382334 397497
rect 382278 397423 382334 397432
rect 382372 397384 382424 397390
rect 382200 397310 382320 397338
rect 382372 397326 382424 397332
rect 382462 397352 382518 397361
rect 382004 395956 382056 395962
rect 382004 395898 382056 395904
rect 382292 394398 382320 397310
rect 382280 394392 382332 394398
rect 382280 394334 382332 394340
rect 382384 392630 382412 397326
rect 382462 397287 382518 397296
rect 382372 392624 382424 392630
rect 382372 392566 382424 392572
rect 381910 315752 381966 315761
rect 381910 315687 381966 315696
rect 381360 312452 381412 312458
rect 381360 312394 381412 312400
rect 382476 311137 382504 397287
rect 382660 397186 382688 399706
rect 382752 397390 382780 399724
rect 383074 399616 383102 400044
rect 383166 399809 383194 400044
rect 383152 399800 383208 399809
rect 383152 399735 383208 399744
rect 383258 399650 383286 400044
rect 383350 399786 383378 400044
rect 383442 399906 383470 400044
rect 383430 399900 383482 399906
rect 383430 399842 383482 399848
rect 383534 399786 383562 400044
rect 383350 399758 383424 399786
rect 382936 399588 383102 399616
rect 383212 399622 383286 399650
rect 382830 399528 382886 399537
rect 382830 399463 382886 399472
rect 382740 397384 382792 397390
rect 382740 397326 382792 397332
rect 382844 397202 382872 399463
rect 382936 398478 382964 399588
rect 383106 399528 383162 399537
rect 383106 399463 383162 399472
rect 383016 398880 383068 398886
rect 383016 398822 383068 398828
rect 382924 398472 382976 398478
rect 382924 398414 382976 398420
rect 382924 397996 382976 398002
rect 382924 397938 382976 397944
rect 382648 397180 382700 397186
rect 382648 397122 382700 397128
rect 382752 397174 382872 397202
rect 382752 397066 382780 397174
rect 382568 397038 382780 397066
rect 382568 312769 382596 397038
rect 382648 396568 382700 396574
rect 382648 396510 382700 396516
rect 382660 363662 382688 396510
rect 382936 393314 382964 397938
rect 382752 393286 382964 393314
rect 382648 363656 382700 363662
rect 382648 363598 382700 363604
rect 382752 315110 382780 393286
rect 382740 315104 382792 315110
rect 382740 315046 382792 315052
rect 382554 312760 382610 312769
rect 382554 312695 382610 312704
rect 382462 311128 382518 311137
rect 382462 311063 382518 311072
rect 381176 310344 381228 310350
rect 380898 310312 380954 310321
rect 381176 310286 381228 310292
rect 380898 310247 380954 310256
rect 380348 303272 380400 303278
rect 383028 303249 383056 398822
rect 383120 391270 383148 399463
rect 383108 391264 383160 391270
rect 383108 391206 383160 391212
rect 383212 308689 383240 399622
rect 383292 399560 383344 399566
rect 383292 399502 383344 399508
rect 383304 397118 383332 399502
rect 383292 397112 383344 397118
rect 383292 397054 383344 397060
rect 383396 396574 383424 399758
rect 383488 399758 383562 399786
rect 383626 399786 383654 400044
rect 383718 399906 383746 400044
rect 383810 399906 383838 400044
rect 383706 399900 383758 399906
rect 383706 399842 383758 399848
rect 383798 399900 383850 399906
rect 383798 399842 383850 399848
rect 383902 399786 383930 400044
rect 383994 399809 384022 400044
rect 383626 399758 383700 399786
rect 383488 397633 383516 399758
rect 383568 399696 383620 399702
rect 383568 399638 383620 399644
rect 383580 398886 383608 399638
rect 383568 398880 383620 398886
rect 383568 398822 383620 398828
rect 383474 397624 383530 397633
rect 383474 397559 383530 397568
rect 383672 396658 383700 399758
rect 383764 399758 383930 399786
rect 383980 399800 384036 399809
rect 383764 397254 383792 399758
rect 383980 399735 384036 399744
rect 383936 399696 383988 399702
rect 383842 399664 383898 399673
rect 384086 399684 384114 400044
rect 384178 399906 384206 400044
rect 384270 399906 384298 400044
rect 384362 399945 384390 400044
rect 384348 399936 384404 399945
rect 384166 399900 384218 399906
rect 384166 399842 384218 399848
rect 384258 399900 384310 399906
rect 384454 399906 384482 400044
rect 384348 399871 384404 399880
rect 384442 399900 384494 399906
rect 384258 399842 384310 399848
rect 384442 399842 384494 399848
rect 383936 399638 383988 399644
rect 384040 399656 384114 399684
rect 384304 399696 384356 399702
rect 383842 399599 383898 399608
rect 383752 397248 383804 397254
rect 383752 397190 383804 397196
rect 383672 396630 383792 396658
rect 383384 396568 383436 396574
rect 383384 396510 383436 396516
rect 383660 395684 383712 395690
rect 383660 395626 383712 395632
rect 383672 388686 383700 395626
rect 383660 388680 383712 388686
rect 383660 388622 383712 388628
rect 383764 310214 383792 396630
rect 383752 310208 383804 310214
rect 383856 310185 383884 399599
rect 383948 396710 383976 399638
rect 383936 396704 383988 396710
rect 383936 396646 383988 396652
rect 383936 396500 383988 396506
rect 383936 396442 383988 396448
rect 383948 320929 383976 396442
rect 384040 322930 384068 399656
rect 384546 399650 384574 400044
rect 384638 399843 384666 400044
rect 384624 399834 384680 399843
rect 384624 399769 384680 399778
rect 384730 399770 384758 400044
rect 384718 399764 384770 399770
rect 384718 399706 384770 399712
rect 384304 399638 384356 399644
rect 384316 397338 384344 399638
rect 384224 397310 384344 397338
rect 384408 399622 384574 399650
rect 384670 399664 384726 399673
rect 384120 396704 384172 396710
rect 384120 396646 384172 396652
rect 384132 323610 384160 396646
rect 384224 329118 384252 397310
rect 384304 397180 384356 397186
rect 384304 397122 384356 397128
rect 384316 367810 384344 397122
rect 384408 395690 384436 399622
rect 384670 399599 384726 399608
rect 384822 399616 384850 400044
rect 384914 399945 384942 400044
rect 384900 399936 384956 399945
rect 384900 399871 384956 399880
rect 385006 399786 385034 400044
rect 385098 399838 385126 400044
rect 385190 399945 385218 400044
rect 385176 399936 385232 399945
rect 385176 399871 385232 399880
rect 384960 399758 385034 399786
rect 385086 399832 385138 399838
rect 385086 399774 385138 399780
rect 384580 399560 384632 399566
rect 384580 399502 384632 399508
rect 384488 398404 384540 398410
rect 384488 398346 384540 398352
rect 384396 395684 384448 395690
rect 384396 395626 384448 395632
rect 384304 367804 384356 367810
rect 384304 367746 384356 367752
rect 384212 329112 384264 329118
rect 384212 329054 384264 329060
rect 384500 324970 384528 398346
rect 384592 397186 384620 399502
rect 384580 397180 384632 397186
rect 384580 397122 384632 397128
rect 384684 396506 384712 399599
rect 384822 399588 384896 399616
rect 384764 399492 384816 399498
rect 384764 399434 384816 399440
rect 384776 398177 384804 399434
rect 384762 398168 384818 398177
rect 384762 398103 384818 398112
rect 384672 396500 384724 396506
rect 384672 396442 384724 396448
rect 384488 324964 384540 324970
rect 384488 324906 384540 324912
rect 384120 323604 384172 323610
rect 384120 323546 384172 323552
rect 384028 322924 384080 322930
rect 384028 322866 384080 322872
rect 383934 320920 383990 320929
rect 383934 320855 383990 320864
rect 383752 310150 383804 310156
rect 383842 310176 383898 310185
rect 383842 310111 383898 310120
rect 384868 308961 384896 399588
rect 384960 394694 384988 399758
rect 385282 399752 385310 400044
rect 385374 399945 385402 400044
rect 385360 399936 385416 399945
rect 385360 399871 385416 399880
rect 385466 399752 385494 400044
rect 385558 399906 385586 400044
rect 385546 399900 385598 399906
rect 385546 399842 385598 399848
rect 385650 399838 385678 400044
rect 385742 399843 385770 400044
rect 385638 399832 385690 399838
rect 385638 399774 385690 399780
rect 385728 399834 385784 399843
rect 385728 399769 385784 399778
rect 385834 399786 385862 400044
rect 385926 399906 385954 400044
rect 386018 399906 386046 400044
rect 385914 399900 385966 399906
rect 385914 399842 385966 399848
rect 386006 399900 386058 399906
rect 386006 399842 386058 399848
rect 385834 399758 386000 399786
rect 385282 399724 385356 399752
rect 385222 399664 385278 399673
rect 385222 399599 385278 399608
rect 385236 397338 385264 399599
rect 385328 397526 385356 399724
rect 385420 399724 385494 399752
rect 385316 397520 385368 397526
rect 385316 397462 385368 397468
rect 385420 397361 385448 399724
rect 385684 399696 385736 399702
rect 385684 399638 385736 399644
rect 385868 399696 385920 399702
rect 385868 399638 385920 399644
rect 385592 399492 385644 399498
rect 385592 399434 385644 399440
rect 385406 397352 385462 397361
rect 385236 397310 385356 397338
rect 385224 396704 385276 396710
rect 385224 396646 385276 396652
rect 384960 394666 385080 394694
rect 385052 315314 385080 394666
rect 385132 394188 385184 394194
rect 385132 394130 385184 394136
rect 385144 315897 385172 394130
rect 385236 316742 385264 396646
rect 385328 330546 385356 397310
rect 385406 397287 385462 397296
rect 385500 396160 385552 396166
rect 385500 396102 385552 396108
rect 385408 395616 385460 395622
rect 385408 395558 385460 395564
rect 385316 330540 385368 330546
rect 385316 330482 385368 330488
rect 385316 327072 385368 327078
rect 385316 327014 385368 327020
rect 385328 325786 385356 327014
rect 385316 325780 385368 325786
rect 385316 325722 385368 325728
rect 385328 325145 385356 325722
rect 385314 325136 385370 325145
rect 385314 325071 385370 325080
rect 385420 323678 385448 395558
rect 385512 325694 385540 396102
rect 385604 327078 385632 399434
rect 385696 398886 385724 399638
rect 385776 399628 385828 399634
rect 385776 399570 385828 399576
rect 385684 398880 385736 398886
rect 385684 398822 385736 398828
rect 385684 397384 385736 397390
rect 385684 397326 385736 397332
rect 385696 334626 385724 397326
rect 385788 394194 385816 399570
rect 385880 396710 385908 399638
rect 385972 397390 386000 399758
rect 386110 399684 386138 400044
rect 386202 399838 386230 400044
rect 386190 399832 386242 399838
rect 386190 399774 386242 399780
rect 386294 399752 386322 400044
rect 386386 399945 386414 400044
rect 386372 399936 386428 399945
rect 386372 399871 386428 399880
rect 386478 399752 386506 400044
rect 386570 399906 386598 400044
rect 386558 399900 386610 399906
rect 386558 399842 386610 399848
rect 386662 399786 386690 400044
rect 386754 399838 386782 400044
rect 386616 399758 386690 399786
rect 386742 399832 386794 399838
rect 386846 399809 386874 400044
rect 386742 399774 386794 399780
rect 386832 399800 386888 399809
rect 386294 399724 386368 399752
rect 386478 399724 386552 399752
rect 386064 399656 386138 399684
rect 385960 397384 386012 397390
rect 385960 397326 386012 397332
rect 385868 396704 385920 396710
rect 385868 396646 385920 396652
rect 385776 394188 385828 394194
rect 385776 394130 385828 394136
rect 386064 394126 386092 399656
rect 386236 399628 386288 399634
rect 386236 399570 386288 399576
rect 386248 396166 386276 399570
rect 386236 396160 386288 396166
rect 386236 396102 386288 396108
rect 386340 395622 386368 399724
rect 386420 399628 386472 399634
rect 386420 399570 386472 399576
rect 386432 397730 386460 399570
rect 386524 398154 386552 399724
rect 386616 398410 386644 399758
rect 386832 399735 386888 399744
rect 386938 399752 386966 400044
rect 387030 399906 387058 400044
rect 387018 399900 387070 399906
rect 387018 399842 387070 399848
rect 387122 399838 387150 400044
rect 387214 399906 387242 400044
rect 387202 399900 387254 399906
rect 387202 399842 387254 399848
rect 387110 399832 387162 399838
rect 387110 399774 387162 399780
rect 386938 399724 387012 399752
rect 386788 399696 386840 399702
rect 386788 399638 386840 399644
rect 386604 398404 386656 398410
rect 386604 398346 386656 398352
rect 386524 398126 386644 398154
rect 386512 398064 386564 398070
rect 386512 398006 386564 398012
rect 386420 397724 386472 397730
rect 386420 397666 386472 397672
rect 386420 397452 386472 397458
rect 386420 397394 386472 397400
rect 386328 395616 386380 395622
rect 386328 395558 386380 395564
rect 386052 394120 386104 394126
rect 386052 394062 386104 394068
rect 386432 388482 386460 397394
rect 386524 393242 386552 398006
rect 386512 393236 386564 393242
rect 386512 393178 386564 393184
rect 386420 388476 386472 388482
rect 386420 388418 386472 388424
rect 385684 334620 385736 334626
rect 385684 334562 385736 334568
rect 385776 330540 385828 330546
rect 385776 330482 385828 330488
rect 385592 327072 385644 327078
rect 385592 327014 385644 327020
rect 385684 325712 385736 325718
rect 385512 325666 385684 325694
rect 385408 323672 385460 323678
rect 385408 323614 385460 323620
rect 385512 317393 385540 325666
rect 385684 325654 385736 325660
rect 385788 322318 385816 330482
rect 385776 322312 385828 322318
rect 385776 322254 385828 322260
rect 386616 321609 386644 398126
rect 386696 397044 386748 397050
rect 386696 396986 386748 396992
rect 386708 326369 386736 396986
rect 386800 330449 386828 399638
rect 386880 399628 386932 399634
rect 386880 399570 386932 399576
rect 386892 345014 386920 399570
rect 386984 398206 387012 399724
rect 387306 399684 387334 400044
rect 387524 399900 387576 399906
rect 387524 399842 387576 399848
rect 387154 399664 387210 399673
rect 387154 399599 387210 399608
rect 387260 399656 387334 399684
rect 386972 398200 387024 398206
rect 386972 398142 387024 398148
rect 386972 398064 387024 398070
rect 386972 398006 387024 398012
rect 386984 355337 387012 398006
rect 386970 355328 387026 355337
rect 386970 355263 387026 355272
rect 386892 344986 387012 345014
rect 386786 330440 386842 330449
rect 386786 330375 386842 330384
rect 386984 329866 387012 344986
rect 386972 329860 387024 329866
rect 386972 329802 387024 329808
rect 386984 329089 387012 329802
rect 386970 329080 387026 329089
rect 386970 329015 387026 329024
rect 386694 326360 386750 326369
rect 386694 326295 386750 326304
rect 386602 321600 386658 321609
rect 386602 321535 386658 321544
rect 387062 321600 387118 321609
rect 387062 321535 387118 321544
rect 385498 317384 385554 317393
rect 385498 317319 385554 317328
rect 385224 316736 385276 316742
rect 385224 316678 385276 316684
rect 385130 315888 385186 315897
rect 385130 315823 385186 315832
rect 385040 315308 385092 315314
rect 385040 315250 385092 315256
rect 384854 308952 384910 308961
rect 384854 308887 384910 308896
rect 383198 308680 383254 308689
rect 383198 308615 383254 308624
rect 380348 303214 380400 303220
rect 383014 303240 383070 303249
rect 383014 303175 383070 303184
rect 378692 299396 378744 299402
rect 378692 299338 378744 299344
rect 382280 248532 382332 248538
rect 382280 248474 382332 248480
rect 380900 142928 380952 142934
rect 380900 142870 380952 142876
rect 380912 16574 380940 142870
rect 382292 16574 382320 248474
rect 385040 244452 385092 244458
rect 385040 244394 385092 244400
rect 383660 138712 383712 138718
rect 383660 138654 383712 138660
rect 383672 16574 383700 138654
rect 385052 16574 385080 244394
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 382292 16546 382412 16574
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 378048 3596 378100 3602
rect 378048 3538 378100 3544
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379978 9480 380034 9489
rect 379978 9415 380034 9424
rect 379992 480 380020 9415
rect 381188 480 381216 16546
rect 382384 480 382412 16546
rect 383568 9036 383620 9042
rect 383568 8978 383620 8984
rect 383580 480 383608 8978
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 387076 3398 387104 321535
rect 387168 310457 387196 399599
rect 387260 397050 387288 399656
rect 387340 397724 387392 397730
rect 387340 397666 387392 397672
rect 387248 397044 387300 397050
rect 387248 396986 387300 396992
rect 387352 312905 387380 397666
rect 387536 397458 387564 399842
rect 387720 398070 387748 400302
rect 390192 400318 390244 400324
rect 387798 400279 387854 400288
rect 387892 400104 387944 400110
rect 387892 400046 387944 400052
rect 390006 400072 390062 400081
rect 387800 399424 387852 399430
rect 387800 399366 387852 399372
rect 387708 398064 387760 398070
rect 387708 398006 387760 398012
rect 387524 397452 387576 397458
rect 387524 397394 387576 397400
rect 387338 312896 387394 312905
rect 387338 312831 387394 312840
rect 387154 310448 387210 310457
rect 387154 310383 387210 310392
rect 387812 309602 387840 399366
rect 387904 312662 387932 400046
rect 387984 400036 388036 400042
rect 390006 400007 390062 400016
rect 387984 399978 388036 399984
rect 387996 314265 388024 399978
rect 389180 399560 389232 399566
rect 388166 399528 388222 399537
rect 389180 399502 389232 399508
rect 388166 399463 388222 399472
rect 388076 398676 388128 398682
rect 388076 398618 388128 398624
rect 388088 314537 388116 398618
rect 388180 320793 388208 399463
rect 388444 368552 388496 368558
rect 388444 368494 388496 368500
rect 388456 325650 388484 368494
rect 388444 325644 388496 325650
rect 388444 325586 388496 325592
rect 388166 320784 388222 320793
rect 388166 320719 388222 320728
rect 388074 314528 388130 314537
rect 388074 314463 388130 314472
rect 387982 314256 388038 314265
rect 387982 314191 388038 314200
rect 387892 312656 387944 312662
rect 387892 312598 387944 312604
rect 387800 309596 387852 309602
rect 387800 309538 387852 309544
rect 389192 289134 389220 399502
rect 389272 398608 389324 398614
rect 389272 398550 389324 398556
rect 389284 313274 389312 398550
rect 389548 398472 389600 398478
rect 389548 398414 389600 398420
rect 389456 397520 389508 397526
rect 389456 397462 389508 397468
rect 389364 397248 389416 397254
rect 389364 397190 389416 397196
rect 389376 314673 389404 397190
rect 389362 314664 389418 314673
rect 389362 314599 389418 314608
rect 389468 314401 389496 397462
rect 389560 317354 389588 398414
rect 390020 396914 390048 400007
rect 390204 399974 390232 400318
rect 390192 399968 390244 399974
rect 390192 399910 390244 399916
rect 390834 399936 390890 399945
rect 390834 399871 390890 399880
rect 390652 398540 390704 398546
rect 390652 398482 390704 398488
rect 390560 398268 390612 398274
rect 390560 398210 390612 398216
rect 390008 396908 390060 396914
rect 390008 396850 390060 396856
rect 389640 394120 389692 394126
rect 389640 394062 389692 394068
rect 389652 333266 389680 394062
rect 389640 333260 389692 333266
rect 389640 333202 389692 333208
rect 389548 317348 389600 317354
rect 389548 317290 389600 317296
rect 389454 314392 389510 314401
rect 389454 314327 389510 314336
rect 389272 313268 389324 313274
rect 389272 313210 389324 313216
rect 390572 303618 390600 398210
rect 390560 303612 390612 303618
rect 390560 303554 390612 303560
rect 390664 303550 390692 398482
rect 390744 395140 390796 395146
rect 390744 395082 390796 395088
rect 390756 309670 390784 395082
rect 390848 314022 390876 399871
rect 392032 398404 392084 398410
rect 392032 398346 392084 398352
rect 391938 398168 391994 398177
rect 391938 398103 391994 398112
rect 390836 314016 390888 314022
rect 390836 313958 390888 313964
rect 390744 309664 390796 309670
rect 390744 309606 390796 309612
rect 390652 303544 390704 303550
rect 391952 303521 391980 398103
rect 392044 311545 392072 398346
rect 392136 311817 392164 400454
rect 394792 400376 394844 400382
rect 394792 400318 394844 400324
rect 392214 399392 392270 399401
rect 392214 399327 392270 399336
rect 392228 313177 392256 399327
rect 394700 398880 394752 398886
rect 394700 398822 394752 398828
rect 392214 313168 392270 313177
rect 392214 313103 392270 313112
rect 392122 311808 392178 311817
rect 392122 311743 392178 311752
rect 392030 311536 392086 311545
rect 392030 311471 392086 311480
rect 394712 311137 394740 398822
rect 394804 312497 394832 400318
rect 394884 396908 394936 396914
rect 394884 396850 394936 396856
rect 394896 317422 394924 396850
rect 580264 386436 580316 386442
rect 580264 386378 580316 386384
rect 580276 378457 580304 386378
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 523684 370660 523736 370666
rect 523684 370602 523736 370608
rect 498200 334008 498252 334014
rect 498200 333950 498252 333956
rect 484400 332648 484452 332654
rect 484400 332590 484452 332596
rect 416778 328536 416834 328545
rect 416778 328471 416834 328480
rect 396080 324964 396132 324970
rect 396080 324906 396132 324912
rect 394884 317416 394936 317422
rect 394884 317358 394936 317364
rect 395988 317416 396040 317422
rect 395988 317358 396040 317364
rect 396000 316742 396028 317358
rect 395988 316736 396040 316742
rect 395988 316678 396040 316684
rect 394790 312488 394846 312497
rect 394790 312423 394846 312432
rect 394698 311128 394754 311137
rect 394698 311063 394754 311072
rect 390652 303486 390704 303492
rect 391938 303512 391994 303521
rect 391938 303447 391994 303456
rect 389180 289128 389232 289134
rect 389180 289070 389232 289076
rect 389180 262880 389232 262886
rect 389180 262822 389232 262828
rect 387800 131776 387852 131782
rect 387800 131718 387852 131724
rect 387154 9344 387210 9353
rect 387154 9279 387210 9288
rect 387064 3392 387116 3398
rect 387064 3334 387116 3340
rect 387168 480 387196 9279
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 131718
rect 389192 16574 389220 262822
rect 391940 257372 391992 257378
rect 391940 257314 391992 257320
rect 390560 133272 390612 133278
rect 390560 133214 390612 133220
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3466 390600 133214
rect 391952 16574 391980 257314
rect 394700 123548 394752 123554
rect 394700 123490 394752 123496
rect 394712 16574 394740 123490
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 390650 6216 390706 6225
rect 390650 6151 390706 6160
rect 390560 3460 390612 3466
rect 390560 3402 390612 3408
rect 390664 480 390692 6151
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 391860 480 391888 3402
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394238 9208 394294 9217
rect 394238 9143 394294 9152
rect 394252 480 394280 9143
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 324906
rect 398930 324456 398986 324465
rect 398930 324391 398986 324400
rect 397460 165640 397512 165646
rect 397460 165582 397512 165588
rect 397472 16574 397500 165582
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398840 3732 398892 3738
rect 398840 3674 398892 3680
rect 398852 1850 398880 3674
rect 398944 3398 398972 324391
rect 402980 291848 403032 291854
rect 402980 291790 403032 291796
rect 400220 79348 400272 79354
rect 400220 79290 400272 79296
rect 400232 16574 400260 79290
rect 402992 16574 403020 291790
rect 414020 263696 414072 263702
rect 414020 263638 414072 263644
rect 407120 248464 407172 248470
rect 407120 248406 407172 248412
rect 405740 137352 405792 137358
rect 405740 137294 405792 137300
rect 404360 112464 404412 112470
rect 404360 112406 404412 112412
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 1822 398972 1850
rect 398944 480 398972 1822
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 3664 402572 3670
rect 402520 3606 402572 3612
rect 402532 480 402560 3606
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 112406
rect 405752 16574 405780 137294
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3210 407160 248406
rect 409880 247172 409932 247178
rect 409880 247114 409932 247120
rect 408500 130416 408552 130422
rect 408500 130358 408552 130364
rect 407210 54496 407266 54505
rect 407210 54431 407266 54440
rect 407224 3398 407252 54431
rect 408512 16574 408540 130358
rect 409892 16574 409920 247114
rect 412638 122088 412694 122097
rect 412638 122023 412694 122032
rect 411258 51776 411314 51785
rect 411258 51711 411314 51720
rect 411272 16574 411300 51711
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 122023
rect 414032 16574 414060 263638
rect 415400 146940 415452 146946
rect 415400 146882 415452 146888
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3534 415440 146882
rect 416792 16574 416820 328471
rect 477498 313984 477554 313993
rect 466460 313948 466512 313954
rect 477498 313919 477554 313928
rect 466460 313890 466512 313896
rect 431960 307080 432012 307086
rect 431960 307022 432012 307028
rect 427820 255332 427872 255338
rect 427820 255274 427872 255280
rect 423772 251320 423824 251326
rect 423772 251262 423824 251268
rect 419540 141568 419592 141574
rect 419540 141510 419592 141516
rect 419552 16574 419580 141510
rect 422944 129124 422996 129130
rect 422944 129066 422996 129072
rect 416792 16546 417464 16574
rect 419552 16546 420224 16574
rect 415490 9072 415546 9081
rect 415490 9007 415546 9016
rect 415400 3528 415452 3534
rect 415400 3470 415452 3476
rect 415504 480 415532 9007
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 416700 480 416728 3470
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418988 8968 419040 8974
rect 418988 8910 419040 8916
rect 419000 480 419028 8910
rect 420196 480 420224 16546
rect 422574 8936 422630 8945
rect 422574 8871 422630 8880
rect 421380 3392 421432 3398
rect 421380 3334 421432 3340
rect 421392 480 421420 3334
rect 422588 480 422616 8871
rect 422956 3534 422984 129066
rect 423784 3670 423812 251262
rect 425060 174004 425112 174010
rect 425060 173946 425112 173952
rect 425072 16574 425100 173946
rect 426438 120728 426494 120737
rect 426438 120663 426494 120672
rect 426452 16574 426480 120663
rect 427832 16574 427860 255274
rect 431222 156632 431278 156641
rect 431222 156567 431278 156576
rect 430578 30968 430634 30977
rect 430578 30903 430634 30912
rect 430592 16574 430620 30903
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 423772 3664 423824 3670
rect 423772 3606 423824 3612
rect 424968 3664 425020 3670
rect 424968 3606 425020 3612
rect 422944 3528 422996 3534
rect 422944 3470 422996 3476
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 423784 480 423812 3470
rect 424980 480 425008 3606
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429200 15904 429252 15910
rect 429200 15846 429252 15852
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 15846
rect 430868 480 430896 16546
rect 431236 4010 431264 156567
rect 431224 4004 431276 4010
rect 431224 3946 431276 3952
rect 431972 3346 432000 307022
rect 445760 263628 445812 263634
rect 445760 263570 445812 263576
rect 441620 258120 441672 258126
rect 441620 258062 441672 258068
rect 438860 250504 438912 250510
rect 438860 250446 438912 250452
rect 434720 245676 434772 245682
rect 434720 245618 434772 245624
rect 432052 173936 432104 173942
rect 432052 173878 432104 173884
rect 432064 3534 432092 173878
rect 434732 16574 434760 245618
rect 436744 144288 436796 144294
rect 436744 144230 436796 144236
rect 434732 16546 435128 16574
rect 434444 4004 434496 4010
rect 434444 3946 434496 3952
rect 432052 3528 432104 3534
rect 432052 3470 432104 3476
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 431972 3318 432092 3346
rect 432064 480 432092 3318
rect 433260 480 433288 3470
rect 434456 480 434484 3946
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 436652 6180 436704 6186
rect 436652 6122 436704 6128
rect 436664 3074 436692 6122
rect 436756 3534 436784 144230
rect 438872 16574 438900 250446
rect 440240 135924 440292 135930
rect 440240 135866 440292 135872
rect 438872 16546 439176 16574
rect 436744 3528 436796 3534
rect 436744 3470 436796 3476
rect 437940 3528 437992 3534
rect 437940 3470 437992 3476
rect 436664 3046 436784 3074
rect 436756 480 436784 3046
rect 437952 480 437980 3470
rect 439148 480 439176 16546
rect 440252 3534 440280 135866
rect 441632 16574 441660 258062
rect 443000 186380 443052 186386
rect 443000 186322 443052 186328
rect 443012 16574 443040 186322
rect 444380 127628 444432 127634
rect 444380 127570 444432 127576
rect 444392 16574 444420 127570
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 440330 11656 440386 11665
rect 440330 11591 440386 11600
rect 440240 3528 440292 3534
rect 440240 3470 440292 3476
rect 440344 480 440372 11591
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 441540 480 441568 3470
rect 442644 480 442672 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 263570
rect 452660 262268 452712 262274
rect 452660 262210 452712 262216
rect 448612 252680 448664 252686
rect 448612 252622 448664 252628
rect 447140 167068 447192 167074
rect 447140 167010 447192 167016
rect 447152 16574 447180 167010
rect 447782 118008 447838 118017
rect 447782 117943 447838 117952
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 447796 3534 447824 117943
rect 448624 3670 448652 252622
rect 451280 149728 451332 149734
rect 451280 149670 451332 149676
rect 449900 142860 449952 142866
rect 449900 142802 449952 142808
rect 449912 16574 449940 142802
rect 451292 16574 451320 149670
rect 452672 16574 452700 262210
rect 459560 247104 459612 247110
rect 459560 247046 459612 247052
rect 456800 244384 456852 244390
rect 456800 244326 456852 244332
rect 455420 134632 455472 134638
rect 455420 134574 455472 134580
rect 454038 98696 454094 98705
rect 454038 98631 454094 98640
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3664 448664 3670
rect 448612 3606 448664 3612
rect 449808 3664 449860 3670
rect 449808 3606 449860 3612
rect 447784 3528 447836 3534
rect 447784 3470 447836 3476
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 448624 480 448652 3470
rect 449820 480 449848 3606
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 98631
rect 455432 16574 455460 134574
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3346 456840 244326
rect 458180 126336 458232 126342
rect 458180 126278 458232 126284
rect 456890 46200 456946 46209
rect 456890 46135 456946 46144
rect 456904 3534 456932 46135
rect 458192 16574 458220 126278
rect 459572 16574 459600 247046
rect 462320 116612 462372 116618
rect 462320 116554 462372 116560
rect 460938 44840 460994 44849
rect 460938 44775 460994 44784
rect 460952 16574 460980 44775
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456812 3318 456932 3346
rect 456904 480 456932 3318
rect 458100 480 458128 3470
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 116554
rect 465078 115152 465134 115161
rect 465078 115087 465134 115096
rect 463976 3596 464028 3602
rect 463976 3538 464028 3544
rect 463988 480 464016 3538
rect 465092 3534 465120 115087
rect 466472 16574 466500 313890
rect 470600 256760 470652 256766
rect 470600 256702 470652 256708
rect 467840 175296 467892 175302
rect 467840 175238 467892 175244
rect 467852 16574 467880 175238
rect 468482 131744 468538 131753
rect 468482 131679 468538 131688
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 465172 13116 465224 13122
rect 465172 13058 465224 13064
rect 465080 3528 465132 3534
rect 465080 3470 465132 3476
rect 465184 480 465212 13058
rect 465908 3528 465960 3534
rect 465908 3470 465960 3476
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465920 354 465948 3470
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 3534 468524 131679
rect 468484 3528 468536 3534
rect 468484 3470 468536 3476
rect 469864 3528 469916 3534
rect 469864 3470 469916 3476
rect 469876 480 469904 3470
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 256702
rect 471244 243024 471296 243030
rect 471244 242966 471296 242972
rect 471256 3602 471284 242966
rect 472622 124808 472678 124817
rect 472622 124743 472678 124752
rect 472256 10328 472308 10334
rect 472256 10270 472308 10276
rect 471244 3596 471296 3602
rect 471244 3538 471296 3544
rect 472268 480 472296 10270
rect 472636 3534 472664 124743
rect 476118 113792 476174 113801
rect 476118 113727 476174 113736
rect 474738 42120 474794 42129
rect 474738 42055 474794 42064
rect 474752 16574 474780 42055
rect 476132 16574 476160 113727
rect 477512 16574 477540 313919
rect 481640 241596 481692 241602
rect 481640 241538 481692 241544
rect 480260 129056 480312 129062
rect 480260 128998 480312 129004
rect 480272 16574 480300 128998
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 474556 3596 474608 3602
rect 474556 3538 474608 3544
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 474568 480 474596 3538
rect 475764 480 475792 16546
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 478880 11756 478932 11762
rect 478880 11698 478932 11704
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 11698
rect 480548 480 480576 16546
rect 481652 6914 481680 241538
rect 481732 169788 481784 169794
rect 481732 169730 481784 169736
rect 481744 16574 481772 169730
rect 483020 153332 483072 153338
rect 483020 153274 483072 153280
rect 483032 16574 483060 153274
rect 484412 16574 484440 332590
rect 495440 273284 495492 273290
rect 495440 273226 495492 273232
rect 491300 251252 491352 251258
rect 491300 251194 491352 251200
rect 488540 241528 488592 241534
rect 488540 241470 488592 241476
rect 485778 109712 485834 109721
rect 485778 109647 485834 109656
rect 485792 16574 485820 109647
rect 487158 37904 487214 37913
rect 487158 37839 487214 37848
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 37839
rect 488552 16574 488580 241470
rect 489920 126268 489972 126274
rect 489920 126210 489972 126216
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3534 489960 126210
rect 490010 18592 490066 18601
rect 490010 18527 490066 18536
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 18527
rect 491312 16574 491340 251194
rect 494060 155304 494112 155310
rect 494060 155246 494112 155252
rect 492680 108316 492732 108322
rect 492680 108258 492732 108264
rect 492692 16574 492720 108258
rect 494072 16574 494100 155246
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 273226
rect 496818 106856 496874 106865
rect 496818 106791 496874 106800
rect 496832 16574 496860 106791
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 3534 498240 333950
rect 513378 329896 513434 329905
rect 513378 329831 513434 329840
rect 502340 312588 502392 312594
rect 502340 312530 502392 312536
rect 498290 151056 498346 151065
rect 498290 150991 498346 151000
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 150991
rect 500958 148472 501014 148481
rect 500958 148407 501014 148416
rect 499580 105596 499632 105602
rect 499580 105538 499632 105544
rect 499592 16574 499620 105538
rect 500972 16574 501000 148407
rect 502352 16574 502380 312530
rect 507124 244316 507176 244322
rect 507124 244258 507176 244264
rect 506480 238876 506532 238882
rect 506480 238818 506532 238824
rect 503720 123480 503772 123486
rect 503720 123422 503772 123428
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 123422
rect 505100 17264 505152 17270
rect 505100 17206 505152 17212
rect 505112 16574 505140 17206
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 238818
rect 506570 104136 506626 104145
rect 506570 104071 506626 104080
rect 506584 16574 506612 104071
rect 506584 16546 507072 16574
rect 507044 490 507072 16546
rect 507136 4078 507164 244258
rect 507860 153264 507912 153270
rect 507860 153206 507912 153212
rect 507872 16574 507900 153206
rect 512000 152584 512052 152590
rect 512000 152526 512052 152532
rect 510620 102808 510672 102814
rect 510620 102750 510672 102756
rect 510632 16574 510660 102750
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 507124 4072 507176 4078
rect 507124 4014 507176 4020
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507044 462 507256 490
rect 508884 480 508912 16546
rect 510068 4072 510120 4078
rect 510068 4014 510120 4020
rect 510080 480 510108 4014
rect 511276 480 511304 16546
rect 507228 354 507256 462
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 152526
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 329831
rect 523696 313274 523724 370602
rect 580724 370592 580776 370598
rect 580724 370534 580776 370540
rect 580356 370524 580408 370530
rect 580356 370466 580408 370472
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580262 364984 580318 364993
rect 580262 364919 580318 364928
rect 569960 329860 570012 329866
rect 569960 329802 570012 329808
rect 547880 325780 547932 325786
rect 547880 325722 547932 325728
rect 527824 316736 527876 316742
rect 527824 316678 527876 316684
rect 523684 313268 523736 313274
rect 523684 313210 523736 313216
rect 516140 276072 516192 276078
rect 516140 276014 516192 276020
rect 514024 145580 514076 145586
rect 514024 145522 514076 145528
rect 514036 3058 514064 145522
rect 514850 101416 514906 101425
rect 514850 101351 514906 101360
rect 514864 6914 514892 101351
rect 516152 16574 516180 276014
rect 527180 253972 527232 253978
rect 527180 253914 527232 253920
rect 523132 252612 523184 252618
rect 523132 252554 523184 252560
rect 520280 242956 520332 242962
rect 520280 242898 520332 242904
rect 518900 155984 518952 155990
rect 518900 155926 518952 155932
rect 517518 71088 517574 71097
rect 517518 71023 517574 71032
rect 517532 16574 517560 71023
rect 518912 16574 518940 155926
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 514772 6886 514892 6914
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 6886
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 242898
rect 522304 155236 522356 155242
rect 522304 155178 522356 155184
rect 520924 122120 520976 122126
rect 520924 122062 520976 122068
rect 520936 3534 520964 122062
rect 522316 3534 522344 155178
rect 523144 16574 523172 252554
rect 525800 36576 525852 36582
rect 525800 36518 525852 36524
rect 524420 28280 524472 28286
rect 524420 28222 524472 28228
rect 524432 16574 524460 28222
rect 525812 16574 525840 36518
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 520924 3528 520976 3534
rect 520924 3470 520976 3476
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 522304 3528 522356 3534
rect 522304 3470 522356 3476
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 521856 480 521884 3470
rect 523052 480 523080 3470
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527192 6914 527220 253914
rect 527836 16574 527864 316678
rect 538220 289128 538272 289134
rect 538220 289070 538272 289076
rect 531320 277432 531372 277438
rect 531320 277374 531372 277380
rect 529938 149696 529994 149705
rect 529938 149631 529994 149640
rect 528558 69592 528614 69601
rect 528558 69527 528614 69536
rect 527836 16546 527956 16574
rect 527192 6886 527864 6914
rect 527836 480 527864 6886
rect 527928 3534 527956 16546
rect 527916 3528 527968 3534
rect 527916 3470 527968 3476
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 69527
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 149631
rect 531332 480 531360 277374
rect 534080 249824 534132 249830
rect 534080 249766 534132 249772
rect 532700 144220 532752 144226
rect 532700 144162 532752 144168
rect 531410 95840 531466 95849
rect 531410 95775 531466 95784
rect 531424 16574 531452 95775
rect 532712 16574 532740 144162
rect 534092 16574 534120 249766
rect 536104 152516 536156 152522
rect 536104 152458 536156 152464
rect 535460 94512 535512 94518
rect 535460 94454 535512 94460
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 535472 6914 535500 94454
rect 536116 16574 536144 152458
rect 536838 119368 536894 119377
rect 536838 119303 536894 119312
rect 536852 16574 536880 119303
rect 536116 16546 536236 16574
rect 536852 16546 537248 16574
rect 535472 6886 536144 6914
rect 536116 480 536144 6886
rect 536208 3058 536236 16546
rect 536196 3052 536248 3058
rect 536196 2994 536248 3000
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 289070
rect 543004 266416 543056 266422
rect 543004 266358 543056 266364
rect 540980 238808 541032 238814
rect 540980 238750 541032 238756
rect 539692 120760 539744 120766
rect 539692 120702 539744 120708
rect 539704 6914 539732 120702
rect 540992 16574 541020 238750
rect 542360 93152 542412 93158
rect 542360 93094 542412 93100
rect 542372 16574 542400 93094
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 539612 6886 539732 6914
rect 539612 480 539640 6886
rect 540796 3052 540848 3058
rect 540796 2994 540848 3000
rect 540808 480 540836 2994
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3126 543044 266358
rect 543738 148336 543794 148345
rect 543738 148271 543794 148280
rect 543752 16574 543780 148271
rect 546500 91792 546552 91798
rect 546500 91734 546552 91740
rect 543752 16546 544424 16574
rect 543004 3120 543056 3126
rect 543004 3062 543056 3068
rect 544396 480 544424 16546
rect 545488 3120 545540 3126
rect 545488 3062 545540 3068
rect 545500 480 545528 3062
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 91734
rect 547892 3602 547920 325722
rect 563060 325712 563112 325718
rect 563060 325654 563112 325660
rect 556250 311128 556306 311137
rect 556250 311063 556306 311072
rect 550640 141432 550692 141438
rect 550640 141374 550692 141380
rect 549904 134564 549956 134570
rect 549904 134506 549956 134512
rect 548522 90400 548578 90409
rect 548522 90335 548578 90344
rect 547970 35184 548026 35193
rect 547970 35119 548026 35128
rect 547880 3596 547932 3602
rect 547880 3538 547932 3544
rect 547984 3482 548012 35119
rect 547892 3454 548012 3482
rect 547892 480 547920 3454
rect 548536 2990 548564 90335
rect 549916 3602 549944 134506
rect 550652 16574 550680 141374
rect 554780 137284 554832 137290
rect 554780 137226 554832 137232
rect 552664 89004 552716 89010
rect 552664 88946 552716 88952
rect 550652 16546 551048 16574
rect 548708 3596 548760 3602
rect 548708 3538 548760 3544
rect 549904 3596 549956 3602
rect 549904 3538 549956 3544
rect 548524 2984 548576 2990
rect 548524 2926 548576 2932
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3538
rect 550272 2984 550324 2990
rect 550272 2926 550324 2932
rect 550284 480 550312 2926
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 3670 552704 88946
rect 553400 87644 553452 87650
rect 553400 87586 553452 87592
rect 553412 16574 553440 87586
rect 553412 16546 553808 16574
rect 552664 3664 552716 3670
rect 552664 3606 552716 3612
rect 552664 3528 552716 3534
rect 552664 3470 552716 3476
rect 552676 480 552704 3470
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 137226
rect 556264 6914 556292 311063
rect 558920 239420 558972 239426
rect 558920 239362 558972 239368
rect 557538 153776 557594 153785
rect 557538 153711 557594 153720
rect 557552 16574 557580 153711
rect 558932 16574 558960 239362
rect 561678 146976 561734 146985
rect 561678 146911 561734 146920
rect 560300 86284 560352 86290
rect 560300 86226 560352 86232
rect 560312 16574 560340 86226
rect 561692 16574 561720 146911
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556172 6886 556292 6914
rect 556172 480 556200 6886
rect 557356 3664 557408 3670
rect 557356 3606 557408 3612
rect 557368 480 557396 3606
rect 558564 480 558592 16546
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 325654
rect 568580 135312 568632 135318
rect 568580 135254 568632 135260
rect 564438 84824 564494 84833
rect 564438 84759 564494 84768
rect 564452 480 564480 84759
rect 567200 82136 567252 82142
rect 567200 82078 567252 82084
rect 564532 33788 564584 33794
rect 564532 33730 564584 33736
rect 564544 16574 564572 33730
rect 567212 16574 567240 82078
rect 568592 16574 568620 135254
rect 569972 16574 570000 329802
rect 579988 325644 580040 325650
rect 579988 325586 580040 325592
rect 580000 325281 580028 325586
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 579620 313268 579672 313274
rect 579620 313210 579672 313216
rect 572810 312488 572866 312497
rect 572810 312423 572866 312432
rect 571982 306504 572038 306513
rect 571982 306439 572038 306448
rect 564544 16546 565216 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566832 3460 566884 3466
rect 566832 3402 566884 3408
rect 566844 480 566872 3402
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 571522 7576 571578 7585
rect 571522 7511 571578 7520
rect 571536 480 571564 7511
rect 571996 4146 572024 306439
rect 572824 16574 572852 312423
rect 579632 312089 579660 313210
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 577504 299532 577556 299538
rect 577504 299474 577556 299480
rect 577516 245614 577544 299474
rect 580172 298784 580224 298790
rect 580170 298752 580172 298761
rect 580224 298752 580226 298761
rect 580170 298687 580226 298696
rect 577504 245608 577556 245614
rect 579620 245608 579672 245614
rect 577504 245550 577556 245556
rect 579618 245576 579620 245585
rect 579672 245576 579674 245585
rect 579618 245511 579674 245520
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579988 209092 580040 209098
rect 579988 209034 580040 209040
rect 580000 205737 580028 209034
rect 579986 205728 580042 205737
rect 579986 205663 580042 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 579896 153196 579948 153202
rect 579896 153138 579948 153144
rect 579908 152697 579936 153138
rect 579894 152688 579950 152697
rect 579894 152623 579950 152632
rect 580276 139369 580304 364919
rect 580368 219065 580396 370466
rect 580632 369164 580684 369170
rect 580632 369106 580684 369112
rect 580446 366344 580502 366353
rect 580446 366279 580502 366288
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 580354 206272 580410 206281
rect 580354 206207 580410 206216
rect 580262 139360 580318 139369
rect 580262 139295 580318 139304
rect 575480 133204 575532 133210
rect 575480 133146 575532 133152
rect 574100 83496 574152 83502
rect 574100 83438 574152 83444
rect 574112 16574 574140 83438
rect 575492 16574 575520 133146
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580264 97300 580316 97306
rect 580264 97242 580316 97248
rect 580276 86193 580304 97242
rect 580262 86184 580318 86193
rect 580262 86119 580318 86128
rect 578240 80708 578292 80714
rect 578240 80650 578292 80656
rect 578252 16574 578280 80650
rect 580264 73840 580316 73846
rect 580264 73782 580316 73788
rect 580276 46345 580304 73782
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580080 20664 580132 20670
rect 580080 20606 580132 20612
rect 580092 19825 580120 20606
rect 580078 19816 580134 19825
rect 580078 19751 580134 19760
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 571984 4140 572036 4146
rect 571984 4082 572036 4088
rect 572720 3596 572772 3602
rect 572720 3538 572772 3544
rect 572732 480 572760 3538
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 578620 480 578648 16546
rect 580368 6633 580396 206207
rect 580460 179217 580488 366279
rect 580538 360904 580594 360913
rect 580538 360839 580594 360848
rect 580552 258913 580580 360839
rect 580644 272241 580672 369106
rect 580736 351937 580764 370534
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580630 272232 580686 272241
rect 580630 272167 580686 272176
rect 580538 258904 580594 258913
rect 580538 258839 580594 258848
rect 580722 209128 580778 209137
rect 580722 209063 580778 209072
rect 580538 208992 580594 209001
rect 580538 208927 580594 208936
rect 580446 179208 580502 179217
rect 580446 179143 580502 179152
rect 580552 126041 580580 208927
rect 580736 165889 580764 209063
rect 580722 165880 580778 165889
rect 580722 165815 580778 165824
rect 580538 126032 580594 126041
rect 580538 125967 580594 125976
rect 580354 6624 580410 6633
rect 580354 6559 580410 6568
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 6918 450472 6974 450528
rect 4066 410488 4122 410544
rect 71778 404232 71834 404288
rect 3422 397432 3478 397488
rect 265806 402056 265862 402112
rect 263322 401784 263378 401840
rect 256606 398112 256662 398168
rect 220450 373224 220506 373280
rect 3238 371320 3294 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 204166 322088 204222 322144
rect 3422 319232 3478 319288
rect 4066 306176 4122 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 158626 241712 158682 241768
rect 151726 241576 151782 241632
rect 3330 241032 3386 241088
rect 150254 228384 150310 228440
rect 3146 214920 3202 214976
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3330 149776 3386 149832
rect 3054 136720 3110 136776
rect 3330 110608 3386 110664
rect 3054 58520 3110 58576
rect 2870 32408 2926 32464
rect 3698 162832 3754 162888
rect 3606 97552 3662 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 19352 3478 19408
rect 6918 153720 6974 153776
rect 3422 6432 3478 6488
rect 16578 146920 16634 146976
rect 31022 148280 31078 148336
rect 33138 144064 33194 144120
rect 32402 130328 32458 130384
rect 44822 113736 44878 113792
rect 44178 112376 44234 112432
rect 51078 152360 51134 152416
rect 52458 131688 52514 131744
rect 59358 137264 59414 137320
rect 62118 138624 62174 138680
rect 71778 153856 71834 153912
rect 71042 149640 71098 149696
rect 80058 139984 80114 140040
rect 89718 147056 89774 147112
rect 88982 145560 89038 145616
rect 93858 145696 93914 145752
rect 100758 149776 100814 149832
rect 103518 148416 103574 148472
rect 107658 144200 107714 144256
rect 110418 141344 110474 141400
rect 116582 148552 116638 148608
rect 121458 140120 121514 140176
rect 127622 149912 127678 149968
rect 126978 134408 127034 134464
rect 129738 111016 129794 111072
rect 131118 153992 131174 154048
rect 136638 126248 136694 126304
rect 146942 209072 146998 209128
rect 143630 135904 143686 135960
rect 149150 159024 149206 159080
rect 150254 159024 150310 159080
rect 147678 141480 147734 141536
rect 151174 160112 151230 160168
rect 151542 160112 151598 160168
rect 150438 158480 150494 158536
rect 150530 140664 150586 140720
rect 150530 139984 150586 140040
rect 151634 158480 151690 158536
rect 151174 148280 151230 148336
rect 154210 240216 154266 240272
rect 153014 239400 153070 239456
rect 151726 140664 151782 140720
rect 151910 150456 151966 150512
rect 152830 159432 152886 159488
rect 154026 158888 154082 158944
rect 153106 147600 153162 147656
rect 155866 241032 155922 241088
rect 154486 240896 154542 240952
rect 154394 233008 154450 233064
rect 154026 149776 154082 149832
rect 154394 146240 154450 146296
rect 154578 153040 154634 153096
rect 154486 146104 154542 146160
rect 155406 160248 155462 160304
rect 155314 158752 155370 158808
rect 155682 159568 155738 159624
rect 155682 158752 155738 158808
rect 157154 239536 157210 239592
rect 155866 158752 155922 158808
rect 155774 157392 155830 157448
rect 155498 156848 155554 156904
rect 155406 153720 155462 153776
rect 155866 153856 155922 153912
rect 155314 149912 155370 149968
rect 156510 149640 156566 149696
rect 156694 156984 156750 157040
rect 156878 159296 156934 159352
rect 156786 156712 156842 156768
rect 156694 152360 156750 152416
rect 158350 228248 158406 228304
rect 157338 157664 157394 157720
rect 157246 157256 157302 157312
rect 157154 156984 157210 157040
rect 157338 153992 157394 154048
rect 156878 148416 156934 148472
rect 158258 157800 158314 157856
rect 158166 157664 158222 157720
rect 158258 153040 158314 153096
rect 158074 148552 158130 148608
rect 159914 241440 159970 241496
rect 159454 235184 159510 235240
rect 158718 158616 158774 158672
rect 158442 157936 158498 157992
rect 159454 159160 159510 159216
rect 159730 160384 159786 160440
rect 159914 158616 159970 158672
rect 160098 158616 160154 158672
rect 159914 158072 159970 158128
rect 159454 150456 159510 150512
rect 161110 158616 161166 158672
rect 161110 158208 161166 158264
rect 160742 157528 160798 157584
rect 164330 292712 164386 292768
rect 162766 292576 162822 292632
rect 165710 282104 165766 282160
rect 164330 212064 164386 212120
rect 166906 212064 166962 212120
rect 169758 209888 169814 209944
rect 170402 209888 170458 209944
rect 176750 289040 176806 289096
rect 180890 288496 180946 288552
rect 182914 235456 182970 235512
rect 182546 210024 182602 210080
rect 186410 288632 186466 288688
rect 187790 289176 187846 289232
rect 189814 289448 189870 289504
rect 190642 290672 190698 290728
rect 190458 289856 190514 289912
rect 190550 272448 190606 272504
rect 192206 290536 192262 290592
rect 192022 290400 192078 290456
rect 191838 289992 191894 290048
rect 190734 242120 190790 242176
rect 192482 232464 192538 232520
rect 194322 232328 194378 232384
rect 198646 210024 198702 210080
rect 164146 209480 164202 209536
rect 184846 209480 184902 209536
rect 189538 209480 189594 209536
rect 194414 209480 194470 209536
rect 195886 209480 195942 209536
rect 198462 209480 198518 209536
rect 199198 209480 199254 209536
rect 199934 209752 199990 209808
rect 199842 209480 199898 209536
rect 205546 321544 205602 321600
rect 205454 316648 205510 316704
rect 204902 307128 204958 307184
rect 204258 209480 204314 209536
rect 205086 238992 205142 239048
rect 206926 318824 206982 318880
rect 206742 318144 206798 318200
rect 206374 308488 206430 308544
rect 205546 233144 205602 233200
rect 206650 236680 206706 236736
rect 206742 219272 206798 219328
rect 206742 218864 206798 218920
rect 205546 209208 205602 209264
rect 207478 174528 207534 174584
rect 162950 159840 163006 159896
rect 162858 159704 162914 159760
rect 162490 157120 162546 157176
rect 163134 159874 163190 159930
rect 163594 159840 163650 159896
rect 163042 157392 163098 157448
rect 163318 158616 163374 158672
rect 163502 157528 163558 157584
rect 163870 159704 163926 159760
rect 164054 159840 164110 159896
rect 164238 159704 164294 159760
rect 164238 158616 164294 158672
rect 164514 159840 164570 159896
rect 164790 158616 164846 158672
rect 164698 158344 164754 158400
rect 164606 157392 164662 157448
rect 165066 159024 165122 159080
rect 165158 158616 165214 158672
rect 164974 157256 165030 157312
rect 165434 159840 165490 159896
rect 165618 159840 165674 159896
rect 165618 159296 165674 159352
rect 165710 158616 165766 158672
rect 165894 159024 165950 159080
rect 166262 159704 166318 159760
rect 166078 158616 166134 158672
rect 166078 158208 166134 158264
rect 166354 156984 166410 157040
rect 166538 159840 166594 159896
rect 166170 137944 166226 138000
rect 166170 137536 166226 137592
rect 166814 159840 166870 159896
rect 166906 159704 166962 159760
rect 166906 159024 166962 159080
rect 166814 158888 166870 158944
rect 166906 158208 166962 158264
rect 166998 157800 167054 157856
rect 166906 157664 166962 157720
rect 167274 156712 167330 156768
rect 167458 156848 167514 156904
rect 167642 159840 167698 159896
rect 167918 159704 167974 159760
rect 167826 159568 167882 159624
rect 167826 159160 167882 159216
rect 167826 158616 167882 158672
rect 167826 157936 167882 157992
rect 168010 158752 168066 158808
rect 168194 159840 168250 159896
rect 168286 158344 168342 158400
rect 168286 157664 168342 157720
rect 168470 159840 168526 159896
rect 168838 159704 168894 159760
rect 168654 158616 168710 158672
rect 168562 158344 168618 158400
rect 168562 157836 168564 157856
rect 168564 157836 168616 157856
rect 168616 157836 168618 157856
rect 168562 157800 168618 157836
rect 168654 139304 168710 139360
rect 169022 159840 169078 159896
rect 169114 158480 169170 158536
rect 169298 159568 169354 159624
rect 169574 159840 169630 159896
rect 169482 159704 169538 159760
rect 169390 158616 169446 158672
rect 169758 158888 169814 158944
rect 169666 158344 169722 158400
rect 169022 139304 169078 139360
rect 168838 139032 168894 139088
rect 169850 158616 169906 158672
rect 169666 144200 169722 144256
rect 169206 139032 169262 139088
rect 170310 159840 170366 159896
rect 170126 159568 170182 159624
rect 170678 159704 170734 159760
rect 171046 159874 171102 159930
rect 171138 159704 171194 159760
rect 170954 159316 171010 159352
rect 170954 159296 170956 159316
rect 170956 159296 171008 159316
rect 171008 159296 171010 159316
rect 171046 157276 171102 157312
rect 171046 157256 171048 157276
rect 171048 157256 171100 157276
rect 171100 157256 171102 157276
rect 171506 159840 171562 159896
rect 171690 159568 171746 159624
rect 171966 159874 172022 159930
rect 171598 159296 171654 159352
rect 171506 159160 171562 159216
rect 171506 158888 171562 158944
rect 171230 155896 171286 155952
rect 171598 158480 171654 158536
rect 171874 158616 171930 158672
rect 172058 159704 172114 159760
rect 172150 158480 172206 158536
rect 171782 131144 171838 131200
rect 172334 158616 172390 158672
rect 172610 159840 172666 159896
rect 172702 159704 172758 159760
rect 172886 159840 172942 159896
rect 172886 159160 172942 159216
rect 172518 157256 172574 157312
rect 173162 159704 173218 159760
rect 173070 158616 173126 158672
rect 173438 159840 173494 159896
rect 172426 142024 172482 142080
rect 172426 140120 172482 140176
rect 172978 147192 173034 147248
rect 173714 159840 173770 159896
rect 173990 159568 174046 159624
rect 173990 159160 174046 159216
rect 174266 159840 174322 159896
rect 174542 159874 174598 159930
rect 174174 159024 174230 159080
rect 173898 158616 173954 158672
rect 173898 146240 173954 146296
rect 174450 157800 174506 157856
rect 174358 157664 174414 157720
rect 174818 159704 174874 159760
rect 175002 159874 175058 159930
rect 174726 159568 174782 159624
rect 174818 158480 174874 158536
rect 174634 143384 174690 143440
rect 175094 159704 175150 159760
rect 175002 158480 175058 158536
rect 175370 158480 175426 158536
rect 175278 158344 175334 158400
rect 175646 158616 175702 158672
rect 175922 159840 175978 159896
rect 176106 159160 176162 159216
rect 176014 158616 176070 158672
rect 175922 158208 175978 158264
rect 176382 159704 176438 159760
rect 176934 157800 176990 157856
rect 177210 157392 177266 157448
rect 177854 157664 177910 157720
rect 177762 157392 177818 157448
rect 178130 159840 178186 159896
rect 178222 157936 178278 157992
rect 178406 157800 178462 157856
rect 178314 157392 178370 157448
rect 178682 159704 178738 159760
rect 178958 159704 179014 159760
rect 178958 157664 179014 157720
rect 179234 158616 179290 158672
rect 179234 157800 179290 157856
rect 179510 157664 179566 157720
rect 179786 158616 179842 158672
rect 180062 159840 180118 159896
rect 179970 157392 180026 157448
rect 180338 157392 180394 157448
rect 180614 159840 180670 159896
rect 180890 159568 180946 159624
rect 180890 157936 180946 157992
rect 180614 157664 180670 157720
rect 180154 136584 180210 136640
rect 181166 159840 181222 159896
rect 181442 157664 181498 157720
rect 181718 157392 181774 157448
rect 181994 158616 182050 158672
rect 181902 157936 181958 157992
rect 182270 158616 182326 158672
rect 182546 159840 182602 159896
rect 182546 159740 182548 159760
rect 182548 159740 182600 159760
rect 182600 159740 182602 159760
rect 182546 159704 182602 159740
rect 183374 159840 183430 159896
rect 183650 157392 183706 157448
rect 183926 159840 183982 159896
rect 184202 159704 184258 159760
rect 184478 159840 184534 159896
rect 185306 159840 185362 159896
rect 185030 157392 185086 157448
rect 186318 158616 186374 158672
rect 186686 158480 186742 158536
rect 186318 139576 186374 139632
rect 186318 138624 186374 138680
rect 187238 158616 187294 158672
rect 187422 159432 187478 159488
rect 187514 158616 187570 158672
rect 187790 158616 187846 158672
rect 187514 140256 187570 140312
rect 187606 140120 187662 140176
rect 187514 139576 187570 139632
rect 186686 139440 186742 139496
rect 187606 139440 187662 139496
rect 188342 159840 188398 159896
rect 188618 158616 188674 158672
rect 188894 158616 188950 158672
rect 189170 158616 189226 158672
rect 189722 159840 189778 159896
rect 189998 158616 190054 158672
rect 190274 158616 190330 158672
rect 189998 140412 190054 140448
rect 189998 140392 190000 140412
rect 190000 140392 190052 140412
rect 190052 140392 190054 140412
rect 190642 158616 190698 158672
rect 191102 159840 191158 159896
rect 190826 158344 190882 158400
rect 191378 158480 191434 158536
rect 191746 159704 191802 159760
rect 191654 157256 191710 157312
rect 191654 140800 191710 140856
rect 192022 158480 192078 158536
rect 191930 158208 191986 158264
rect 192022 157936 192078 157992
rect 192206 159840 192262 159896
rect 192206 158072 192262 158128
rect 192114 151136 192170 151192
rect 192390 158752 192446 158808
rect 192482 158480 192538 158536
rect 192758 158616 192814 158672
rect 193034 159024 193090 159080
rect 193218 158208 193274 158264
rect 193126 158072 193182 158128
rect 193586 159840 193642 159896
rect 193494 156576 193550 156632
rect 193402 151680 193458 151736
rect 193862 159840 193918 159896
rect 194138 158616 194194 158672
rect 194414 158616 194470 158672
rect 194322 158344 194378 158400
rect 194506 158480 194562 158536
rect 194690 158344 194746 158400
rect 194966 159704 195022 159760
rect 195242 159840 195298 159896
rect 195518 159840 195574 159896
rect 195794 159840 195850 159896
rect 195518 158616 195574 158672
rect 195702 155080 195758 155136
rect 195426 140256 195482 140312
rect 195426 139712 195482 139768
rect 195886 158480 195942 158536
rect 196070 158616 196126 158672
rect 196346 159704 196402 159760
rect 196622 159840 196678 159896
rect 196622 157936 196678 157992
rect 196806 158072 196862 158128
rect 197082 159160 197138 159216
rect 197266 158616 197322 158672
rect 197266 153176 197322 153232
rect 197174 151408 197230 151464
rect 196622 120808 196678 120864
rect 197542 154536 197598 154592
rect 197726 159704 197782 159760
rect 198002 159840 198058 159896
rect 198186 159568 198242 159624
rect 198278 158616 198334 158672
rect 198186 157256 198242 157312
rect 198554 159840 198610 159896
rect 198462 159568 198518 159624
rect 198370 153856 198426 153912
rect 198830 159840 198886 159896
rect 199106 159840 199162 159896
rect 198922 158888 198978 158944
rect 198646 158616 198702 158672
rect 198738 158344 198794 158400
rect 198646 139712 198702 139768
rect 198002 24112 198058 24168
rect 199382 159840 199438 159896
rect 199198 158480 199254 158536
rect 199106 158208 199162 158264
rect 199474 158616 199530 158672
rect 199474 158072 199530 158128
rect 199290 157936 199346 157992
rect 198922 148688 198978 148744
rect 199658 159704 199714 159760
rect 199842 156984 199898 157040
rect 200026 158208 200082 158264
rect 200210 159840 200266 159896
rect 200302 158480 200358 158536
rect 200210 157392 200266 157448
rect 200118 156712 200174 156768
rect 200486 158344 200542 158400
rect 200670 157392 200726 157448
rect 200394 155896 200450 155952
rect 200946 159296 201002 159352
rect 200946 158888 201002 158944
rect 201038 158616 201094 158672
rect 200946 155080 201002 155136
rect 201222 159704 201278 159760
rect 201314 158072 201370 158128
rect 201130 151544 201186 151600
rect 201498 155352 201554 155408
rect 201406 148824 201462 148880
rect 200210 143384 200266 143440
rect 201314 143384 201370 143440
rect 201314 142976 201370 143032
rect 201866 158480 201922 158536
rect 202418 159704 202474 159760
rect 202326 159024 202382 159080
rect 202142 158616 202198 158672
rect 202234 158208 202290 158264
rect 202142 157800 202198 157856
rect 202142 157528 202198 157584
rect 202050 157120 202106 157176
rect 202694 159704 202750 159760
rect 202878 159840 202934 159896
rect 202786 158208 202842 158264
rect 202786 158092 202842 158128
rect 202786 158072 202788 158092
rect 202788 158072 202840 158092
rect 202840 158072 202842 158092
rect 202786 148552 202842 148608
rect 202694 143384 202750 143440
rect 203246 159874 203302 159930
rect 203154 154128 203210 154184
rect 203522 158344 203578 158400
rect 203430 155080 203486 155136
rect 203798 158616 203854 158672
rect 203706 158072 203762 158128
rect 203614 150320 203670 150376
rect 202970 144744 203026 144800
rect 204074 159840 204130 159896
rect 203982 158888 204038 158944
rect 203982 158752 204038 158808
rect 203890 144744 203946 144800
rect 204258 159840 204314 159896
rect 204166 158480 204222 158536
rect 204074 155080 204130 155136
rect 204258 154536 204314 154592
rect 204166 152768 204222 152824
rect 204626 159704 204682 159760
rect 204534 158208 204590 158264
rect 204902 159840 204958 159896
rect 204994 158616 205050 158672
rect 205178 159840 205234 159896
rect 205086 158344 205142 158400
rect 205178 154400 205234 154456
rect 205454 159840 205510 159896
rect 205362 155488 205418 155544
rect 204718 148960 204774 149016
rect 205638 157392 205694 157448
rect 204258 91704 204314 91760
rect 206006 159160 206062 159216
rect 205914 158752 205970 158808
rect 206006 158072 206062 158128
rect 205914 154264 205970 154320
rect 206282 159840 206338 159896
rect 206558 158616 206614 158672
rect 206466 158480 206522 158536
rect 206558 158072 206614 158128
rect 206098 147600 206154 147656
rect 206466 155216 206522 155272
rect 206834 159704 206890 159760
rect 206742 159160 206798 159216
rect 206742 157528 206798 157584
rect 206650 157392 206706 157448
rect 207018 159704 207074 159760
rect 207294 159840 207350 159896
rect 207938 241304 207994 241360
rect 208214 238040 208270 238096
rect 208122 233008 208178 233064
rect 209410 238856 209466 238912
rect 207846 188264 207902 188320
rect 207938 184184 207994 184240
rect 208030 176024 208086 176080
rect 208030 168952 208086 169008
rect 207754 161200 207810 161256
rect 207386 159704 207442 159760
rect 207202 158072 207258 158128
rect 208858 164736 208914 164792
rect 206926 155216 206982 155272
rect 208122 158072 208178 158128
rect 208950 160384 209006 160440
rect 209042 158344 209098 158400
rect 208674 157936 208730 157992
rect 208490 156576 208546 156632
rect 209594 315288 209650 315344
rect 211066 319504 211122 319560
rect 210790 318008 210846 318064
rect 210238 307808 210294 307864
rect 210238 233688 210294 233744
rect 209686 224848 209742 224904
rect 209594 222808 209650 222864
rect 209502 158208 209558 158264
rect 209778 164736 209834 164792
rect 210238 161200 210294 161256
rect 210238 160248 210294 160304
rect 208674 153584 208730 153640
rect 203890 3576 203946 3632
rect 210606 240896 210662 240952
rect 210698 239536 210754 239592
rect 210698 239264 210754 239320
rect 210698 238584 210754 238640
rect 210882 315696 210938 315752
rect 210790 238176 210846 238232
rect 211066 239808 211122 239864
rect 210974 238584 211030 238640
rect 210882 235456 210938 235512
rect 211066 238176 211122 238232
rect 211066 237360 211122 237416
rect 211066 234504 211122 234560
rect 211066 233688 211122 233744
rect 210974 157664 211030 157720
rect 211986 298696 212042 298752
rect 211986 237224 212042 237280
rect 211710 155896 211766 155952
rect 219346 321680 219402 321736
rect 212906 239536 212962 239592
rect 211894 146920 211950 146976
rect 215206 319640 215262 319696
rect 213274 240352 213330 240408
rect 213090 236816 213146 236872
rect 213458 240080 213514 240136
rect 213458 239400 213514 239456
rect 212538 146240 212594 146296
rect 212538 144064 212594 144120
rect 213550 236000 213606 236056
rect 215114 316784 215170 316840
rect 214930 315832 214986 315888
rect 213642 235864 213698 235920
rect 213642 235320 213698 235376
rect 213826 236952 213882 237008
rect 213458 152224 213514 152280
rect 214194 222808 214250 222864
rect 214102 149776 214158 149832
rect 215390 236000 215446 236056
rect 215666 235184 215722 235240
rect 217874 320184 217930 320240
rect 217138 291760 217194 291816
rect 217138 240352 217194 240408
rect 216586 236680 216642 236736
rect 216586 236000 216642 236056
rect 216310 156848 216366 156904
rect 215298 149912 215354 149968
rect 214194 145832 214250 145888
rect 217414 241440 217470 241496
rect 217322 239128 217378 239184
rect 215942 144200 215998 144256
rect 216678 139848 216734 139904
rect 218978 308352 219034 308408
rect 218702 292168 218758 292224
rect 218978 240760 219034 240816
rect 218978 240352 219034 240408
rect 218518 209616 218574 209672
rect 218518 209072 218574 209128
rect 217598 152360 217654 152416
rect 218794 236816 218850 236872
rect 218058 145968 218114 146024
rect 219346 241304 219402 241360
rect 220174 306992 220230 307048
rect 220266 291896 220322 291952
rect 220358 240896 220414 240952
rect 222106 374040 222162 374096
rect 222014 369824 222070 369880
rect 221646 305632 221702 305688
rect 220726 291624 220782 291680
rect 220726 290300 220728 290320
rect 220728 290300 220780 290320
rect 220780 290300 220782 290320
rect 220726 290264 220782 290300
rect 220910 285132 220912 285152
rect 220912 285132 220964 285152
rect 220964 285132 220966 285152
rect 220910 285096 220966 285132
rect 221554 285096 221610 285152
rect 220910 276684 220966 276720
rect 220910 276664 220912 276684
rect 220912 276664 220964 276684
rect 220964 276664 220966 276684
rect 220818 240624 220874 240680
rect 221094 240080 221150 240136
rect 221278 240896 221334 240952
rect 219990 155624 220046 155680
rect 218058 145560 218114 145616
rect 218794 145560 218850 145616
rect 217414 144336 217470 144392
rect 221278 238176 221334 238232
rect 220726 237088 220782 237144
rect 220450 235184 220506 235240
rect 220450 155216 220506 155272
rect 221646 227024 221702 227080
rect 221462 142704 221518 142760
rect 221830 290128 221886 290184
rect 222014 276664 222070 276720
rect 222014 240080 222070 240136
rect 225602 360848 225658 360904
rect 224222 292848 224278 292904
rect 225694 359352 225750 359408
rect 224682 292848 224738 292904
rect 224590 291896 224646 291952
rect 224406 291624 224462 291680
rect 224590 291624 224646 291680
rect 225786 330384 225842 330440
rect 225878 318688 225934 318744
rect 225878 298016 225934 298072
rect 225786 292576 225842 292632
rect 225510 291216 225566 291272
rect 226154 291216 226210 291272
rect 227074 369144 227130 369200
rect 227626 290264 227682 290320
rect 229742 368872 229798 368928
rect 228546 322224 228602 322280
rect 229926 323584 229982 323640
rect 229466 291760 229522 291816
rect 230202 318552 230258 318608
rect 230202 294616 230258 294672
rect 229926 291760 229982 291816
rect 231306 294616 231362 294672
rect 231306 294344 231362 294400
rect 226062 289584 226118 289640
rect 244278 317056 244334 317112
rect 248418 367648 248474 367704
rect 247682 363568 247738 363624
rect 246394 289584 246450 289640
rect 247038 315152 247094 315208
rect 247774 352552 247830 352608
rect 247682 289856 247738 289912
rect 248326 290672 248382 290728
rect 251822 369008 251878 369064
rect 250626 366288 250682 366344
rect 249154 291624 249210 291680
rect 249706 290672 249762 290728
rect 251178 292032 251234 292088
rect 250810 291896 250866 291952
rect 250626 291488 250682 291544
rect 249706 290128 249762 290184
rect 251546 291352 251602 291408
rect 251178 290264 251234 290320
rect 251914 360984 251970 361040
rect 251914 291352 251970 291408
rect 251914 290400 251970 290456
rect 251822 290264 251878 290320
rect 251730 289992 251786 290048
rect 252098 290264 252154 290320
rect 248970 289720 249026 289776
rect 248142 289584 248198 289640
rect 252558 292168 252614 292224
rect 252834 290536 252890 290592
rect 253754 316920 253810 316976
rect 257066 318416 257122 318472
rect 257158 310392 257214 310448
rect 257158 309440 257214 309496
rect 259366 397976 259422 398032
rect 257894 310392 257950 310448
rect 260654 389816 260710 389872
rect 260470 388320 260526 388376
rect 259274 310392 259330 310448
rect 259274 309576 259330 309632
rect 260562 386960 260618 387016
rect 260470 322904 260526 322960
rect 262034 391176 262090 391232
rect 260654 310120 260710 310176
rect 261482 292032 261538 292088
rect 262126 302096 262182 302152
rect 262126 301552 262182 301608
rect 265622 401648 265678 401704
rect 264886 398248 264942 398304
rect 263506 391312 263562 391368
rect 263690 318144 263746 318200
rect 263690 317600 263746 317656
rect 263506 308488 263562 308544
rect 264886 317600 264942 317656
rect 264794 315988 264850 316024
rect 264794 315968 264796 315988
rect 264796 315968 264848 315988
rect 264848 315968 264850 315988
rect 266266 401920 266322 401976
rect 266174 389952 266230 390008
rect 267002 400288 267058 400344
rect 266266 307128 266322 307184
rect 270130 396888 270186 396944
rect 270038 396752 270094 396808
rect 267186 291896 267242 291952
rect 267094 290400 267150 290456
rect 247038 289448 247094 289504
rect 248050 289448 248106 289504
rect 252466 289448 252522 289504
rect 253662 289448 253718 289504
rect 237930 289312 237986 289368
rect 241242 289312 241298 289368
rect 269026 391448 269082 391504
rect 268658 390088 268714 390144
rect 268842 388456 268898 388512
rect 268750 385600 268806 385656
rect 269486 320456 269542 320512
rect 268566 315696 268622 315752
rect 268566 315152 268622 315208
rect 269578 315968 269634 316024
rect 269026 314472 269082 314528
rect 269026 313656 269082 313712
rect 267462 288496 267518 288552
rect 267554 257216 267610 257272
rect 267554 249192 267610 249248
rect 268014 250552 268070 250608
rect 267738 247560 267794 247616
rect 222014 236408 222070 236464
rect 222980 239842 223036 239898
rect 222750 239672 222806 239728
rect 223670 239828 223726 239864
rect 223670 239808 223672 239828
rect 223672 239808 223724 239828
rect 223724 239808 223726 239828
rect 223394 239708 223396 239728
rect 223396 239708 223448 239728
rect 223448 239708 223450 239728
rect 223394 239672 223450 239708
rect 223118 239400 223174 239456
rect 222014 150048 222070 150104
rect 221646 142568 221702 142624
rect 223394 238720 223450 238776
rect 223946 239672 224002 239728
rect 224038 239400 224094 239456
rect 223946 238720 224002 238776
rect 223578 220632 223634 220688
rect 223670 220088 223726 220144
rect 223118 141208 223174 141264
rect 224130 238992 224186 239048
rect 224130 238448 224186 238504
rect 224498 239400 224554 239456
rect 224406 238312 224462 238368
rect 224222 222944 224278 223000
rect 223946 184184 224002 184240
rect 224314 221584 224370 221640
rect 224774 236000 224830 236056
rect 224958 239692 225014 239728
rect 224958 239672 224960 239692
rect 224960 239672 225012 239692
rect 225012 239672 225014 239692
rect 225280 239808 225336 239864
rect 225464 239844 225466 239864
rect 225466 239844 225518 239864
rect 225518 239844 225520 239864
rect 225464 239808 225520 239844
rect 224866 235048 224922 235104
rect 224682 224848 224738 224904
rect 225234 239436 225236 239456
rect 225236 239436 225288 239456
rect 225288 239436 225290 239456
rect 225234 239400 225290 239436
rect 225050 238992 225106 239048
rect 225234 238448 225290 238504
rect 224590 219272 224646 219328
rect 225694 239672 225750 239728
rect 225786 238720 225842 238776
rect 225878 238448 225934 238504
rect 225418 218592 225474 218648
rect 224958 168952 225014 169008
rect 224314 141344 224370 141400
rect 223578 135904 223634 135960
rect 225878 238040 225934 238096
rect 226292 239808 226348 239864
rect 226430 239808 226486 239864
rect 226338 239400 226394 239456
rect 226430 239264 226486 239320
rect 226522 238992 226578 239048
rect 226890 239672 226946 239728
rect 226798 239400 226854 239456
rect 226338 238040 226394 238096
rect 226246 231512 226302 231568
rect 226338 231240 226394 231296
rect 225970 220632 226026 220688
rect 226338 145560 226394 145616
rect 226522 231104 226578 231160
rect 227120 239808 227176 239864
rect 227166 239708 227168 239728
rect 227168 239708 227220 239728
rect 227220 239708 227222 239728
rect 227166 239672 227222 239708
rect 227580 239808 227636 239864
rect 227350 239264 227406 239320
rect 227258 238584 227314 238640
rect 227350 236272 227406 236328
rect 227258 226208 227314 226264
rect 226430 138896 226486 138952
rect 227442 230968 227498 231024
rect 227626 239400 227682 239456
rect 227994 239828 228050 239864
rect 227994 239808 227996 239828
rect 227996 239808 228048 239828
rect 228048 239808 228050 239828
rect 227994 239672 228050 239728
rect 228086 238584 228142 238640
rect 227994 238312 228050 238368
rect 227718 231376 227774 231432
rect 227626 218728 227682 218784
rect 227350 158072 227406 158128
rect 227258 147056 227314 147112
rect 228178 238448 228234 238504
rect 228960 239808 229016 239864
rect 228454 238856 228510 238912
rect 228454 237224 228510 237280
rect 228270 229744 228326 229800
rect 228086 224168 228142 224224
rect 228730 239672 228786 239728
rect 228730 239400 228786 239456
rect 228730 238856 228786 238912
rect 229006 238448 229062 238504
rect 229282 239128 229338 239184
rect 229098 237632 229154 237688
rect 228822 231784 228878 231840
rect 229006 231240 229062 231296
rect 228546 224168 228602 224224
rect 228454 220224 228510 220280
rect 227166 137944 227222 138000
rect 226430 130328 226486 130384
rect 228638 144472 228694 144528
rect 229696 239808 229752 239864
rect 229650 239400 229706 239456
rect 229834 238584 229890 238640
rect 230340 239808 230396 239864
rect 230616 239808 230672 239864
rect 230156 239672 230212 239728
rect 230110 239128 230166 239184
rect 229558 237496 229614 237552
rect 229834 235592 229890 235648
rect 229558 229880 229614 229936
rect 229650 217912 229706 217968
rect 229650 217640 229706 217696
rect 229282 216960 229338 217016
rect 229006 124072 229062 124128
rect 229006 122848 229062 122904
rect 229926 220224 229982 220280
rect 230892 239808 230948 239864
rect 230662 238584 230718 238640
rect 230478 237360 230534 237416
rect 230386 217912 230442 217968
rect 230938 239672 230994 239728
rect 230846 231784 230902 231840
rect 230478 217096 230534 217152
rect 230202 214512 230258 214568
rect 230110 160520 230166 160576
rect 231122 239708 231124 239728
rect 231124 239708 231176 239728
rect 231176 239708 231178 239728
rect 231122 239672 231178 239708
rect 231030 238312 231086 238368
rect 231214 239400 231270 239456
rect 231398 239692 231454 239728
rect 231398 239672 231400 239692
rect 231400 239672 231452 239692
rect 231452 239672 231454 239692
rect 231306 238584 231362 238640
rect 231214 237496 231270 237552
rect 231996 239808 232052 239864
rect 231858 239708 231860 239728
rect 231860 239708 231912 239728
rect 231912 239708 231914 239728
rect 231858 239672 231914 239708
rect 231950 239400 232006 239456
rect 232042 239128 232098 239184
rect 231674 238076 231676 238096
rect 231676 238076 231728 238096
rect 231728 238076 231730 238096
rect 231674 238040 231730 238076
rect 231582 237904 231638 237960
rect 230846 217776 230902 217832
rect 231214 221720 231270 221776
rect 231858 234096 231914 234152
rect 233192 239808 233248 239864
rect 233514 239828 233570 239864
rect 233514 239808 233516 239828
rect 233516 239808 233568 239828
rect 233568 239808 233570 239828
rect 233790 239828 233846 239864
rect 233790 239808 233792 239828
rect 233792 239808 233844 239828
rect 233844 239808 233846 239828
rect 232686 238312 232742 238368
rect 231950 217504 232006 217560
rect 231398 217368 231454 217424
rect 231306 188264 231362 188320
rect 229926 139984 229982 140040
rect 230478 122848 230534 122904
rect 232594 147192 232650 147248
rect 232778 226208 232834 226264
rect 233238 239692 233294 239728
rect 233238 239672 233240 239692
rect 233240 239672 233292 239692
rect 233292 239672 233294 239692
rect 233146 239436 233148 239456
rect 233148 239436 233200 239456
rect 233200 239436 233202 239456
rect 233146 239400 233202 239436
rect 233330 239264 233386 239320
rect 233606 239672 233662 239728
rect 232686 143112 232742 143168
rect 233514 236544 233570 236600
rect 233882 239672 233938 239728
rect 234250 239828 234306 239864
rect 234250 239808 234252 239828
rect 234252 239808 234304 239828
rect 234304 239808 234306 239828
rect 233974 239264 234030 239320
rect 233790 235456 233846 235512
rect 233882 232600 233938 232656
rect 233790 221448 233846 221504
rect 233054 217232 233110 217288
rect 232778 141616 232834 141672
rect 234480 239842 234536 239898
rect 234250 239264 234306 239320
rect 234066 231104 234122 231160
rect 234618 239708 234620 239728
rect 234620 239708 234672 239728
rect 234672 239708 234674 239728
rect 234618 239672 234674 239708
rect 234618 239400 234674 239456
rect 234434 232736 234490 232792
rect 234342 224848 234398 224904
rect 234986 237088 235042 237144
rect 235262 239400 235318 239456
rect 235446 236272 235502 236328
rect 235354 236000 235410 236056
rect 234986 213152 235042 213208
rect 234342 151136 234398 151192
rect 235354 220360 235410 220416
rect 234158 147464 234214 147520
rect 233882 126928 233938 126984
rect 233882 126248 233938 126304
rect 235998 235864 236054 235920
rect 236182 239708 236184 239728
rect 236184 239708 236236 239728
rect 236236 239708 236238 239728
rect 236182 239672 236238 239708
rect 236090 232736 236146 232792
rect 236780 239842 236836 239898
rect 236826 239708 236828 239728
rect 236828 239708 236880 239728
rect 236880 239708 236882 239728
rect 236826 239672 236882 239708
rect 236642 237632 236698 237688
rect 236734 236952 236790 237008
rect 237102 239400 237158 239456
rect 237194 238720 237250 238776
rect 237102 238448 237158 238504
rect 237608 239808 237664 239864
rect 237424 239672 237480 239728
rect 238712 239842 238768 239898
rect 237194 236680 237250 236736
rect 236826 227432 236882 227488
rect 236642 153856 236698 153912
rect 236826 155488 236882 155544
rect 235354 141480 235410 141536
rect 237470 239400 237526 239456
rect 237654 239672 237710 239728
rect 239264 239842 239320 239898
rect 238206 239672 238262 239728
rect 237746 236408 237802 236464
rect 237930 231784 237986 231840
rect 238390 239672 238446 239728
rect 238390 237768 238446 237824
rect 237470 220768 237526 220824
rect 237378 213832 237434 213888
rect 238666 239672 238722 239728
rect 238850 239420 238906 239456
rect 238850 239400 238852 239420
rect 238852 239400 238904 239420
rect 238904 239400 238906 239420
rect 238758 238720 238814 238776
rect 238482 213696 238538 213752
rect 239034 235320 239090 235376
rect 239632 239842 239688 239898
rect 239218 239672 239274 239728
rect 240276 239842 240332 239898
rect 240644 239842 240700 239898
rect 239816 239706 239872 239762
rect 239218 233960 239274 234016
rect 239678 238992 239734 239048
rect 239678 235456 239734 235512
rect 239678 235048 239734 235104
rect 238850 213016 238906 213072
rect 238758 211792 238814 211848
rect 240138 239400 240194 239456
rect 239954 236816 240010 236872
rect 239862 231240 239918 231296
rect 240322 239672 240378 239728
rect 240138 234368 240194 234424
rect 240782 239672 240838 239728
rect 239494 220088 239550 220144
rect 238206 151272 238262 151328
rect 238022 141752 238078 141808
rect 241564 239808 241620 239864
rect 241334 239436 241336 239456
rect 241336 239436 241388 239456
rect 241388 239436 241390 239456
rect 241334 239400 241390 239436
rect 241518 238992 241574 239048
rect 242116 239842 242172 239898
rect 240874 234776 240930 234832
rect 241610 237924 241666 237960
rect 241610 237904 241612 237924
rect 241612 237904 241664 237924
rect 241664 237904 241666 237924
rect 241150 235864 241206 235920
rect 239954 218048 240010 218104
rect 239954 211928 240010 211984
rect 239770 156712 239826 156768
rect 239678 152496 239734 152552
rect 239494 137264 239550 137320
rect 241702 236000 241758 236056
rect 241978 239692 242034 239728
rect 241978 239672 241980 239692
rect 241980 239672 242032 239692
rect 242032 239672 242034 239692
rect 241978 239400 242034 239456
rect 241886 235864 241942 235920
rect 241886 235728 241942 235784
rect 241978 230016 242034 230072
rect 242806 239692 242862 239728
rect 242806 239672 242808 239692
rect 242808 239672 242860 239692
rect 242860 239672 242862 239692
rect 242622 234504 242678 234560
rect 243266 235592 243322 235648
rect 243450 235048 243506 235104
rect 242254 219000 242310 219056
rect 242254 218728 242310 218784
rect 244048 239808 244104 239864
rect 244784 239808 244840 239864
rect 243450 226888 243506 226944
rect 244002 239692 244058 239728
rect 244002 239672 244004 239692
rect 244004 239672 244056 239692
rect 244056 239672 244058 239692
rect 243910 235456 243966 235512
rect 244370 239420 244426 239456
rect 244370 239400 244372 239420
rect 244372 239400 244424 239420
rect 244424 239400 244426 239420
rect 244370 238720 244426 238776
rect 244462 238584 244518 238640
rect 244186 234232 244242 234288
rect 244002 218184 244058 218240
rect 243818 218048 243874 218104
rect 243818 213288 243874 213344
rect 245888 239842 245944 239898
rect 246578 239808 246634 239864
rect 244462 230152 244518 230208
rect 245106 237632 245162 237688
rect 245198 236952 245254 237008
rect 245382 238720 245438 238776
rect 245382 238584 245438 238640
rect 244278 126248 244334 126304
rect 245566 239128 245622 239184
rect 245934 239128 245990 239184
rect 246118 239536 246174 239592
rect 246578 239672 246634 239728
rect 246394 239128 246450 239184
rect 246394 228656 246450 228712
rect 247176 239808 247232 239864
rect 247038 239536 247094 239592
rect 247314 239536 247370 239592
rect 247728 239842 247784 239898
rect 247406 239128 247462 239184
rect 247406 238720 247462 238776
rect 247498 238584 247554 238640
rect 247222 236000 247278 236056
rect 247406 236816 247462 236872
rect 247222 226072 247278 226128
rect 247774 236000 247830 236056
rect 248050 239536 248106 239592
rect 248050 238856 248106 238912
rect 247774 222808 247830 222864
rect 248556 239808 248612 239864
rect 248970 239808 249026 239864
rect 249752 239842 249808 239898
rect 248602 239536 248658 239592
rect 248510 239264 248566 239320
rect 248418 238584 248474 238640
rect 248510 237904 248566 237960
rect 248050 227296 248106 227352
rect 248050 225528 248106 225584
rect 247774 162288 247830 162344
rect 249154 239128 249210 239184
rect 248694 230016 248750 230072
rect 249706 239572 249708 239592
rect 249708 239572 249760 239592
rect 249760 239572 249762 239592
rect 249706 239536 249762 239572
rect 249706 239264 249762 239320
rect 249706 234640 249762 234696
rect 249982 237360 250038 237416
rect 250258 239400 250314 239456
rect 249430 220768 249486 220824
rect 249154 159568 249210 159624
rect 249430 210296 249486 210352
rect 247682 112376 247738 112432
rect 250534 239808 250590 239864
rect 250626 239536 250682 239592
rect 250534 238856 250590 238912
rect 250534 238720 250590 238776
rect 250718 236000 250774 236056
rect 250902 239536 250958 239592
rect 250902 238856 250958 238912
rect 250534 234096 250590 234152
rect 251960 239842 252016 239898
rect 251362 239264 251418 239320
rect 251086 232872 251142 232928
rect 251178 228656 251234 228712
rect 251546 237632 251602 237688
rect 252006 234096 252062 234152
rect 252006 232464 252062 232520
rect 252190 239264 252246 239320
rect 252190 234096 252246 234152
rect 251822 221040 251878 221096
rect 253064 239842 253120 239898
rect 252558 233028 252614 233064
rect 252558 233008 252560 233028
rect 252560 233008 252612 233028
rect 252612 233008 252614 233028
rect 252282 220360 252338 220416
rect 252834 239556 252890 239592
rect 252834 239536 252836 239556
rect 252836 239536 252888 239556
rect 252888 239536 252890 239556
rect 253248 239808 253304 239864
rect 253294 237360 253350 237416
rect 253294 237244 253350 237280
rect 253294 237224 253296 237244
rect 253296 237224 253348 237244
rect 253348 237224 253350 237244
rect 253570 239808 253626 239864
rect 253708 239808 253764 239864
rect 253478 236408 253534 236464
rect 253386 231920 253442 231976
rect 253662 231920 253718 231976
rect 253846 230424 253902 230480
rect 253386 224712 253442 224768
rect 251270 98776 251326 98832
rect 253478 222128 253534 222184
rect 253478 152632 253534 152688
rect 253294 137672 253350 137728
rect 254352 239842 254408 239898
rect 254720 239842 254776 239898
rect 254904 239842 254960 239898
rect 254398 239672 254454 239728
rect 254490 237632 254546 237688
rect 254398 237244 254454 237280
rect 254398 237224 254400 237244
rect 254400 237224 254452 237244
rect 254452 237224 254454 237244
rect 254858 239672 254914 239728
rect 254490 231648 254546 231704
rect 255548 239808 255604 239864
rect 255134 239708 255136 239728
rect 255136 239708 255188 239728
rect 255188 239708 255190 239728
rect 255134 239672 255190 239708
rect 255134 236544 255190 236600
rect 255410 239400 255466 239456
rect 255318 238992 255374 239048
rect 255134 229880 255190 229936
rect 254122 219952 254178 220008
rect 255134 214784 255190 214840
rect 255318 214648 255374 214704
rect 255502 234776 255558 234832
rect 255962 239672 256018 239728
rect 255962 239400 256018 239456
rect 255870 238992 255926 239048
rect 255778 236816 255834 236872
rect 256054 234776 256110 234832
rect 255870 234504 255926 234560
rect 256330 236952 256386 237008
rect 256514 236272 256570 236328
rect 256422 234368 256478 234424
rect 257204 239844 257206 239864
rect 257206 239844 257258 239864
rect 257258 239844 257260 239864
rect 257204 239808 257260 239844
rect 256514 220224 256570 220280
rect 256238 163512 256294 163568
rect 256146 150184 256202 150240
rect 254582 137808 254638 137864
rect 256882 239400 256938 239456
rect 256882 238584 256938 238640
rect 257066 239672 257122 239728
rect 257250 239672 257306 239728
rect 258124 239842 258180 239898
rect 258308 239808 258364 239864
rect 258584 239808 258640 239864
rect 258768 239808 258824 239864
rect 257802 239672 257858 239728
rect 257710 233416 257766 233472
rect 256974 224168 257030 224224
rect 257526 221720 257582 221776
rect 257526 210432 257582 210488
rect 258078 238720 258134 238776
rect 258262 233824 258318 233880
rect 258170 231648 258226 231704
rect 258538 239400 258594 239456
rect 258722 239400 258778 239456
rect 258630 238584 258686 238640
rect 258630 238312 258686 238368
rect 258630 238176 258686 238232
rect 258630 237632 258686 237688
rect 258630 237360 258686 237416
rect 258078 215464 258134 215520
rect 258814 238720 258870 238776
rect 258906 238176 258962 238232
rect 258722 225936 258778 225992
rect 259504 239842 259560 239898
rect 259642 239672 259698 239728
rect 259458 236272 259514 236328
rect 259550 235320 259606 235376
rect 259550 234912 259606 234968
rect 259918 239400 259974 239456
rect 259734 237768 259790 237824
rect 259734 235320 259790 235376
rect 260286 237768 260342 237824
rect 260792 239808 260848 239864
rect 261160 239842 261216 239898
rect 260378 237360 260434 237416
rect 259090 226344 259146 226400
rect 257618 151408 257674 151464
rect 258814 215328 258870 215384
rect 259366 216552 259422 216608
rect 259366 215464 259422 215520
rect 258998 162152 259054 162208
rect 259090 161064 259146 161120
rect 258906 160928 258962 160984
rect 260102 159296 260158 159352
rect 258722 139168 258778 139224
rect 255318 127608 255374 127664
rect 258722 124752 258778 124808
rect 260378 223488 260434 223544
rect 260838 239692 260894 239728
rect 260838 239672 260840 239692
rect 260840 239672 260892 239692
rect 260892 239672 260894 239692
rect 260746 237360 260802 237416
rect 261528 239808 261584 239864
rect 262034 239808 262090 239864
rect 261022 236816 261078 236872
rect 261574 233552 261630 233608
rect 261482 229744 261538 229800
rect 260378 207576 260434 207632
rect 261482 176024 261538 176080
rect 260838 142180 260894 142216
rect 260838 142160 260840 142180
rect 260840 142160 260892 142180
rect 260892 142160 260894 142180
rect 262218 239692 262274 239728
rect 262218 239672 262220 239692
rect 262220 239672 262272 239692
rect 262272 239672 262274 239692
rect 262218 239400 262274 239456
rect 262126 239128 262182 239184
rect 261942 236544 261998 236600
rect 261758 231532 261814 231568
rect 261758 231512 261760 231532
rect 261760 231512 261812 231532
rect 261812 231512 261814 231532
rect 262632 239808 262688 239864
rect 262678 239672 262734 239728
rect 263092 239808 263148 239864
rect 263322 239808 263378 239864
rect 263552 239842 263608 239898
rect 262770 239400 262826 239456
rect 262494 236952 262550 237008
rect 262954 238856 263010 238912
rect 262954 238756 262956 238776
rect 262956 238756 263008 238776
rect 263008 238756 263010 238776
rect 262954 238720 263010 238756
rect 262218 223488 262274 223544
rect 263138 233008 263194 233064
rect 263138 223216 263194 223272
rect 263322 223488 263378 223544
rect 263322 223080 263378 223136
rect 263690 237088 263746 237144
rect 264472 239808 264528 239864
rect 264242 239264 264298 239320
rect 264426 238992 264482 239048
rect 263966 238584 264022 238640
rect 263874 238448 263930 238504
rect 263966 238040 264022 238096
rect 263874 233688 263930 233744
rect 264518 238584 264574 238640
rect 264242 230424 264298 230480
rect 264150 230152 264206 230208
rect 265392 239808 265448 239864
rect 265760 239808 265816 239864
rect 266036 239842 266092 239898
rect 264978 238992 265034 239048
rect 264978 238756 264980 238776
rect 264980 238756 265032 238776
rect 265032 238756 265034 238776
rect 264978 238720 265034 238756
rect 264886 237768 264942 237824
rect 266588 239808 266644 239864
rect 265438 238992 265494 239048
rect 265254 238584 265310 238640
rect 265714 239264 265770 239320
rect 265530 238720 265586 238776
rect 264702 227432 264758 227488
rect 264610 227160 264666 227216
rect 263690 170312 263746 170368
rect 263598 167592 263654 167648
rect 263138 161880 263194 161936
rect 265070 165008 265126 165064
rect 264426 164872 264482 164928
rect 264242 161200 264298 161256
rect 263046 159024 263102 159080
rect 262954 154128 263010 154184
rect 262862 152768 262918 152824
rect 263598 142860 263654 142896
rect 263598 142840 263600 142860
rect 263600 142840 263652 142860
rect 263652 142840 263654 142860
rect 265806 238720 265862 238776
rect 266634 239708 266636 239728
rect 266636 239708 266688 239728
rect 266688 239708 266690 239728
rect 266082 239264 266138 239320
rect 265898 238312 265954 238368
rect 265806 237904 265862 237960
rect 265714 237224 265770 237280
rect 265714 228792 265770 228848
rect 265714 179968 265770 180024
rect 266358 235184 266414 235240
rect 266634 239672 266690 239708
rect 266634 239436 266636 239456
rect 266636 239436 266688 239456
rect 266688 239436 266690 239456
rect 266634 239400 266690 239436
rect 266910 238448 266966 238504
rect 267278 239264 267334 239320
rect 267646 239808 267702 239864
rect 267462 235864 267518 235920
rect 267094 231240 267150 231296
rect 266726 228928 266782 228984
rect 267002 228928 267058 228984
rect 266726 174528 266782 174584
rect 266082 166232 266138 166288
rect 265898 163376 265954 163432
rect 265622 161336 265678 161392
rect 267186 227432 267242 227488
rect 267186 204856 267242 204912
rect 267462 182824 267518 182880
rect 267094 171672 267150 171728
rect 268106 240352 268162 240408
rect 267646 162016 267702 162072
rect 267002 159160 267058 159216
rect 265622 122168 265678 122224
rect 267922 235184 267978 235240
rect 268014 234776 268070 234832
rect 268382 238720 268438 238776
rect 268842 247832 268898 247888
rect 268658 243072 268714 243128
rect 268658 242936 268714 242992
rect 268658 240080 268714 240136
rect 268290 237496 268346 237552
rect 268658 238040 268714 238096
rect 268474 234912 268530 234968
rect 268934 237360 268990 237416
rect 269118 247696 269174 247752
rect 269210 240624 269266 240680
rect 269210 240352 269266 240408
rect 268750 234232 268806 234288
rect 268658 232872 268714 232928
rect 268566 231240 268622 231296
rect 268014 158888 268070 158944
rect 269670 308624 269726 308680
rect 269578 239536 269634 239592
rect 269394 237360 269450 237416
rect 269578 237360 269634 237416
rect 269854 317328 269910 317384
rect 269854 315696 269910 315752
rect 270038 320456 270094 320512
rect 270222 396616 270278 396672
rect 271234 395256 271290 395312
rect 270406 394032 270462 394088
rect 270130 311616 270186 311672
rect 270038 240760 270094 240816
rect 271142 320320 271198 320376
rect 271050 315832 271106 315888
rect 270406 310256 270462 310312
rect 270222 257488 270278 257544
rect 270222 241576 270278 241632
rect 270406 246336 270462 246392
rect 270498 240080 270554 240136
rect 270406 238312 270462 238368
rect 270314 238176 270370 238232
rect 269946 234504 270002 234560
rect 270130 233960 270186 234016
rect 269762 226208 269818 226264
rect 269210 160792 269266 160848
rect 269118 148688 269174 148744
rect 269762 148552 269818 148608
rect 270590 237904 270646 237960
rect 270774 245384 270830 245440
rect 270866 240760 270922 240816
rect 270866 238992 270922 239048
rect 270866 238176 270922 238232
rect 270774 236680 270830 236736
rect 270682 231784 270738 231840
rect 270590 156984 270646 157040
rect 271418 317192 271474 317248
rect 271602 314472 271658 314528
rect 271602 313792 271658 313848
rect 274178 397024 274234 397080
rect 272890 395528 272946 395584
rect 271786 395392 271842 395448
rect 271694 311752 271750 311808
rect 271694 241576 271750 241632
rect 271234 239264 271290 239320
rect 271694 237360 271750 237416
rect 270866 158752 270922 158808
rect 270774 155080 270830 155136
rect 271786 234368 271842 234424
rect 272614 318280 272670 318336
rect 272154 243752 272210 243808
rect 272154 236680 272210 236736
rect 272154 236408 272210 236464
rect 272338 242528 272394 242584
rect 272338 236272 272394 236328
rect 272890 319232 272946 319288
rect 273718 393896 273774 393952
rect 272706 288632 272762 288688
rect 272062 142296 272118 142352
rect 272982 236680 273038 236736
rect 273626 315832 273682 315888
rect 273902 387232 273958 387288
rect 273902 320592 273958 320648
rect 273350 152904 273406 152960
rect 272246 136604 272302 136640
rect 272246 136584 272248 136604
rect 272248 136584 272300 136604
rect 272300 136584 272302 136604
rect 274086 314336 274142 314392
rect 280066 454008 280122 454064
rect 278318 448568 278374 448624
rect 275098 320728 275154 320784
rect 274454 317056 274510 317112
rect 274546 241984 274602 242040
rect 274546 241884 274548 241904
rect 274548 241884 274600 241904
rect 274600 241884 274602 241904
rect 274546 241848 274602 241884
rect 274454 232736 274510 232792
rect 274914 239128 274970 239184
rect 274638 148824 274694 148880
rect 275374 320728 275430 320784
rect 275558 239944 275614 240000
rect 276018 368600 276074 368656
rect 276478 368600 276534 368656
rect 275926 314608 275982 314664
rect 274914 157120 274970 157176
rect 276110 154400 276166 154456
rect 276662 322088 276718 322144
rect 276754 321000 276810 321056
rect 278042 390224 278098 390280
rect 277766 371728 277822 371784
rect 277858 320864 277914 320920
rect 277858 320184 277914 320240
rect 277306 318824 277362 318880
rect 276754 315288 276810 315344
rect 277122 245112 277178 245168
rect 277306 231376 277362 231432
rect 278042 361664 278098 361720
rect 278318 373380 278374 373416
rect 278318 373360 278320 373380
rect 278320 373360 278372 373380
rect 278372 373360 278374 373380
rect 278318 371728 278374 371784
rect 278226 320592 278282 320648
rect 278226 320184 278282 320240
rect 278318 319504 278374 319560
rect 278410 318960 278466 319016
rect 278318 318824 278374 318880
rect 278318 317464 278374 317520
rect 277490 160656 277546 160712
rect 276294 153040 276350 153096
rect 273626 3440 273682 3496
rect 279238 321816 279294 321872
rect 279238 321544 279294 321600
rect 278778 243752 278834 243808
rect 278778 242936 278834 242992
rect 278686 233960 278742 234016
rect 279514 321272 279570 321328
rect 279698 318824 279754 318880
rect 279606 318552 279662 318608
rect 279606 317464 279662 317520
rect 279882 361800 279938 361856
rect 280618 451968 280674 452024
rect 280618 372000 280674 372056
rect 280066 371864 280122 371920
rect 278870 144744 278926 144800
rect 280158 320728 280214 320784
rect 280894 451560 280950 451616
rect 280802 373904 280858 373960
rect 280894 373224 280950 373280
rect 280802 372952 280858 373008
rect 281078 316104 281134 316160
rect 282826 451696 282882 451752
rect 282182 448704 282238 448760
rect 281170 245248 281226 245304
rect 281630 319912 281686 319968
rect 281998 363568 282054 363624
rect 282182 361664 282238 361720
rect 282090 322904 282146 322960
rect 281906 322088 281962 322144
rect 281998 321680 282054 321736
rect 281998 321136 282054 321192
rect 281998 320592 282054 320648
rect 281814 319640 281870 319696
rect 281538 240216 281594 240272
rect 285954 448840 286010 448896
rect 282918 391992 282974 392048
rect 282826 371320 282882 371376
rect 284114 373904 284170 373960
rect 284206 373224 284262 373280
rect 284114 371592 284170 371648
rect 285080 369824 285136 369880
rect 290462 447888 290518 447944
rect 286322 447752 286378 447808
rect 286046 372680 286102 372736
rect 285954 369960 286010 370016
rect 286414 370096 286470 370152
rect 286184 369688 286240 369744
rect 289082 376760 289138 376816
rect 287150 374448 287206 374504
rect 287702 374448 287758 374504
rect 287150 374040 287206 374096
rect 287058 369960 287114 370016
rect 286920 369688 286976 369744
rect 287058 369688 287114 369744
rect 284482 369416 284538 369472
rect 286782 369416 286838 369472
rect 287794 371864 287850 371920
rect 288254 371456 288310 371512
rect 291842 443536 291898 443592
rect 289726 372136 289782 372192
rect 290002 371728 290058 371784
rect 289726 371320 289782 371376
rect 287288 369416 287344 369472
rect 295338 397160 295394 397216
rect 297546 401240 297602 401296
rect 300214 449112 300270 449168
rect 300398 400968 300454 401024
rect 301594 399744 301650 399800
rect 308402 454144 308458 454200
rect 304262 439456 304318 439512
rect 303526 401104 303582 401160
rect 303618 384240 303674 384296
rect 305734 399608 305790 399664
rect 303480 369688 303536 369744
rect 303986 369688 304042 369744
rect 307666 449928 307722 449984
rect 307666 404232 307722 404288
rect 309138 450472 309194 450528
rect 309598 375400 309654 375456
rect 308770 371456 308826 371512
rect 309874 450064 309930 450120
rect 310058 375400 310114 375456
rect 312542 448976 312598 449032
rect 311254 401512 311310 401568
rect 310518 372544 310574 372600
rect 310242 371728 310298 371784
rect 311346 372544 311402 372600
rect 306286 369416 306342 369472
rect 307666 369416 307722 369472
rect 311806 369416 311862 369472
rect 312312 369416 312368 369472
rect 313186 370096 313242 370152
rect 314106 400832 314162 400888
rect 315394 399880 315450 399936
rect 317694 385736 317750 385792
rect 315854 369824 315910 369880
rect 319442 369824 319498 369880
rect 319810 369552 319866 369608
rect 322478 399472 322534 399528
rect 331494 449520 331550 449576
rect 331494 448704 331550 448760
rect 314382 369416 314438 369472
rect 318430 369416 318486 369472
rect 319902 369416 319958 369472
rect 321374 369416 321430 369472
rect 322846 369416 322902 369472
rect 288024 369280 288080 369336
rect 289128 369280 289184 369336
rect 312312 369280 312368 369336
rect 327722 360848 327778 360904
rect 327722 359352 327778 359408
rect 327446 355272 327502 355328
rect 282458 352552 282514 352608
rect 327538 330384 327594 330440
rect 282366 321544 282422 321600
rect 282458 321408 282514 321464
rect 282458 321000 282514 321056
rect 282688 320728 282744 320784
rect 283976 320728 284032 320784
rect 284344 320728 284400 320784
rect 285540 320728 285596 320784
rect 288392 320728 288448 320784
rect 289128 320728 289184 320784
rect 289312 320728 289368 320784
rect 289864 320728 289920 320784
rect 291428 320728 291484 320784
rect 295384 320728 295440 320784
rect 297040 320728 297096 320784
rect 301272 320728 301328 320784
rect 304032 320728 304088 320784
rect 304768 320728 304824 320784
rect 307528 320728 307584 320784
rect 311116 320728 311172 320784
rect 314796 320748 314852 320784
rect 314796 320728 314798 320748
rect 314798 320728 314850 320748
rect 314850 320728 314852 320748
rect 315808 320728 315864 320784
rect 318476 320728 318532 320784
rect 321696 320728 321752 320784
rect 322432 320728 322488 320784
rect 324088 320728 324144 320784
rect 324640 320728 324696 320784
rect 325192 320728 325248 320784
rect 326480 320728 326536 320784
rect 327400 320728 327456 320784
rect 284712 320592 284768 320648
rect 285080 320592 285136 320648
rect 288300 320592 288356 320648
rect 292164 320592 292220 320648
rect 293452 320592 293508 320648
rect 294096 320592 294152 320648
rect 298144 320592 298200 320648
rect 298512 320592 298568 320648
rect 299248 320592 299304 320648
rect 304492 320592 304548 320648
rect 305320 320592 305376 320648
rect 307620 320612 307676 320648
rect 307620 320592 307622 320612
rect 307622 320592 307674 320612
rect 307674 320592 307676 320612
rect 313784 320592 313840 320648
rect 317832 320592 317888 320648
rect 326756 320592 326812 320648
rect 327308 320592 327364 320648
rect 299984 320456 300040 320512
rect 300536 320456 300592 320512
rect 302100 320456 302156 320512
rect 305504 320456 305560 320512
rect 312588 320456 312644 320512
rect 313508 320456 313564 320512
rect 319672 320456 319728 320512
rect 322984 320456 323040 320512
rect 324364 320456 324420 320512
rect 325008 320456 325064 320512
rect 308724 320320 308780 320376
rect 309460 320320 309516 320376
rect 310932 320320 310988 320376
rect 311484 320320 311540 320376
rect 323536 320320 323592 320376
rect 325468 320320 325524 320376
rect 326296 320320 326352 320376
rect 284528 320184 284584 320240
rect 284896 320184 284952 320240
rect 285448 320184 285504 320240
rect 286828 320184 286884 320240
rect 287288 320184 287344 320240
rect 288024 320184 288080 320240
rect 290324 320184 290380 320240
rect 291980 320184 292036 320240
rect 292440 320184 292496 320240
rect 293728 320184 293784 320240
rect 294280 320184 294336 320240
rect 294648 320184 294704 320240
rect 295016 320184 295072 320240
rect 296028 320184 296084 320240
rect 296488 320184 296544 320240
rect 296948 320184 297004 320240
rect 298696 320184 298752 320240
rect 299156 320184 299212 320240
rect 300168 320184 300224 320240
rect 302744 320184 302800 320240
rect 305136 320184 305192 320240
rect 306240 320184 306296 320240
rect 307068 320184 307124 320240
rect 308448 320184 308504 320240
rect 308632 320184 308688 320240
rect 309644 320184 309700 320240
rect 312496 320184 312552 320240
rect 314152 320184 314208 320240
rect 314980 320184 315036 320240
rect 316912 320184 316968 320240
rect 319120 320184 319176 320240
rect 319856 320184 319912 320240
rect 320592 320184 320648 320240
rect 282872 320048 282928 320104
rect 282504 319776 282560 319832
rect 283332 320048 283388 320104
rect 282918 319232 282974 319288
rect 282642 317736 282698 317792
rect 282366 316784 282422 316840
rect 277122 3304 277178 3360
rect 280710 6024 280766 6080
rect 282458 240216 282514 240272
rect 283102 319640 283158 319696
rect 283010 307672 283066 307728
rect 283608 320048 283664 320104
rect 283792 319878 283848 319934
rect 284068 320048 284124 320104
rect 283654 319368 283710 319424
rect 283838 318960 283894 319016
rect 283562 317464 283618 317520
rect 284252 319878 284308 319934
rect 284022 319640 284078 319696
rect 284022 319368 284078 319424
rect 284298 319640 284354 319696
rect 283930 317872 283986 317928
rect 283654 314608 283710 314664
rect 283378 241304 283434 241360
rect 283010 230288 283066 230344
rect 282458 148960 282514 149016
rect 282458 148280 282514 148336
rect 283746 310528 283802 310584
rect 283930 305768 283986 305824
rect 283930 298968 283986 299024
rect 284298 318416 284354 318472
rect 284482 319232 284538 319288
rect 284390 317328 284446 317384
rect 284114 316648 284170 316704
rect 284758 318960 284814 319016
rect 284666 317600 284722 317656
rect 284022 295024 284078 295080
rect 285632 320048 285688 320104
rect 285034 318960 285090 319016
rect 285586 319776 285642 319832
rect 284942 317464 284998 317520
rect 284850 315968 284906 316024
rect 285126 317464 285182 317520
rect 284298 241032 284354 241088
rect 284022 151680 284078 151736
rect 284022 151136 284078 151192
rect 285770 319776 285826 319832
rect 286276 320048 286332 320104
rect 286184 319776 286240 319832
rect 286460 319878 286516 319934
rect 285402 297064 285458 297120
rect 285678 309304 285734 309360
rect 286230 318280 286286 318336
rect 286230 317600 286286 317656
rect 286138 310120 286194 310176
rect 285494 242664 285550 242720
rect 285586 241168 285642 241224
rect 286920 320048 286976 320104
rect 286506 318688 286562 318744
rect 286782 319640 286838 319696
rect 286506 317600 286562 317656
rect 286230 242800 286286 242856
rect 285402 222672 285458 222728
rect 284942 217776 284998 217832
rect 284482 151544 284538 151600
rect 284482 151000 284538 151056
rect 284298 6840 284354 6896
rect 286414 298016 286470 298072
rect 286414 296928 286470 296984
rect 287196 320048 287252 320104
rect 287058 319232 287114 319288
rect 287242 319776 287298 319832
rect 287472 320048 287528 320104
rect 287242 319096 287298 319152
rect 287242 318960 287298 319016
rect 287426 319640 287482 319696
rect 287334 318008 287390 318064
rect 287334 317636 287336 317656
rect 287336 317636 287388 317656
rect 287388 317636 287390 317656
rect 287334 317600 287390 317636
rect 286782 298016 286838 298072
rect 286782 297608 286838 297664
rect 287334 302096 287390 302152
rect 287840 320048 287896 320104
rect 287610 319640 287666 319696
rect 287610 318008 287666 318064
rect 288116 320048 288172 320104
rect 288484 320048 288540 320104
rect 288668 320048 288724 320104
rect 287932 319776 287988 319832
rect 287978 319640 288034 319696
rect 287702 313792 287758 313848
rect 287610 295976 287666 296032
rect 287518 233824 287574 233880
rect 286782 221856 286838 221912
rect 288070 319232 288126 319288
rect 287978 317872 288034 317928
rect 287886 309576 287942 309632
rect 287702 229880 287758 229936
rect 288346 318688 288402 318744
rect 288622 319776 288678 319832
rect 288530 319640 288586 319696
rect 288254 309440 288310 309496
rect 288070 298152 288126 298208
rect 288438 317056 288494 317112
rect 288346 296248 288402 296304
rect 288346 236544 288402 236600
rect 288944 319878 289000 319934
rect 289220 320048 289276 320104
rect 289174 319776 289230 319832
rect 288898 319232 288954 319288
rect 289082 319232 289138 319288
rect 289082 318552 289138 318608
rect 288806 298832 288862 298888
rect 288714 296112 288770 296168
rect 288622 294888 288678 294944
rect 289174 317872 289230 317928
rect 289772 320048 289828 320104
rect 289818 319776 289874 319832
rect 290416 320048 290472 320104
rect 289542 318144 289598 318200
rect 289726 318960 289782 319016
rect 288530 238992 288586 239048
rect 288438 217912 288494 217968
rect 289358 310392 289414 310448
rect 289450 297200 289506 297256
rect 289358 222944 289414 223000
rect 289818 318280 289874 318336
rect 290692 320048 290748 320104
rect 290968 320048 291024 320104
rect 291152 320048 291208 320104
rect 290600 319776 290656 319832
rect 290370 319640 290426 319696
rect 290186 311208 290242 311264
rect 290002 298968 290058 299024
rect 289910 294752 289966 294808
rect 289726 294616 289782 294672
rect 290738 319640 290794 319696
rect 290554 318008 290610 318064
rect 290462 310392 290518 310448
rect 289450 221720 289506 221776
rect 290554 294752 290610 294808
rect 291106 319776 291162 319832
rect 291704 320048 291760 320104
rect 290922 318008 290978 318064
rect 291106 311344 291162 311400
rect 291106 311208 291162 311264
rect 290738 295024 290794 295080
rect 290646 229744 290702 229800
rect 290554 216280 290610 216336
rect 291750 318960 291806 319016
rect 291842 309712 291898 309768
rect 291014 294480 291070 294536
rect 290738 216416 290794 216472
rect 290646 157256 290702 157312
rect 291106 157256 291162 157312
rect 291106 156576 291162 156632
rect 291382 6704 291438 6760
rect 292118 319368 292174 319424
rect 292302 319776 292358 319832
rect 292532 319776 292588 319832
rect 292808 320048 292864 320104
rect 292578 319540 292580 319560
rect 292580 319540 292632 319560
rect 292632 319540 292634 319560
rect 292578 319504 292634 319540
rect 292486 318960 292542 319016
rect 292670 319232 292726 319288
rect 292670 318960 292726 319016
rect 292026 311752 292082 311808
rect 292210 295160 292266 295216
rect 292026 228384 292082 228440
rect 293084 320048 293140 320104
rect 293038 319368 293094 319424
rect 292946 319252 293002 319288
rect 292946 319232 292948 319252
rect 292948 319232 293000 319252
rect 293000 319232 293002 319252
rect 292762 313656 292818 313712
rect 293222 314336 293278 314392
rect 293406 318008 293462 318064
rect 293682 318960 293738 319016
rect 294004 320048 294060 320104
rect 294234 319776 294290 319832
rect 294234 319232 294290 319288
rect 292854 299240 292910 299296
rect 292854 298696 292910 298752
rect 294510 319368 294566 319424
rect 294602 318688 294658 318744
rect 294970 319640 295026 319696
rect 294694 312568 294750 312624
rect 294050 236952 294106 237008
rect 294050 236000 294106 236056
rect 294878 305768 294934 305824
rect 295062 236000 295118 236056
rect 295844 320048 295900 320104
rect 296212 320048 296268 320104
rect 295338 310528 295394 310584
rect 295798 319368 295854 319424
rect 296074 319232 296130 319288
rect 295706 318960 295762 319016
rect 295798 318552 295854 318608
rect 296258 305904 296314 305960
rect 296166 302096 296222 302152
rect 296074 238856 296130 238912
rect 295338 147600 295394 147656
rect 295338 146920 295394 146976
rect 292578 125432 292634 125488
rect 293222 125432 293278 125488
rect 292578 124752 292634 124808
rect 294878 6568 294934 6624
rect 297224 320048 297280 320104
rect 296718 319232 296774 319288
rect 296626 316648 296682 316704
rect 296534 312432 296590 312488
rect 296902 319232 296958 319288
rect 296902 318824 296958 318880
rect 297592 320048 297648 320104
rect 297776 320048 297832 320104
rect 297454 319232 297510 319288
rect 297362 318960 297418 319016
rect 297362 318552 297418 318608
rect 297362 318144 297418 318200
rect 297730 319368 297786 319424
rect 297546 318960 297602 319016
rect 297730 318960 297786 319016
rect 297546 318416 297602 318472
rect 296626 231512 296682 231568
rect 296350 227160 296406 227216
rect 296166 218592 296222 218648
rect 296074 146920 296130 146976
rect 297730 306176 297786 306232
rect 298420 320048 298476 320104
rect 299064 320048 299120 320104
rect 298742 318960 298798 319016
rect 298650 316512 298706 316568
rect 298374 316376 298430 316432
rect 297914 293256 297970 293312
rect 298190 237088 298246 237144
rect 298558 316240 298614 316296
rect 298374 297472 298430 297528
rect 299110 309712 299166 309768
rect 298926 298832 298982 298888
rect 298834 237088 298890 237144
rect 299432 320048 299488 320104
rect 300076 320048 300132 320104
rect 300260 320048 300316 320104
rect 299386 318960 299442 319016
rect 299294 315968 299350 316024
rect 299202 302096 299258 302152
rect 299662 318844 299718 318880
rect 299662 318824 299664 318844
rect 299664 318824 299716 318844
rect 299716 318824 299718 318844
rect 299478 316104 299534 316160
rect 299478 313928 299534 313984
rect 299938 319368 299994 319424
rect 299386 299376 299442 299432
rect 300214 318996 300216 319016
rect 300216 318996 300268 319016
rect 300268 318996 300270 319016
rect 300214 318960 300270 318996
rect 300122 318824 300178 318880
rect 300214 318008 300270 318064
rect 300122 317464 300178 317520
rect 300490 319368 300546 319424
rect 300030 302776 300086 302832
rect 298926 222808 298982 222864
rect 298190 150320 298246 150376
rect 299386 150320 299442 150376
rect 299386 149640 299442 149696
rect 300904 320048 300960 320104
rect 300582 318688 300638 318744
rect 300582 317736 300638 317792
rect 301502 319368 301558 319424
rect 301410 317464 301466 317520
rect 301410 308760 301466 308816
rect 301410 308352 301466 308408
rect 300766 301552 300822 301608
rect 300582 293120 300638 293176
rect 301686 318960 301742 319016
rect 301778 317464 301834 317520
rect 302054 317736 302110 317792
rect 302836 320048 302892 320104
rect 302238 318416 302294 318472
rect 302606 317464 302662 317520
rect 302790 318144 302846 318200
rect 301870 302776 301926 302832
rect 303664 320048 303720 320104
rect 303158 317464 303214 317520
rect 302146 238176 302202 238232
rect 303342 317736 303398 317792
rect 303802 317872 303858 317928
rect 304262 317736 304318 317792
rect 303250 289312 303306 289368
rect 304538 307400 304594 307456
rect 305182 319504 305238 319560
rect 305872 320048 305928 320104
rect 305366 302912 305422 302968
rect 305550 318960 305606 319016
rect 305734 319504 305790 319560
rect 306102 319504 306158 319560
rect 306194 317736 306250 317792
rect 306976 320048 307032 320104
rect 306378 318688 306434 318744
rect 306470 318416 306526 318472
rect 306378 317872 306434 317928
rect 306286 317464 306342 317520
rect 306378 314628 306434 314664
rect 306378 314608 306380 314628
rect 306380 314608 306432 314628
rect 306432 314608 306434 314628
rect 306746 319504 306802 319560
rect 306654 319368 306710 319424
rect 306838 317464 306894 317520
rect 306838 306312 306894 306368
rect 306654 303320 306710 303376
rect 306654 302232 306710 302288
rect 307344 320048 307400 320104
rect 307298 319368 307354 319424
rect 308080 320048 308136 320104
rect 307942 319504 307998 319560
rect 307942 319368 307998 319424
rect 307758 317464 307814 317520
rect 307298 306312 307354 306368
rect 307114 304952 307170 305008
rect 307114 302232 307170 302288
rect 306102 289040 306158 289096
rect 307666 304952 307722 305008
rect 307758 303592 307814 303648
rect 307574 297064 307630 297120
rect 308126 319504 308182 319560
rect 308218 318960 308274 319016
rect 308310 318280 308366 318336
rect 308494 318688 308550 318744
rect 309828 320048 309884 320104
rect 308862 317736 308918 317792
rect 309230 319504 309286 319560
rect 308678 306040 308734 306096
rect 309046 298016 309102 298072
rect 309046 297644 309048 297664
rect 309048 297644 309100 297664
rect 309100 297644 309102 297664
rect 309046 297608 309102 297644
rect 308954 297064 309010 297120
rect 310288 320048 310344 320104
rect 309782 319504 309838 319560
rect 309690 319368 309746 319424
rect 309690 318824 309746 318880
rect 309782 317464 309838 317520
rect 309966 317464 310022 317520
rect 310058 315696 310114 315752
rect 309782 313112 309838 313168
rect 309690 312296 309746 312352
rect 310518 315560 310574 315616
rect 310518 312840 310574 312896
rect 309506 305904 309562 305960
rect 308494 227296 308550 227352
rect 310058 298152 310114 298208
rect 310334 299412 310336 299432
rect 310336 299412 310388 299432
rect 310388 299412 310390 299432
rect 310334 299376 310390 299412
rect 310978 319368 311034 319424
rect 311668 320048 311724 320104
rect 311162 315560 311218 315616
rect 310518 228656 310574 228712
rect 312128 320048 312184 320104
rect 311898 317464 311954 317520
rect 312082 318960 312138 319016
rect 312772 320048 312828 320104
rect 312266 319368 312322 319424
rect 311622 298832 311678 298888
rect 311714 287680 311770 287736
rect 312910 317736 312966 317792
rect 312450 314608 312506 314664
rect 312818 314472 312874 314528
rect 312542 313112 312598 313168
rect 312358 307400 312414 307456
rect 312266 307264 312322 307320
rect 312174 306176 312230 306232
rect 311530 233688 311586 233744
rect 312726 307264 312782 307320
rect 313876 320048 313932 320104
rect 313646 318688 313702 318744
rect 313094 314608 313150 314664
rect 313830 317464 313886 317520
rect 313462 307808 313518 307864
rect 314014 319504 314070 319560
rect 314198 319368 314254 319424
rect 312634 234096 312690 234152
rect 312542 225936 312598 225992
rect 311346 224848 311402 224904
rect 311162 105440 311218 105496
rect 314014 308352 314070 308408
rect 314014 307808 314070 307864
rect 314658 318280 314714 318336
rect 314474 317464 314530 317520
rect 315532 320048 315588 320104
rect 314934 318008 314990 318064
rect 314842 317056 314898 317112
rect 314474 306992 314530 307048
rect 315302 316920 315358 316976
rect 314842 306992 314898 307048
rect 314750 305768 314806 305824
rect 315302 296792 315358 296848
rect 315486 306992 315542 307048
rect 316636 320048 316692 320104
rect 315670 304272 315726 304328
rect 315578 257352 315634 257408
rect 316682 316784 316738 316840
rect 316406 311344 316462 311400
rect 316406 310528 316462 310584
rect 317142 319504 317198 319560
rect 317142 318008 317198 318064
rect 317050 315968 317106 316024
rect 316866 297472 316922 297528
rect 316866 296792 316922 296848
rect 316774 267008 316830 267064
rect 317326 317736 317382 317792
rect 317142 312724 317198 312760
rect 317142 312704 317144 312724
rect 317144 312704 317196 312724
rect 317196 312704 317198 312724
rect 317142 310528 317198 310584
rect 317786 317736 317842 317792
rect 318292 320048 318348 320104
rect 318154 317872 318210 317928
rect 318062 317464 318118 317520
rect 317694 311616 317750 311672
rect 317510 303456 317566 303512
rect 317510 302776 317566 302832
rect 318844 320048 318900 320104
rect 319488 320048 319544 320104
rect 318706 318008 318762 318064
rect 318982 319368 319038 319424
rect 318890 318280 318946 318336
rect 318798 317872 318854 317928
rect 318890 317736 318946 317792
rect 318062 311480 318118 311536
rect 318062 310936 318118 310992
rect 316774 224576 316830 224632
rect 317418 223352 317474 223408
rect 315578 221992 315634 222048
rect 318154 260072 318210 260128
rect 319350 318552 319406 318608
rect 320040 320048 320096 320104
rect 319258 315288 319314 315344
rect 319166 314608 319222 314664
rect 320500 320048 320556 320104
rect 319626 318960 319682 319016
rect 319534 314064 319590 314120
rect 318706 300736 318762 300792
rect 318706 298832 318762 298888
rect 318706 297200 318762 297256
rect 319718 318824 319774 318880
rect 319994 318960 320050 319016
rect 319902 314608 319958 314664
rect 319902 313928 319958 313984
rect 319534 242392 319590 242448
rect 320086 318416 320142 318472
rect 320362 318688 320418 318744
rect 320270 318008 320326 318064
rect 320638 319504 320694 319560
rect 320730 318280 320786 318336
rect 321328 320048 321384 320104
rect 321098 318688 321154 318744
rect 321006 317872 321062 317928
rect 320914 317464 320970 317520
rect 321098 317464 321154 317520
rect 320822 313248 320878 313304
rect 320546 309984 320602 310040
rect 320454 304680 320510 304736
rect 320086 242528 320142 242584
rect 320914 304952 320970 305008
rect 321098 309984 321154 310040
rect 321282 304680 321338 304736
rect 321742 316648 321798 316704
rect 322018 318416 322074 318472
rect 322018 317600 322074 317656
rect 322202 317600 322258 317656
rect 321558 315152 321614 315208
rect 321558 313248 321614 313304
rect 322478 317192 322534 317248
rect 322478 316648 322534 316704
rect 322800 320048 322856 320104
rect 323352 320048 323408 320104
rect 322662 317464 322718 317520
rect 322386 316104 322442 316160
rect 322294 314608 322350 314664
rect 321742 310256 321798 310312
rect 322202 307536 322258 307592
rect 321006 253136 321062 253192
rect 320914 242120 320970 242176
rect 315302 113872 315358 113928
rect 318798 119448 318854 119504
rect 322662 314608 322718 314664
rect 322846 317872 322902 317928
rect 322662 310256 322718 310312
rect 322386 304544 322442 304600
rect 322386 258712 322442 258768
rect 322202 249056 322258 249112
rect 323122 312976 323178 313032
rect 323490 319504 323546 319560
rect 323490 317600 323546 317656
rect 324180 320048 324236 320104
rect 324456 320048 324512 320104
rect 323766 319504 323822 319560
rect 323674 316240 323730 316296
rect 323766 316104 323822 316160
rect 323122 309032 323178 309088
rect 323030 303184 323086 303240
rect 323582 313112 323638 313168
rect 323582 312704 323638 312760
rect 323674 309032 323730 309088
rect 323674 308624 323730 308680
rect 324042 318280 324098 318336
rect 324042 316376 324098 316432
rect 324226 315424 324282 315480
rect 323858 313792 323914 313848
rect 324226 313112 324282 313168
rect 324134 312976 324190 313032
rect 324134 312568 324190 312624
rect 323950 303456 324006 303512
rect 324042 303184 324098 303240
rect 323674 247560 323730 247616
rect 323582 246200 323638 246256
rect 324594 318960 324650 319016
rect 324502 318824 324558 318880
rect 324410 318588 324412 318608
rect 324412 318588 324464 318608
rect 324464 318588 324466 318608
rect 324410 318552 324466 318588
rect 324318 312432 324374 312488
rect 324916 320048 324972 320104
rect 325560 320048 325616 320104
rect 325054 318824 325110 318880
rect 324962 317872 325018 317928
rect 324594 311616 324650 311672
rect 324502 310120 324558 310176
rect 324410 308896 324466 308952
rect 325054 317328 325110 317384
rect 325330 319504 325386 319560
rect 325330 314472 325386 314528
rect 325514 318688 325570 318744
rect 325422 314336 325478 314392
rect 325146 311616 325202 311672
rect 325054 310120 325110 310176
rect 324962 309304 325018 309360
rect 325146 271088 325202 271144
rect 325054 250416 325110 250472
rect 325606 308896 325662 308952
rect 325882 318144 325938 318200
rect 325882 317872 325938 317928
rect 325882 317464 325938 317520
rect 326572 320048 326628 320104
rect 326250 317464 326306 317520
rect 326066 315832 326122 315888
rect 326940 320048 326996 320104
rect 326618 319504 326674 319560
rect 326526 317328 326582 317384
rect 326526 315696 326582 315752
rect 326434 314200 326490 314256
rect 326526 312976 326582 313032
rect 325790 311208 325846 311264
rect 325698 246336 325754 246392
rect 325514 244976 325570 245032
rect 326434 310392 326490 310448
rect 326802 317464 326858 317520
rect 327814 357992 327870 358048
rect 327906 351056 327962 351112
rect 327630 320728 327686 320784
rect 327538 319912 327594 319968
rect 327722 320592 327778 320648
rect 327722 320456 327778 320512
rect 327722 319912 327778 319968
rect 326986 319504 327042 319560
rect 326986 316648 327042 316704
rect 326894 312976 326950 313032
rect 326618 312840 326674 312896
rect 326986 311480 327042 311536
rect 326986 311208 327042 311264
rect 326710 264152 326766 264208
rect 327262 318552 327318 318608
rect 327446 319504 327502 319560
rect 327354 317872 327410 317928
rect 327722 319368 327778 319424
rect 327446 317736 327502 317792
rect 327446 317620 327502 317656
rect 327446 317600 327448 317620
rect 327448 317600 327500 317620
rect 327500 317600 327502 317620
rect 327262 316240 327318 316296
rect 327078 257216 327134 257272
rect 326526 250552 326582 250608
rect 326434 247696 326490 247752
rect 326342 244840 326398 244896
rect 327906 317328 327962 317384
rect 327446 308488 327502 308544
rect 327262 303456 327318 303512
rect 327170 229880 327226 229936
rect 328366 365608 328422 365664
rect 328182 323584 328238 323640
rect 328090 318280 328146 318336
rect 328366 321408 328422 321464
rect 328366 320456 328422 320512
rect 328366 318960 328422 319016
rect 328274 318008 328330 318064
rect 328458 315696 328514 315752
rect 328458 311072 328514 311128
rect 327814 225800 327870 225856
rect 328918 315696 328974 315752
rect 328918 315152 328974 315208
rect 328734 237904 328790 237960
rect 329562 317872 329618 317928
rect 330390 321816 330446 321872
rect 330114 318688 330170 318744
rect 329930 318144 329986 318200
rect 329838 318008 329894 318064
rect 330114 316648 330170 316704
rect 330022 314200 330078 314256
rect 330206 314472 330262 314528
rect 330206 314200 330262 314256
rect 330114 307128 330170 307184
rect 330942 398384 330998 398440
rect 330850 314608 330906 314664
rect 330850 313792 330906 313848
rect 331218 322904 331274 322960
rect 331310 322088 331366 322144
rect 330758 310936 330814 310992
rect 328826 230424 328882 230480
rect 331402 318552 331458 318608
rect 331402 235864 331458 235920
rect 331954 395936 332010 395992
rect 333242 397160 333298 397216
rect 332690 321952 332746 322008
rect 331770 300056 331826 300112
rect 331310 235184 331366 235240
rect 332782 238720 332838 238776
rect 331218 229744 331274 229800
rect 333886 450200 333942 450256
rect 334162 398520 334218 398576
rect 334162 398248 334218 398304
rect 334806 452648 334862 452704
rect 333886 368736 333942 368792
rect 333978 319912 334034 319968
rect 333150 237224 333206 237280
rect 334070 233008 334126 233064
rect 333978 227568 334034 227624
rect 328458 223216 328514 223272
rect 322938 68176 322994 68232
rect 332690 102720 332746 102776
rect 334806 395800 334862 395856
rect 335818 452104 335874 452160
rect 335818 451696 335874 451752
rect 336002 449248 336058 449304
rect 336002 448840 336058 448896
rect 336094 402192 336150 402248
rect 335266 329160 335322 329216
rect 335174 318416 335230 318472
rect 335818 321272 335874 321328
rect 335450 320184 335506 320240
rect 335818 320184 335874 320240
rect 335358 316512 335414 316568
rect 335910 316512 335966 316568
rect 336278 397568 336334 397624
rect 336462 326440 336518 326496
rect 337474 397296 337530 397352
rect 337382 368464 337438 368520
rect 336830 320456 336886 320512
rect 337198 320456 337254 320512
rect 336738 317056 336794 317112
rect 335542 304272 335598 304328
rect 336462 304272 336518 304328
rect 336922 315288 336978 315344
rect 337934 327664 337990 327720
rect 338118 325216 338174 325272
rect 337934 317056 337990 317112
rect 338210 321680 338266 321736
rect 338118 316784 338174 316840
rect 338854 394712 338910 394768
rect 338762 368600 338818 368656
rect 339866 396208 339922 396264
rect 340234 451424 340290 451480
rect 340234 398248 340290 398304
rect 340050 365608 340106 365664
rect 340050 364928 340106 364984
rect 339498 317056 339554 317112
rect 339498 223488 339554 223544
rect 340326 396480 340382 396536
rect 350722 454008 350778 454064
rect 340878 451288 340934 451344
rect 340970 438232 341026 438288
rect 341706 438232 341762 438288
rect 341338 401784 341394 401840
rect 341430 400696 341486 400752
rect 340970 391448 341026 391504
rect 341154 390496 341210 390552
rect 341614 400288 341670 400344
rect 341890 400152 341946 400208
rect 341890 399744 341946 399800
rect 341430 398928 341486 398984
rect 341890 398792 341946 398848
rect 341338 395664 341394 395720
rect 340786 364928 340842 364984
rect 340694 337320 340750 337376
rect 340970 323720 341026 323776
rect 340694 317056 340750 317112
rect 339590 222128 339646 222184
rect 341798 391992 341854 392048
rect 344466 452104 344522 452160
rect 344098 451696 344154 451752
rect 345202 451968 345258 452024
rect 345064 450200 345120 450256
rect 347778 451832 347834 451888
rect 345938 451424 345994 451480
rect 347042 451288 347098 451344
rect 352194 451560 352250 451616
rect 352930 450200 352986 450256
rect 352930 449928 352986 449984
rect 356702 451288 356758 451344
rect 356978 451288 357034 451344
rect 346536 449520 346592 449576
rect 343822 449384 343878 449440
rect 345800 449384 345856 449440
rect 349986 449384 350042 449440
rect 359784 449384 359840 449440
rect 360934 451424 360990 451480
rect 360750 451288 360806 451344
rect 360382 449928 360438 449984
rect 361118 451424 361174 451480
rect 361486 451288 361542 451344
rect 360658 449792 360714 449848
rect 363510 451288 363566 451344
rect 363602 449928 363658 449984
rect 364154 451288 364210 451344
rect 365718 450472 365774 450528
rect 365074 449928 365130 449984
rect 368018 454144 368074 454200
rect 369122 452648 369178 452704
rect 368570 451288 368626 451344
rect 368984 450200 369040 450256
rect 369490 451288 369546 451344
rect 370456 450064 370512 450120
rect 370594 449420 370596 449440
rect 370596 449420 370648 449440
rect 370648 449420 370650 449440
rect 370594 449384 370650 449420
rect 373170 449384 373226 449440
rect 374458 452512 374514 452568
rect 377586 451288 377642 451344
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580354 511264 580410 511320
rect 580170 484608 580226 484664
rect 580078 471416 580134 471472
rect 580170 458088 580226 458144
rect 375010 449520 375066 449576
rect 374274 449384 374330 449440
rect 385314 449384 385370 449440
rect 346904 449248 346960 449304
rect 347640 449248 347696 449304
rect 359784 449248 359840 449304
rect 371192 449248 371248 449304
rect 371928 449248 371984 449304
rect 382232 449248 382288 449304
rect 383704 449248 383760 449304
rect 342442 439456 342498 439512
rect 580170 431568 580226 431624
rect 580262 418240 580318 418296
rect 580170 404912 580226 404968
rect 342258 401920 342314 401976
rect 342258 400560 342314 400616
rect 343040 399880 343096 399936
rect 342948 399744 343004 399800
rect 343224 399744 343280 399800
rect 341982 329296 342038 329352
rect 342258 320320 342314 320376
rect 342534 319232 342590 319288
rect 343178 398656 343234 398712
rect 340878 220768 340934 220824
rect 343776 399880 343832 399936
rect 344098 399744 344154 399800
rect 344328 399880 344384 399936
rect 344696 399880 344752 399936
rect 343546 393488 343602 393544
rect 343454 321000 343510 321056
rect 343822 381656 343878 381712
rect 344098 393352 344154 393408
rect 344006 319640 344062 319696
rect 344190 387232 344246 387288
rect 343546 312432 343602 312488
rect 345064 399880 345120 399936
rect 344742 398656 344798 398712
rect 344650 398520 344706 398576
rect 344650 398112 344706 398168
rect 344742 391312 344798 391368
rect 344558 389816 344614 389872
rect 344374 381928 344430 381984
rect 343638 301688 343694 301744
rect 345616 399880 345672 399936
rect 345386 397976 345442 398032
rect 345018 389000 345074 389056
rect 344926 378528 344982 378584
rect 346076 399880 346132 399936
rect 345892 399744 345948 399800
rect 346444 399880 346500 399936
rect 345662 398792 345718 398848
rect 345570 388320 345626 388376
rect 345018 325760 345074 325816
rect 344926 325352 344982 325408
rect 344926 301688 344982 301744
rect 343638 232600 343694 232656
rect 345846 389952 345902 390008
rect 345938 389816 345994 389872
rect 346306 391176 346362 391232
rect 346214 388184 346270 388240
rect 346398 387504 346454 387560
rect 347272 399880 347328 399936
rect 347456 399880 347512 399936
rect 347732 399846 347788 399902
rect 346766 399064 346822 399120
rect 346122 321136 346178 321192
rect 346306 326576 346362 326632
rect 346306 325760 346362 325816
rect 347410 399744 347466 399800
rect 348008 399880 348064 399936
rect 348376 399880 348432 399936
rect 346766 319776 346822 319832
rect 346950 319096 347006 319152
rect 347318 399200 347374 399256
rect 347962 399744 348018 399800
rect 347502 388456 347558 388512
rect 347778 399200 347834 399256
rect 347778 398792 347834 398848
rect 347870 388864 347926 388920
rect 347226 381656 347282 381712
rect 349204 399880 349260 399936
rect 349112 399744 349168 399800
rect 348422 399064 348478 399120
rect 347962 374720 348018 374776
rect 348698 399064 348754 399120
rect 348698 398248 348754 398304
rect 348514 393352 348570 393408
rect 348882 377848 348938 377904
rect 350032 399744 350088 399800
rect 349342 393352 349398 393408
rect 349526 379208 349582 379264
rect 349434 378664 349490 378720
rect 349342 357992 349398 358048
rect 350400 399880 350456 399936
rect 350768 399880 350824 399936
rect 351044 399880 351100 399936
rect 350538 397432 350594 397488
rect 350170 390088 350226 390144
rect 349986 382064 350042 382120
rect 350078 377984 350134 378040
rect 351596 399880 351652 399936
rect 351780 399880 351836 399936
rect 351826 399744 351882 399800
rect 350906 395936 350962 395992
rect 351550 398556 351552 398576
rect 351552 398556 351604 398576
rect 351604 398556 351606 398576
rect 351550 398520 351606 398556
rect 351090 390224 351146 390280
rect 350906 379344 350962 379400
rect 350998 379072 351054 379128
rect 350814 378800 350870 378856
rect 350722 359352 350778 359408
rect 352470 399744 352526 399800
rect 352378 396752 352434 396808
rect 352378 396344 352434 396400
rect 352286 395392 352342 395448
rect 351550 381792 351606 381848
rect 352286 378936 352342 378992
rect 352884 399744 352940 399800
rect 353436 399880 353492 399936
rect 352930 397432 352986 397488
rect 353298 399336 353354 399392
rect 353988 399880 354044 399936
rect 354172 399880 354228 399936
rect 353482 399336 353538 399392
rect 353482 397160 353538 397216
rect 353482 396752 353538 396808
rect 353022 391040 353078 391096
rect 353574 381520 353630 381576
rect 352746 317192 352802 317248
rect 354034 399064 354090 399120
rect 354402 399200 354458 399256
rect 354586 399200 354642 399256
rect 355368 399880 355424 399936
rect 354678 395936 354734 395992
rect 355414 399608 355470 399664
rect 355782 398656 355838 398712
rect 355598 394304 355654 394360
rect 355598 393760 355654 393816
rect 356150 399336 356206 399392
rect 356334 398792 356390 398848
rect 356518 397432 356574 397488
rect 356426 394576 356482 394632
rect 356886 399608 356942 399664
rect 356334 375944 356390 376000
rect 356242 374584 356298 374640
rect 357162 398792 357218 398848
rect 356978 396888 357034 396944
rect 357346 399336 357402 399392
rect 357622 399608 357678 399664
rect 357530 397976 357586 398032
rect 357438 397432 357494 397488
rect 357898 399608 357954 399664
rect 357622 387368 357678 387424
rect 357898 399200 357954 399256
rect 357530 384376 357586 384432
rect 358082 399336 358138 399392
rect 358082 397296 358138 397352
rect 358266 399200 358322 399256
rect 358450 398112 358506 398168
rect 358358 397840 358414 397896
rect 357898 393216 357954 393272
rect 358082 392536 358138 392592
rect 359462 399608 359518 399664
rect 358910 396888 358966 396944
rect 359922 396344 359978 396400
rect 359922 394032 359978 394088
rect 360290 396480 360346 396536
rect 360750 399744 360806 399800
rect 361716 399744 361772 399800
rect 360474 393216 360530 393272
rect 360566 392808 360622 392864
rect 360474 385872 360530 385928
rect 361394 397704 361450 397760
rect 361302 392944 361358 393000
rect 361762 396344 361818 396400
rect 362544 399744 362600 399800
rect 362038 396616 362094 396672
rect 361946 396072 362002 396128
rect 363050 396888 363106 396944
rect 362866 392672 362922 392728
rect 362774 392400 362830 392456
rect 363924 399744 363980 399800
rect 364062 399336 364118 399392
rect 364062 398928 364118 398984
rect 363694 312568 363750 312624
rect 364614 399336 364670 399392
rect 364890 399200 364946 399256
rect 365258 397296 365314 397352
rect 365856 399880 365912 399936
rect 366316 399880 366372 399936
rect 365810 399608 365866 399664
rect 365626 397568 365682 397624
rect 366408 399744 366464 399800
rect 366776 399880 366832 399936
rect 365902 393080 365958 393136
rect 366822 399608 366878 399664
rect 366638 393896 366694 393952
rect 367236 399744 367292 399800
rect 367696 399880 367752 399936
rect 367282 393216 367338 393272
rect 367282 392808 367338 392864
rect 367650 399744 367706 399800
rect 367558 399236 367560 399256
rect 367560 399236 367612 399256
rect 367612 399236 367614 399256
rect 367558 399200 367614 399236
rect 368064 399880 368120 399936
rect 367650 395800 367706 395856
rect 367650 392944 367706 393000
rect 367282 377440 367338 377496
rect 367098 315560 367154 315616
rect 336738 66816 336794 66872
rect 340970 65456 341026 65512
rect 343638 115232 343694 115288
rect 350538 64096 350594 64152
rect 354678 62736 354734 62792
rect 357530 40568 357586 40624
rect 367926 397296 367982 397352
rect 368018 393216 368074 393272
rect 368386 395120 368442 395176
rect 369444 399880 369500 399936
rect 369720 399880 369776 399936
rect 369030 397160 369086 397216
rect 368846 395528 368902 395584
rect 368938 394576 368994 394632
rect 369490 398248 369546 398304
rect 369582 393488 369638 393544
rect 371008 399880 371064 399936
rect 370824 399744 370880 399800
rect 371100 399744 371156 399800
rect 371376 399846 371432 399902
rect 370134 393080 370190 393136
rect 370502 399064 370558 399120
rect 371744 399880 371800 399936
rect 371928 399880 371984 399936
rect 372204 399880 372260 399936
rect 372572 399880 372628 399936
rect 371238 398384 371294 398440
rect 371054 396480 371110 396536
rect 365810 6432 365866 6488
rect 372158 399744 372214 399800
rect 372388 399744 372444 399800
rect 372940 399880 372996 399936
rect 372250 397568 372306 397624
rect 372342 397160 372398 397216
rect 373952 399846 374008 399902
rect 372434 389680 372490 389736
rect 372986 399608 373042 399664
rect 372986 399472 373042 399528
rect 373078 397296 373134 397352
rect 373400 399744 373456 399800
rect 374136 399846 374192 399902
rect 373354 399608 373410 399664
rect 373446 395392 373502 395448
rect 373538 393896 373594 393952
rect 373906 390904 373962 390960
rect 374090 399608 374146 399664
rect 374872 399744 374928 399800
rect 374458 399200 374514 399256
rect 374090 393760 374146 393816
rect 373906 389136 373962 389192
rect 373906 383696 373962 383752
rect 373906 383560 373962 383616
rect 373906 374040 373962 374096
rect 373906 373904 373962 373960
rect 373906 364384 373962 364440
rect 373906 364248 373962 364304
rect 373906 354728 373962 354784
rect 373906 354592 373962 354648
rect 374182 351056 374238 351112
rect 373906 345072 373962 345128
rect 373906 344936 373962 344992
rect 373906 340720 373962 340776
rect 373906 331200 373962 331256
rect 373906 325760 373962 325816
rect 375332 399880 375388 399936
rect 374826 399472 374882 399528
rect 374918 397296 374974 397352
rect 375194 395392 375250 395448
rect 376252 399880 376308 399936
rect 375470 398928 375526 398984
rect 375378 396888 375434 396944
rect 374734 377304 374790 377360
rect 376022 370504 376078 370560
rect 375930 369008 375986 369064
rect 375562 311344 375618 311400
rect 376298 397976 376354 398032
rect 376988 399880 377044 399936
rect 377264 399880 377320 399936
rect 377632 399880 377688 399936
rect 377908 399880 377964 399936
rect 376666 399472 376722 399528
rect 376942 399064 376998 399120
rect 376942 395256 376998 395312
rect 377310 399064 377366 399120
rect 377034 315968 377090 316024
rect 377586 390360 377642 390416
rect 377310 304680 377366 304736
rect 377862 399608 377918 399664
rect 378368 399880 378424 399936
rect 377770 323584 377826 323640
rect 378046 396752 378102 396808
rect 378230 399472 378286 399528
rect 378322 395120 378378 395176
rect 378138 393488 378194 393544
rect 378138 389272 378194 389328
rect 378046 321680 378102 321736
rect 376022 151136 376078 151192
rect 376482 6296 376538 6352
rect 378828 399880 378884 399936
rect 378598 399508 378600 399528
rect 378600 399508 378652 399528
rect 378652 399508 378654 399528
rect 378598 399472 378654 399508
rect 378966 399608 379022 399664
rect 379288 399880 379344 399936
rect 379472 399880 379528 399936
rect 379656 399846 379712 399902
rect 379242 399200 379298 399256
rect 379334 396616 379390 396672
rect 379932 399880 379988 399936
rect 380208 399880 380264 399936
rect 380116 399744 380172 399800
rect 379978 399608 380034 399664
rect 380162 399472 380218 399528
rect 379702 396616 379758 396672
rect 379794 314064 379850 314120
rect 380254 395664 380310 395720
rect 381036 399880 381092 399936
rect 380806 399200 380862 399256
rect 380714 397840 380770 397896
rect 380530 395256 380586 395312
rect 381680 399880 381736 399936
rect 381174 399608 381230 399664
rect 381174 396480 381230 396536
rect 381542 394168 381598 394224
rect 381818 397704 381874 397760
rect 382094 397568 382150 397624
rect 382692 399880 382748 399936
rect 382968 399744 383024 399800
rect 382278 397432 382334 397488
rect 382462 397296 382518 397352
rect 381910 315696 381966 315752
rect 383152 399744 383208 399800
rect 382830 399472 382886 399528
rect 383106 399472 383162 399528
rect 382554 312704 382610 312760
rect 382462 311072 382518 311128
rect 380898 310256 380954 310312
rect 383474 397568 383530 397624
rect 383980 399744 384036 399800
rect 383842 399608 383898 399664
rect 384348 399880 384404 399936
rect 384624 399778 384680 399834
rect 384670 399608 384726 399664
rect 384900 399880 384956 399936
rect 385176 399880 385232 399936
rect 384762 398112 384818 398168
rect 383934 320864 383990 320920
rect 383842 310120 383898 310176
rect 385360 399880 385416 399936
rect 385728 399778 385784 399834
rect 385222 399608 385278 399664
rect 385406 397296 385462 397352
rect 385314 325080 385370 325136
rect 386372 399880 386428 399936
rect 386832 399744 386888 399800
rect 387154 399608 387210 399664
rect 386970 355272 387026 355328
rect 386786 330384 386842 330440
rect 386970 329024 387026 329080
rect 386694 326304 386750 326360
rect 386602 321544 386658 321600
rect 387062 321544 387118 321600
rect 385498 317328 385554 317384
rect 385130 315832 385186 315888
rect 384854 308896 384910 308952
rect 383198 308624 383254 308680
rect 383014 303184 383070 303240
rect 379978 9424 380034 9480
rect 387798 400288 387854 400344
rect 387338 312840 387394 312896
rect 387154 310392 387210 310448
rect 390006 400016 390062 400072
rect 388166 399472 388222 399528
rect 388166 320728 388222 320784
rect 388074 314472 388130 314528
rect 387982 314200 388038 314256
rect 389362 314608 389418 314664
rect 390834 399880 390890 399936
rect 389454 314336 389510 314392
rect 391938 398112 391994 398168
rect 392214 399336 392270 399392
rect 392214 313112 392270 313168
rect 392122 311752 392178 311808
rect 392030 311480 392086 311536
rect 580262 378392 580318 378448
rect 416778 328480 416834 328536
rect 394790 312432 394846 312488
rect 394698 311072 394754 311128
rect 391938 303456 391994 303512
rect 387154 9288 387210 9344
rect 390650 6160 390706 6216
rect 394238 9152 394294 9208
rect 398930 324400 398986 324456
rect 407210 54440 407266 54496
rect 412638 122032 412694 122088
rect 411258 51720 411314 51776
rect 477498 313928 477554 313984
rect 415490 9016 415546 9072
rect 422574 8880 422630 8936
rect 426438 120672 426494 120728
rect 431222 156576 431278 156632
rect 430578 30912 430634 30968
rect 440330 11600 440386 11656
rect 447782 117952 447838 118008
rect 454038 98640 454094 98696
rect 456890 46144 456946 46200
rect 460938 44784 460994 44840
rect 465078 115096 465134 115152
rect 468482 131688 468538 131744
rect 472622 124752 472678 124808
rect 476118 113736 476174 113792
rect 474738 42064 474794 42120
rect 485778 109656 485834 109712
rect 487158 37848 487214 37904
rect 490010 18536 490066 18592
rect 496818 106800 496874 106856
rect 513378 329840 513434 329896
rect 498290 151000 498346 151056
rect 500958 148416 501014 148472
rect 506570 104080 506626 104136
rect 580170 365064 580226 365120
rect 580262 364928 580318 364984
rect 514850 101360 514906 101416
rect 517518 71032 517574 71088
rect 529938 149640 529994 149696
rect 528558 69536 528614 69592
rect 531410 95784 531466 95840
rect 536838 119312 536894 119368
rect 543738 148280 543794 148336
rect 556250 311072 556306 311128
rect 548522 90344 548578 90400
rect 547970 35128 548026 35184
rect 557538 153720 557594 153776
rect 561678 146920 561734 146976
rect 564438 84768 564494 84824
rect 579986 325216 580042 325272
rect 572810 312432 572866 312488
rect 571982 306448 572038 306504
rect 571522 7520 571578 7576
rect 579618 312024 579674 312080
rect 580170 298732 580172 298752
rect 580172 298732 580224 298752
rect 580224 298732 580226 298752
rect 580170 298696 580226 298732
rect 579618 245556 579620 245576
rect 579620 245556 579672 245576
rect 579672 245556 579674 245576
rect 579618 245520 579674 245556
rect 579618 232328 579674 232384
rect 579986 205672 580042 205728
rect 580170 192480 580226 192536
rect 579894 152632 579950 152688
rect 580446 366288 580502 366344
rect 580354 219000 580410 219056
rect 580354 206216 580410 206272
rect 580262 139304 580318 139360
rect 580170 99456 580226 99512
rect 580262 86128 580318 86184
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580078 19760 580134 19816
rect 580538 360848 580594 360904
rect 580722 351872 580778 351928
rect 580630 272176 580686 272232
rect 580538 258848 580594 258904
rect 580722 209072 580778 209128
rect 580538 208936 580594 208992
rect 580446 179152 580502 179208
rect 580722 165824 580778 165880
rect 580538 125976 580594 126032
rect 580354 6568 580410 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580349 511322 580415 511325
rect 583520 511322 584960 511412
rect 580349 511320 584960 511322
rect 580349 511264 580354 511320
rect 580410 511264 584960 511320
rect 580349 511262 584960 511264
rect 580349 511259 580415 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580073 471474 580139 471477
rect 583520 471474 584960 471564
rect 580073 471472 584960 471474
rect 580073 471416 580078 471472
rect 580134 471416 584960 471472
rect 580073 471414 584960 471416
rect 580073 471411 580139 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 308397 454202 308463 454205
rect 368013 454202 368079 454205
rect 308397 454200 368079 454202
rect 308397 454144 308402 454200
rect 308458 454144 368018 454200
rect 368074 454144 368079 454200
rect 308397 454142 368079 454144
rect 308397 454139 308463 454142
rect 368013 454139 368079 454142
rect 280061 454066 280127 454069
rect 350717 454066 350783 454069
rect 280061 454064 350783 454066
rect 280061 454008 280066 454064
rect 280122 454008 350722 454064
rect 350778 454008 350783 454064
rect 280061 454006 350783 454008
rect 280061 454003 280127 454006
rect 350717 454003 350783 454006
rect 334801 452706 334867 452709
rect 369117 452706 369183 452709
rect 334801 452704 369183 452706
rect 334801 452648 334806 452704
rect 334862 452648 369122 452704
rect 369178 452648 369183 452704
rect 334801 452646 369183 452648
rect 334801 452643 334867 452646
rect 369117 452643 369183 452646
rect 374126 452508 374132 452572
rect 374196 452570 374202 452572
rect 374453 452570 374519 452573
rect 374196 452568 374519 452570
rect 374196 452512 374458 452568
rect 374514 452512 374519 452568
rect 374196 452510 374519 452512
rect 374196 452508 374202 452510
rect 374453 452507 374519 452510
rect 335813 452162 335879 452165
rect 344461 452162 344527 452165
rect 335813 452160 344527 452162
rect 335813 452104 335818 452160
rect 335874 452104 344466 452160
rect 344522 452104 344527 452160
rect 335813 452102 344527 452104
rect 335813 452099 335879 452102
rect 344461 452099 344527 452102
rect 280613 452026 280679 452029
rect 345197 452026 345263 452029
rect 280613 452024 345263 452026
rect 280613 451968 280618 452024
rect 280674 451968 345202 452024
rect 345258 451968 345263 452024
rect 280613 451966 345263 451968
rect 280613 451963 280679 451966
rect 345197 451963 345263 451966
rect 278630 451828 278636 451892
rect 278700 451890 278706 451892
rect 347773 451890 347839 451893
rect 278700 451888 347839 451890
rect 278700 451832 347778 451888
rect 347834 451832 347839 451888
rect 278700 451830 347839 451832
rect 278700 451828 278706 451830
rect 347773 451827 347839 451830
rect 282821 451754 282887 451757
rect 335813 451754 335879 451757
rect 344093 451754 344159 451757
rect 282821 451752 335879 451754
rect 282821 451696 282826 451752
rect 282882 451696 335818 451752
rect 335874 451696 335879 451752
rect 282821 451694 335879 451696
rect 282821 451691 282887 451694
rect 335813 451691 335879 451694
rect 340830 451752 344159 451754
rect 340830 451696 344098 451752
rect 344154 451696 344159 451752
rect 340830 451694 344159 451696
rect 280889 451618 280955 451621
rect 340830 451618 340890 451694
rect 344093 451691 344159 451694
rect 280889 451616 340890 451618
rect 280889 451560 280894 451616
rect 280950 451560 340890 451616
rect 280889 451558 340890 451560
rect 280889 451555 280955 451558
rect 343950 451556 343956 451620
rect 344020 451618 344026 451620
rect 352189 451618 352255 451621
rect 344020 451616 352255 451618
rect 344020 451560 352194 451616
rect 352250 451560 352255 451616
rect 344020 451558 352255 451560
rect 344020 451556 344026 451558
rect 352189 451555 352255 451558
rect 340229 451482 340295 451485
rect 345933 451482 345999 451485
rect 340229 451480 345999 451482
rect 340229 451424 340234 451480
rect 340290 451424 345938 451480
rect 345994 451424 345999 451480
rect 340229 451422 345999 451424
rect 340229 451419 340295 451422
rect 345933 451419 345999 451422
rect 360929 451482 360995 451485
rect 361113 451482 361179 451485
rect 360929 451480 361179 451482
rect 360929 451424 360934 451480
rect 360990 451424 361118 451480
rect 361174 451424 361179 451480
rect 360929 451422 361179 451424
rect 360929 451419 360995 451422
rect 361113 451419 361179 451422
rect 340873 451346 340939 451349
rect 347037 451346 347103 451349
rect 340873 451344 347103 451346
rect 340873 451288 340878 451344
rect 340934 451288 347042 451344
rect 347098 451288 347103 451344
rect 340873 451286 347103 451288
rect 340873 451283 340939 451286
rect 347037 451283 347103 451286
rect 355174 451284 355180 451348
rect 355244 451346 355250 451348
rect 356697 451346 356763 451349
rect 356973 451346 357039 451349
rect 355244 451344 357039 451346
rect 355244 451288 356702 451344
rect 356758 451288 356978 451344
rect 357034 451288 357039 451344
rect 355244 451286 357039 451288
rect 355244 451284 355250 451286
rect 356697 451283 356763 451286
rect 356973 451283 357039 451286
rect 360745 451346 360811 451349
rect 361481 451346 361547 451349
rect 360745 451344 361547 451346
rect 360745 451288 360750 451344
rect 360806 451288 361486 451344
rect 361542 451288 361547 451344
rect 360745 451286 361547 451288
rect 360745 451283 360811 451286
rect 361481 451283 361547 451286
rect 362902 451284 362908 451348
rect 362972 451346 362978 451348
rect 363505 451346 363571 451349
rect 364149 451346 364215 451349
rect 362972 451344 364215 451346
rect 362972 451288 363510 451344
rect 363566 451288 364154 451344
rect 364210 451288 364215 451344
rect 362972 451286 364215 451288
rect 362972 451284 362978 451286
rect 363505 451283 363571 451286
rect 364149 451283 364215 451286
rect 368238 451284 368244 451348
rect 368308 451346 368314 451348
rect 368565 451346 368631 451349
rect 369485 451346 369551 451349
rect 368308 451344 369551 451346
rect 368308 451288 368570 451344
rect 368626 451288 369490 451344
rect 369546 451288 369551 451344
rect 368308 451286 369551 451288
rect 368308 451284 368314 451286
rect 368565 451283 368631 451286
rect 369485 451283 369551 451286
rect 376886 451284 376892 451348
rect 376956 451346 376962 451348
rect 377581 451346 377647 451349
rect 376956 451344 377647 451346
rect 376956 451288 377586 451344
rect 377642 451288 377647 451344
rect 376956 451286 377647 451288
rect 376956 451284 376962 451286
rect 377581 451283 377647 451286
rect 6913 450530 6979 450533
rect 309133 450530 309199 450533
rect 365713 450530 365779 450533
rect 6913 450528 365779 450530
rect 6913 450472 6918 450528
rect 6974 450472 309138 450528
rect 309194 450472 365718 450528
rect 365774 450472 365779 450528
rect 6913 450470 365779 450472
rect 6913 450467 6979 450470
rect 309133 450467 309199 450470
rect 365713 450467 365779 450470
rect 333881 450258 333947 450261
rect 345059 450258 345125 450261
rect 333881 450256 345125 450258
rect 333881 450200 333886 450256
rect 333942 450200 345064 450256
rect 345120 450200 345125 450256
rect 333881 450198 345125 450200
rect 333881 450195 333947 450198
rect 345059 450195 345125 450198
rect 352925 450258 352991 450261
rect 368979 450258 369045 450261
rect 352925 450256 369045 450258
rect 352925 450200 352930 450256
rect 352986 450200 368984 450256
rect 369040 450200 369045 450256
rect 352925 450198 369045 450200
rect 352925 450195 352991 450198
rect 368979 450195 369045 450198
rect 309869 450122 309935 450125
rect 370451 450122 370517 450125
rect 309869 450120 370517 450122
rect 309869 450064 309874 450120
rect 309930 450064 370456 450120
rect 370512 450064 370517 450120
rect 309869 450062 370517 450064
rect 309869 450059 309935 450062
rect 370451 450059 370517 450062
rect 307661 449986 307727 449989
rect 352925 449986 352991 449989
rect 360377 449988 360443 449989
rect 307661 449984 352991 449986
rect 307661 449928 307666 449984
rect 307722 449928 352930 449984
rect 352986 449928 352991 449984
rect 307661 449926 352991 449928
rect 307661 449923 307727 449926
rect 352925 449923 352991 449926
rect 360326 449924 360332 449988
rect 360396 449986 360443 449988
rect 360396 449984 360488 449986
rect 360438 449928 360488 449984
rect 360396 449926 360488 449928
rect 360396 449924 360443 449926
rect 363270 449924 363276 449988
rect 363340 449986 363346 449988
rect 363597 449986 363663 449989
rect 363340 449984 363663 449986
rect 363340 449928 363602 449984
rect 363658 449928 363663 449984
rect 363340 449926 363663 449928
rect 363340 449924 363346 449926
rect 360377 449923 360443 449924
rect 363597 449923 363663 449926
rect 364374 449924 364380 449988
rect 364444 449986 364450 449988
rect 365069 449986 365135 449989
rect 364444 449984 365135 449986
rect 364444 449928 365074 449984
rect 365130 449928 365135 449984
rect 364444 449926 365135 449928
rect 364444 449924 364450 449926
rect 365069 449923 365135 449926
rect 360510 449788 360516 449852
rect 360580 449850 360586 449852
rect 360653 449850 360719 449853
rect 360580 449848 360719 449850
rect 360580 449792 360658 449848
rect 360714 449792 360719 449848
rect 360580 449790 360719 449792
rect 360580 449788 360586 449790
rect 360653 449787 360719 449790
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 331489 449578 331555 449581
rect 346531 449578 346597 449581
rect 331489 449576 346597 449578
rect 331489 449520 331494 449576
rect 331550 449520 346536 449576
rect 346592 449520 346597 449576
rect 331489 449518 346597 449520
rect 331489 449515 331555 449518
rect 346531 449515 346597 449518
rect 374126 449516 374132 449580
rect 374196 449578 374202 449580
rect 375005 449578 375071 449581
rect 374196 449576 375071 449578
rect 374196 449520 375010 449576
rect 375066 449520 375071 449576
rect 374196 449518 375071 449520
rect 374196 449516 374202 449518
rect 375005 449515 375071 449518
rect 343817 449444 343883 449445
rect 345795 449444 345861 449445
rect 343766 449442 343772 449444
rect 343726 449382 343772 449442
rect 343836 449440 343883 449444
rect 345790 449442 345796 449444
rect 343878 449384 343883 449440
rect 343766 449380 343772 449382
rect 343836 449380 343883 449384
rect 345704 449382 345796 449442
rect 345790 449380 345796 449382
rect 345860 449380 345866 449444
rect 347446 449380 347452 449444
rect 347516 449442 347522 449444
rect 349981 449442 350047 449445
rect 347516 449440 350047 449442
rect 347516 449384 349986 449440
rect 350042 449384 350047 449440
rect 347516 449382 350047 449384
rect 347516 449380 347522 449382
rect 343817 449379 343883 449380
rect 345795 449379 345861 449380
rect 349981 449379 350047 449382
rect 359779 449440 359845 449445
rect 359779 449384 359784 449440
rect 359840 449384 359845 449440
rect 359779 449379 359845 449384
rect 370446 449380 370452 449444
rect 370516 449442 370522 449444
rect 370589 449442 370655 449445
rect 373165 449444 373231 449445
rect 374269 449444 374335 449445
rect 373165 449442 373212 449444
rect 370516 449440 370655 449442
rect 370516 449384 370594 449440
rect 370650 449384 370655 449440
rect 370516 449382 370655 449384
rect 373120 449440 373212 449442
rect 373120 449384 373170 449440
rect 373120 449382 373212 449384
rect 370516 449380 370522 449382
rect 370589 449379 370655 449382
rect 373165 449380 373212 449382
rect 373276 449380 373282 449444
rect 374269 449442 374316 449444
rect 374224 449440 374316 449442
rect 374224 449384 374274 449440
rect 374224 449382 374316 449384
rect 374269 449380 374316 449382
rect 374380 449380 374386 449444
rect 384982 449380 384988 449444
rect 385052 449442 385058 449444
rect 385309 449442 385375 449445
rect 385052 449440 385375 449442
rect 385052 449384 385314 449440
rect 385370 449384 385375 449440
rect 385052 449382 385375 449384
rect 385052 449380 385058 449382
rect 373165 449379 373231 449380
rect 374269 449379 374335 449380
rect 385309 449379 385375 449382
rect 359782 449309 359842 449379
rect 335997 449306 336063 449309
rect 346899 449306 346965 449309
rect 347635 449308 347701 449309
rect 347630 449306 347636 449308
rect 335997 449304 346965 449306
rect 335997 449248 336002 449304
rect 336058 449248 346904 449304
rect 346960 449248 346965 449304
rect 335997 449246 346965 449248
rect 347544 449246 347636 449306
rect 335997 449243 336063 449246
rect 346899 449243 346965 449246
rect 347630 449244 347636 449246
rect 347700 449244 347706 449308
rect 359779 449304 359845 449309
rect 371187 449308 371253 449309
rect 371182 449306 371188 449308
rect 359779 449248 359784 449304
rect 359840 449248 359845 449304
rect 347635 449243 347701 449244
rect 359779 449243 359845 449248
rect 371096 449246 371188 449306
rect 371182 449244 371188 449246
rect 371252 449244 371258 449308
rect 371923 449304 371989 449309
rect 382227 449308 382293 449309
rect 383699 449308 383765 449309
rect 382222 449306 382228 449308
rect 371923 449248 371928 449304
rect 371984 449248 371989 449304
rect 371187 449243 371253 449244
rect 371923 449243 371989 449248
rect 382136 449246 382228 449306
rect 382222 449244 382228 449246
rect 382292 449244 382298 449308
rect 383694 449244 383700 449308
rect 383764 449306 383770 449308
rect 383764 449246 383856 449306
rect 383764 449244 383770 449246
rect 382227 449243 382293 449244
rect 383699 449243 383765 449244
rect 300209 449170 300275 449173
rect 359782 449170 359842 449243
rect 300209 449168 359842 449170
rect 300209 449112 300214 449168
rect 300270 449112 359842 449168
rect 300209 449110 359842 449112
rect 300209 449107 300275 449110
rect 312537 449034 312603 449037
rect 371926 449034 371986 449243
rect 312537 449032 371986 449034
rect 312537 448976 312542 449032
rect 312598 448976 371986 449032
rect 312537 448974 371986 448976
rect 312537 448971 312603 448974
rect 285949 448898 286015 448901
rect 335997 448898 336063 448901
rect 285949 448896 336063 448898
rect 285949 448840 285954 448896
rect 286010 448840 336002 448896
rect 336058 448840 336063 448896
rect 285949 448838 336063 448840
rect 285949 448835 286015 448838
rect 335997 448835 336063 448838
rect 282177 448762 282243 448765
rect 331489 448762 331555 448765
rect 282177 448760 331555 448762
rect 282177 448704 282182 448760
rect 282238 448704 331494 448760
rect 331550 448704 331555 448760
rect 282177 448702 331555 448704
rect 282177 448699 282243 448702
rect 331489 448699 331555 448702
rect 278313 448626 278379 448629
rect 347630 448626 347636 448628
rect 278313 448624 347636 448626
rect 278313 448568 278318 448624
rect 278374 448568 347636 448624
rect 278313 448566 347636 448568
rect 278313 448563 278379 448566
rect 347630 448564 347636 448566
rect 347700 448564 347706 448628
rect 290457 447946 290523 447949
rect 347446 447946 347452 447948
rect 290457 447944 347452 447946
rect 290457 447888 290462 447944
rect 290518 447888 347452 447944
rect 290457 447886 347452 447888
rect 290457 447883 290523 447886
rect 347446 447884 347452 447886
rect 347516 447884 347522 447948
rect 286317 447810 286383 447813
rect 345790 447810 345796 447812
rect 286317 447808 345796 447810
rect 286317 447752 286322 447808
rect 286378 447752 345796 447808
rect 286317 447750 345796 447752
rect 286317 447747 286383 447750
rect 345790 447748 345796 447750
rect 345860 447748 345866 447812
rect 360142 447476 360148 447540
rect 360212 447538 360218 447540
rect 360510 447538 360516 447540
rect 360212 447478 360516 447538
rect 360212 447476 360218 447478
rect 360510 447476 360516 447478
rect 360580 447476 360586 447540
rect 583520 444668 584960 444908
rect 291837 443594 291903 443597
rect 343950 443594 343956 443596
rect 291837 443592 343956 443594
rect 291837 443536 291842 443592
rect 291898 443536 343956 443592
rect 291837 443534 343956 443536
rect 291837 443531 291903 443534
rect 343950 443532 343956 443534
rect 344020 443532 344026 443596
rect 304257 439514 304323 439517
rect 342437 439514 342503 439517
rect 304257 439512 342503 439514
rect 304257 439456 304262 439512
rect 304318 439456 342442 439512
rect 342498 439456 342503 439512
rect 304257 439454 342503 439456
rect 304257 439451 304323 439454
rect 342437 439451 342503 439454
rect 340965 438290 341031 438293
rect 341701 438290 341767 438293
rect 340965 438288 341767 438290
rect 340965 438232 340970 438288
rect 341026 438232 341706 438288
rect 341762 438232 341767 438288
rect 340965 438230 341767 438232
rect 340965 438227 341031 438230
rect 341701 438227 341767 438230
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 4061 410546 4127 410549
rect -960 410544 4127 410546
rect -960 410488 4066 410544
rect 4122 410488 4127 410544
rect -960 410486 4127 410488
rect -960 410396 480 410486
rect 4061 410483 4127 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 71773 404290 71839 404293
rect 307661 404292 307727 404293
rect 307661 404290 307708 404292
rect 71773 404288 307708 404290
rect 307772 404290 307778 404292
rect 71773 404232 71778 404288
rect 71834 404232 307666 404288
rect 71773 404230 307708 404232
rect 71773 404227 71839 404230
rect 307661 404228 307708 404230
rect 307772 404230 307854 404290
rect 307772 404228 307778 404230
rect 307661 404227 307727 404228
rect 336089 402250 336155 402253
rect 343950 402250 343956 402252
rect 336089 402248 343956 402250
rect 336089 402192 336094 402248
rect 336150 402192 343956 402248
rect 336089 402190 343956 402192
rect 336089 402187 336155 402190
rect 343950 402188 343956 402190
rect 344020 402188 344026 402252
rect 265801 402114 265867 402117
rect 343030 402114 343036 402116
rect 265801 402112 343036 402114
rect 265801 402056 265806 402112
rect 265862 402056 343036 402112
rect 265801 402054 343036 402056
rect 265801 402051 265867 402054
rect 343030 402052 343036 402054
rect 343100 402052 343106 402116
rect 266261 401978 266327 401981
rect 342253 401978 342319 401981
rect 266261 401976 342319 401978
rect 266261 401920 266266 401976
rect 266322 401920 342258 401976
rect 342314 401920 342319 401976
rect 266261 401918 342319 401920
rect 266261 401915 266327 401918
rect 342253 401915 342319 401918
rect 360142 401916 360148 401980
rect 360212 401978 360218 401980
rect 360510 401978 360516 401980
rect 360212 401918 360516 401978
rect 360212 401916 360218 401918
rect 360510 401916 360516 401918
rect 360580 401916 360586 401980
rect 263317 401842 263383 401845
rect 341333 401842 341399 401845
rect 263317 401840 341399 401842
rect 263317 401784 263322 401840
rect 263378 401784 341338 401840
rect 341394 401784 341399 401840
rect 263317 401782 341399 401784
rect 263317 401779 263383 401782
rect 341333 401779 341399 401782
rect 265617 401706 265683 401709
rect 347630 401706 347636 401708
rect 265617 401704 347636 401706
rect 265617 401648 265622 401704
rect 265678 401648 347636 401704
rect 265617 401646 347636 401648
rect 265617 401643 265683 401646
rect 347630 401644 347636 401646
rect 347700 401644 347706 401708
rect 311249 401570 311315 401573
rect 371182 401570 371188 401572
rect 311249 401568 371188 401570
rect 311249 401512 311254 401568
rect 311310 401512 371188 401568
rect 311249 401510 371188 401512
rect 311249 401507 311315 401510
rect 371182 401508 371188 401510
rect 371252 401508 371258 401572
rect 297541 401298 297607 401301
rect 355174 401298 355180 401300
rect 297541 401296 355180 401298
rect 297541 401240 297546 401296
rect 297602 401240 355180 401296
rect 297541 401238 355180 401240
rect 297541 401235 297607 401238
rect 355174 401236 355180 401238
rect 355244 401236 355250 401300
rect 303521 401162 303587 401165
rect 362902 401162 362908 401164
rect 303521 401160 362908 401162
rect 303521 401104 303526 401160
rect 303582 401104 362908 401160
rect 303521 401102 362908 401104
rect 303521 401099 303587 401102
rect 362902 401100 362908 401102
rect 362972 401100 362978 401164
rect 300393 401026 300459 401029
rect 360326 401026 360332 401028
rect 300393 401024 360332 401026
rect 300393 400968 300398 401024
rect 300454 400968 360332 401024
rect 300393 400966 360332 400968
rect 300393 400963 300459 400966
rect 360326 400964 360332 400966
rect 360396 400964 360402 401028
rect 314101 400890 314167 400893
rect 374310 400890 374316 400892
rect 314101 400888 374316 400890
rect 314101 400832 314106 400888
rect 314162 400832 374316 400888
rect 314101 400830 374316 400832
rect 314101 400827 314167 400830
rect 374310 400828 374316 400830
rect 374380 400828 374386 400892
rect 341425 400754 341491 400757
rect 352414 400754 352420 400756
rect 341425 400752 352420 400754
rect 341425 400696 341430 400752
rect 341486 400696 352420 400752
rect 341425 400694 352420 400696
rect 341425 400691 341491 400694
rect 352414 400692 352420 400694
rect 352484 400692 352490 400756
rect 342253 400618 342319 400621
rect 355358 400618 355364 400620
rect 342253 400616 355364 400618
rect 342253 400560 342258 400616
rect 342314 400560 355364 400616
rect 342253 400558 355364 400560
rect 342253 400555 342319 400558
rect 355358 400556 355364 400558
rect 355428 400556 355434 400620
rect 343766 400482 343772 400484
rect 340830 400422 343772 400482
rect 266997 400346 267063 400349
rect 340830 400346 340890 400422
rect 343766 400420 343772 400422
rect 343836 400420 343842 400484
rect 266997 400344 340890 400346
rect 266997 400288 267002 400344
rect 267058 400288 340890 400344
rect 266997 400286 340890 400288
rect 341609 400346 341675 400349
rect 345790 400346 345796 400348
rect 341609 400344 345796 400346
rect 341609 400288 341614 400344
rect 341670 400288 345796 400344
rect 341609 400286 345796 400288
rect 266997 400283 267063 400286
rect 341609 400283 341675 400286
rect 345790 400284 345796 400286
rect 345860 400284 345866 400348
rect 354070 400346 354076 400348
rect 346350 400286 354076 400346
rect 341885 400210 341951 400213
rect 346350 400210 346410 400286
rect 354070 400284 354076 400286
rect 354140 400284 354146 400348
rect 387793 400346 387859 400349
rect 378228 400344 387859 400346
rect 378228 400288 387798 400344
rect 387854 400288 387859 400344
rect 378228 400286 387859 400288
rect 355542 400210 355548 400212
rect 341885 400208 346410 400210
rect 341885 400152 341890 400208
rect 341946 400152 346410 400208
rect 341885 400150 346410 400152
rect 348420 400150 355548 400210
rect 341885 400147 341951 400150
rect 348420 400074 348480 400150
rect 355542 400148 355548 400150
rect 355612 400148 355618 400212
rect 357382 400148 357388 400212
rect 357452 400210 357458 400212
rect 370446 400210 370452 400212
rect 357452 400150 370452 400210
rect 357452 400148 357458 400150
rect 370446 400148 370452 400150
rect 370516 400148 370522 400212
rect 354438 400074 354444 400076
rect 338070 400014 348480 400074
rect 351594 400014 354444 400074
rect 315389 399938 315455 399941
rect 338070 399938 338130 400014
rect 351594 399941 351654 400014
rect 354438 400012 354444 400014
rect 354508 400012 354514 400076
rect 354622 400012 354628 400076
rect 354692 400074 354698 400076
rect 354692 400014 355058 400074
rect 354692 400012 354698 400014
rect 343035 399940 343101 399941
rect 343771 399940 343837 399941
rect 343030 399938 343036 399940
rect 315389 399936 338130 399938
rect 315389 399880 315394 399936
rect 315450 399880 338130 399936
rect 315389 399878 338130 399880
rect 342944 399878 343036 399938
rect 315389 399875 315455 399878
rect 343030 399876 343036 399878
rect 343100 399876 343106 399940
rect 343766 399938 343772 399940
rect 343680 399878 343772 399938
rect 343766 399876 343772 399878
rect 343836 399876 343842 399940
rect 344323 399938 344389 399941
rect 344691 399940 344757 399941
rect 345059 399940 345125 399941
rect 344686 399938 344692 399940
rect 344142 399936 344389 399938
rect 344142 399880 344328 399936
rect 344384 399880 344389 399936
rect 344142 399878 344389 399880
rect 344600 399878 344692 399938
rect 343035 399875 343101 399876
rect 343771 399875 343837 399876
rect 344142 399805 344202 399878
rect 344323 399875 344389 399878
rect 344686 399876 344692 399878
rect 344756 399876 344762 399940
rect 345054 399876 345060 399940
rect 345124 399938 345130 399940
rect 345124 399878 345216 399938
rect 345124 399876 345130 399878
rect 345422 399876 345428 399940
rect 345492 399938 345498 399940
rect 345611 399938 345677 399941
rect 345492 399936 345677 399938
rect 345492 399880 345616 399936
rect 345672 399880 345677 399936
rect 345492 399878 345677 399880
rect 345492 399876 345498 399878
rect 344691 399875 344757 399876
rect 345059 399875 345125 399876
rect 345611 399875 345677 399878
rect 345790 399876 345796 399940
rect 345860 399938 345866 399940
rect 346071 399938 346137 399941
rect 346439 399938 346505 399941
rect 347267 399940 347333 399941
rect 347262 399938 347268 399940
rect 345860 399936 346137 399938
rect 345860 399880 346076 399936
rect 346132 399880 346137 399936
rect 345860 399878 346137 399880
rect 345860 399876 345866 399878
rect 346071 399875 346137 399878
rect 346304 399936 346505 399938
rect 346304 399880 346444 399936
rect 346500 399880 346505 399936
rect 346304 399878 346505 399880
rect 347176 399878 347268 399938
rect 301589 399802 301655 399805
rect 341885 399802 341951 399805
rect 301589 399800 341951 399802
rect 301589 399744 301594 399800
rect 301650 399744 341890 399800
rect 341946 399744 341951 399800
rect 301589 399742 341951 399744
rect 301589 399739 301655 399742
rect 341885 399739 341951 399742
rect 342294 399740 342300 399804
rect 342364 399802 342370 399804
rect 342943 399802 343009 399805
rect 343219 399804 343285 399805
rect 343214 399802 343220 399804
rect 342364 399800 343009 399802
rect 342364 399744 342948 399800
rect 343004 399744 343009 399800
rect 342364 399742 343009 399744
rect 343128 399742 343220 399802
rect 342364 399740 342370 399742
rect 342943 399739 343009 399742
rect 343214 399740 343220 399742
rect 343284 399740 343290 399804
rect 344093 399800 344202 399805
rect 344093 399744 344098 399800
rect 344154 399744 344202 399800
rect 344093 399742 344202 399744
rect 343219 399739 343285 399740
rect 344093 399739 344159 399742
rect 345238 399740 345244 399804
rect 345308 399802 345314 399804
rect 345887 399802 345953 399805
rect 345308 399800 345953 399802
rect 345308 399744 345892 399800
rect 345948 399744 345953 399800
rect 345308 399742 345953 399744
rect 346304 399804 346364 399878
rect 346439 399875 346505 399878
rect 347262 399876 347268 399878
rect 347332 399876 347338 399940
rect 347451 399936 347517 399941
rect 348003 399940 348069 399941
rect 348371 399940 348437 399941
rect 347451 399880 347456 399936
rect 347512 399880 347517 399936
rect 347267 399875 347333 399876
rect 347451 399875 347517 399880
rect 347630 399876 347636 399940
rect 347700 399938 347706 399940
rect 347998 399938 348004 399940
rect 347700 399907 347744 399938
rect 347700 399902 347793 399907
rect 347700 399876 347732 399902
rect 347454 399805 347514 399875
rect 347684 399846 347732 399876
rect 347788 399846 347793 399902
rect 347912 399878 348004 399938
rect 347998 399876 348004 399878
rect 348068 399876 348074 399940
rect 348366 399938 348372 399940
rect 348280 399878 348372 399938
rect 348366 399876 348372 399878
rect 348436 399876 348442 399940
rect 348550 399876 348556 399940
rect 348620 399938 348626 399940
rect 349199 399938 349265 399941
rect 350395 399940 350461 399941
rect 350390 399938 350396 399940
rect 348620 399936 349265 399938
rect 348620 399880 349204 399936
rect 349260 399880 349265 399936
rect 348620 399878 349265 399880
rect 350304 399878 350396 399938
rect 348620 399876 348626 399878
rect 348003 399875 348069 399876
rect 348371 399875 348437 399876
rect 349199 399875 349265 399878
rect 350390 399876 350396 399878
rect 350460 399876 350466 399940
rect 350574 399876 350580 399940
rect 350644 399938 350650 399940
rect 350763 399938 350829 399941
rect 350644 399936 350829 399938
rect 350644 399880 350768 399936
rect 350824 399880 350829 399936
rect 350644 399878 350829 399880
rect 350644 399876 350650 399878
rect 350395 399875 350461 399876
rect 350763 399875 350829 399878
rect 351039 399938 351105 399941
rect 351039 399936 351378 399938
rect 351039 399880 351044 399936
rect 351100 399880 351378 399936
rect 351039 399878 351378 399880
rect 351039 399875 351105 399878
rect 347684 399844 347793 399846
rect 347727 399841 347793 399844
rect 346304 399742 346348 399804
rect 345308 399740 345314 399742
rect 345887 399739 345953 399742
rect 346342 399740 346348 399742
rect 346412 399740 346418 399804
rect 347405 399800 347514 399805
rect 347405 399744 347410 399800
rect 347466 399744 347514 399800
rect 347405 399742 347514 399744
rect 347957 399802 348023 399805
rect 349107 399802 349173 399805
rect 350027 399804 350093 399805
rect 350022 399802 350028 399804
rect 347957 399800 349173 399802
rect 347957 399744 347962 399800
rect 348018 399744 349112 399800
rect 349168 399744 349173 399800
rect 347957 399742 349173 399744
rect 349936 399742 350028 399802
rect 347405 399739 347471 399742
rect 347957 399739 348023 399742
rect 349107 399739 349173 399742
rect 350022 399740 350028 399742
rect 350092 399740 350098 399804
rect 351318 399802 351378 399878
rect 351591 399936 351657 399941
rect 351591 399880 351596 399936
rect 351652 399880 351657 399936
rect 351591 399875 351657 399880
rect 351775 399938 351841 399941
rect 351775 399936 352114 399938
rect 351775 399880 351780 399936
rect 351836 399880 352114 399936
rect 351775 399878 352114 399880
rect 351775 399875 351841 399878
rect 351678 399802 351684 399804
rect 351318 399742 351684 399802
rect 351678 399740 351684 399742
rect 351748 399740 351754 399804
rect 351821 399802 351887 399805
rect 352054 399802 352114 399878
rect 352230 399876 352236 399940
rect 352300 399938 352306 399940
rect 353431 399938 353497 399941
rect 352300 399936 353497 399938
rect 352300 399880 353436 399936
rect 353492 399880 353497 399936
rect 352300 399878 353497 399880
rect 352300 399876 352306 399878
rect 353431 399875 353497 399878
rect 353702 399876 353708 399940
rect 353772 399938 353778 399940
rect 353983 399938 354049 399941
rect 353772 399936 354049 399938
rect 353772 399880 353988 399936
rect 354044 399880 354049 399936
rect 353772 399878 354049 399880
rect 353772 399876 353778 399878
rect 353983 399875 354049 399878
rect 354167 399938 354233 399941
rect 354622 399938 354628 399940
rect 354167 399936 354628 399938
rect 354167 399880 354172 399936
rect 354228 399880 354628 399936
rect 354167 399878 354628 399880
rect 354167 399875 354233 399878
rect 354622 399876 354628 399878
rect 354692 399876 354698 399940
rect 354998 399938 355058 400014
rect 355174 400012 355180 400076
rect 355244 400074 355250 400076
rect 364374 400074 364380 400076
rect 355244 400014 364380 400074
rect 355244 400012 355250 400014
rect 364374 400012 364380 400014
rect 364444 400012 364450 400076
rect 374126 400074 374132 400076
rect 365670 400014 374132 400074
rect 355363 399938 355429 399941
rect 354998 399936 355429 399938
rect 354998 399880 355368 399936
rect 355424 399880 355429 399936
rect 354998 399878 355429 399880
rect 355363 399875 355429 399878
rect 355542 399876 355548 399940
rect 355612 399938 355618 399940
rect 365670 399938 365730 400014
rect 374126 400012 374132 400014
rect 374196 400012 374202 400076
rect 376710 400014 377920 400074
rect 355612 399878 365730 399938
rect 365851 399936 365917 399941
rect 365851 399880 365856 399936
rect 365912 399880 365917 399936
rect 355612 399876 355618 399878
rect 365851 399875 365917 399880
rect 366311 399938 366377 399941
rect 366771 399940 366837 399941
rect 366582 399938 366588 399940
rect 366311 399936 366588 399938
rect 366311 399880 366316 399936
rect 366372 399880 366588 399936
rect 366311 399878 366588 399880
rect 366311 399875 366377 399878
rect 366582 399876 366588 399878
rect 366652 399876 366658 399940
rect 366766 399876 366772 399940
rect 366836 399938 366842 399940
rect 367691 399938 367757 399941
rect 368059 399940 368125 399941
rect 366836 399878 366928 399938
rect 367648 399936 367757 399938
rect 367648 399880 367696 399936
rect 367752 399880 367757 399936
rect 366836 399876 366842 399878
rect 366771 399875 366837 399876
rect 367648 399875 367757 399880
rect 368054 399876 368060 399940
rect 368124 399938 368130 399940
rect 368124 399878 368216 399938
rect 368124 399876 368130 399878
rect 368422 399876 368428 399940
rect 368492 399938 368498 399940
rect 369439 399938 369505 399941
rect 369715 399940 369781 399941
rect 371003 399940 371069 399941
rect 371739 399940 371805 399941
rect 369710 399938 369716 399940
rect 368492 399936 369505 399938
rect 368492 399880 369444 399936
rect 369500 399880 369505 399936
rect 368492 399878 369505 399880
rect 369624 399878 369716 399938
rect 368492 399876 368498 399878
rect 368059 399875 368125 399876
rect 369439 399875 369505 399878
rect 369710 399876 369716 399878
rect 369780 399876 369786 399940
rect 370998 399938 371004 399940
rect 370912 399878 371004 399938
rect 370998 399876 371004 399878
rect 371068 399876 371074 399940
rect 371182 399938 371188 399940
rect 371144 399876 371188 399938
rect 371252 399876 371258 399940
rect 371734 399938 371740 399940
rect 371371 399902 371437 399907
rect 369715 399875 369781 399876
rect 371003 399875 371069 399876
rect 352465 399804 352531 399805
rect 351821 399800 352114 399802
rect 351821 399744 351826 399800
rect 351882 399744 352114 399800
rect 351821 399742 352114 399744
rect 350027 399739 350093 399740
rect 351821 399739 351887 399742
rect 352414 399740 352420 399804
rect 352484 399802 352531 399804
rect 352879 399802 352945 399805
rect 353150 399802 353156 399804
rect 352484 399800 352576 399802
rect 352526 399744 352576 399800
rect 352484 399742 352576 399744
rect 352879 399800 353156 399802
rect 352879 399744 352884 399800
rect 352940 399744 353156 399800
rect 352879 399742 353156 399744
rect 352484 399740 352531 399742
rect 352465 399739 352531 399740
rect 352879 399739 352945 399742
rect 353150 399740 353156 399742
rect 353220 399740 353226 399804
rect 354070 399740 354076 399804
rect 354140 399802 354146 399804
rect 360510 399802 360516 399804
rect 354140 399742 360516 399802
rect 354140 399740 354146 399742
rect 360510 399740 360516 399742
rect 360580 399740 360586 399804
rect 360745 399802 360811 399805
rect 360878 399802 360884 399804
rect 360745 399800 360884 399802
rect 360745 399744 360750 399800
rect 360806 399744 360884 399800
rect 360745 399742 360884 399744
rect 360745 399739 360811 399742
rect 360878 399740 360884 399742
rect 360948 399740 360954 399804
rect 361711 399802 361777 399805
rect 362539 399804 362605 399805
rect 362534 399802 362540 399804
rect 361070 399800 361777 399802
rect 361070 399744 361716 399800
rect 361772 399744 361777 399800
rect 361070 399742 361777 399744
rect 362448 399742 362540 399802
rect 305729 399666 305795 399669
rect 355409 399668 355475 399669
rect 355174 399666 355180 399668
rect 305729 399664 355180 399666
rect 305729 399608 305734 399664
rect 305790 399608 355180 399664
rect 305729 399606 355180 399608
rect 305729 399603 305795 399606
rect 355174 399604 355180 399606
rect 355244 399604 355250 399668
rect 355358 399666 355364 399668
rect 355318 399606 355364 399666
rect 355428 399664 355475 399668
rect 355470 399608 355475 399664
rect 355358 399604 355364 399606
rect 355428 399604 355475 399608
rect 355542 399604 355548 399668
rect 355612 399666 355618 399668
rect 356881 399666 356947 399669
rect 355612 399664 356947 399666
rect 355612 399608 356886 399664
rect 356942 399608 356947 399664
rect 355612 399606 356947 399608
rect 355612 399604 355618 399606
rect 355409 399603 355475 399604
rect 356881 399603 356947 399606
rect 357617 399666 357683 399669
rect 357893 399666 357959 399669
rect 357617 399664 357959 399666
rect 357617 399608 357622 399664
rect 357678 399608 357898 399664
rect 357954 399608 357959 399664
rect 357617 399606 357959 399608
rect 357617 399603 357683 399606
rect 357893 399603 357959 399606
rect 358670 399604 358676 399668
rect 358740 399666 358746 399668
rect 359457 399666 359523 399669
rect 358740 399664 359523 399666
rect 358740 399608 359462 399664
rect 359518 399608 359523 399664
rect 358740 399606 359523 399608
rect 358740 399604 358746 399606
rect 359457 399603 359523 399606
rect 360694 399604 360700 399668
rect 360764 399666 360770 399668
rect 361070 399666 361130 399742
rect 361711 399739 361777 399742
rect 362534 399740 362540 399742
rect 362604 399740 362610 399804
rect 363086 399740 363092 399804
rect 363156 399802 363162 399804
rect 363919 399802 363985 399805
rect 363156 399800 363985 399802
rect 363156 399744 363924 399800
rect 363980 399744 363985 399800
rect 363156 399742 363985 399744
rect 363156 399740 363162 399742
rect 362539 399739 362605 399740
rect 363919 399739 363985 399742
rect 364190 399740 364196 399804
rect 364260 399802 364266 399804
rect 365854 399802 365914 399875
rect 367648 399805 367708 399875
rect 371144 399805 371204 399876
rect 371371 399846 371376 399902
rect 371432 399846 371437 399902
rect 371648 399878 371740 399938
rect 371734 399876 371740 399878
rect 371804 399876 371810 399940
rect 371923 399936 371989 399941
rect 372199 399938 372265 399941
rect 371923 399880 371928 399936
rect 371984 399880 371989 399936
rect 371739 399875 371805 399876
rect 371923 399875 371989 399880
rect 372156 399936 372265 399938
rect 372156 399880 372204 399936
rect 372260 399880 372265 399936
rect 372156 399875 372265 399880
rect 372567 399936 372633 399941
rect 372567 399880 372572 399936
rect 372628 399880 372633 399936
rect 372567 399875 372633 399880
rect 372935 399938 373001 399941
rect 372935 399936 373044 399938
rect 372935 399880 372940 399936
rect 372996 399880 373044 399936
rect 372935 399875 373044 399880
rect 371371 399841 371437 399846
rect 364260 399742 365914 399802
rect 366403 399802 366469 399805
rect 366582 399802 366588 399804
rect 366403 399800 366588 399802
rect 366403 399744 366408 399800
rect 366464 399744 366588 399800
rect 366403 399742 366588 399744
rect 364260 399740 364266 399742
rect 366403 399739 366469 399742
rect 366582 399740 366588 399742
rect 366652 399740 366658 399804
rect 367231 399802 367297 399805
rect 367502 399802 367508 399804
rect 367231 399800 367508 399802
rect 367231 399744 367236 399800
rect 367292 399744 367508 399800
rect 367231 399742 367508 399744
rect 367231 399739 367297 399742
rect 367502 399740 367508 399742
rect 367572 399740 367578 399804
rect 367645 399800 367711 399805
rect 367645 399744 367650 399800
rect 367706 399744 367711 399800
rect 367645 399739 367711 399744
rect 369894 399740 369900 399804
rect 369964 399802 369970 399804
rect 370819 399802 370885 399805
rect 369964 399800 370885 399802
rect 369964 399744 370824 399800
rect 370880 399744 370885 399800
rect 369964 399742 370885 399744
rect 369964 399740 369970 399742
rect 370819 399739 370885 399742
rect 371095 399800 371204 399805
rect 371095 399744 371100 399800
rect 371156 399744 371204 399800
rect 371095 399742 371204 399744
rect 371095 399739 371161 399742
rect 360764 399606 361130 399666
rect 365805 399666 365871 399669
rect 366214 399666 366220 399668
rect 365805 399664 366220 399666
rect 365805 399608 365810 399664
rect 365866 399608 366220 399664
rect 365805 399606 366220 399608
rect 360764 399604 360770 399606
rect 365805 399603 365871 399606
rect 366214 399604 366220 399606
rect 366284 399604 366290 399668
rect 366817 399666 366883 399669
rect 368238 399666 368244 399668
rect 366817 399664 368244 399666
rect 366817 399608 366822 399664
rect 366878 399608 368244 399664
rect 366817 399606 368244 399608
rect 366817 399603 366883 399606
rect 368238 399604 368244 399606
rect 368308 399604 368314 399668
rect 322473 399530 322539 399533
rect 322473 399528 369870 399530
rect 322473 399472 322478 399528
rect 322534 399472 369870 399528
rect 322473 399470 369870 399472
rect 322473 399467 322539 399470
rect 343950 399332 343956 399396
rect 344020 399394 344026 399396
rect 353293 399394 353359 399397
rect 344020 399392 353359 399394
rect 344020 399336 353298 399392
rect 353354 399336 353359 399392
rect 344020 399334 353359 399336
rect 344020 399332 344026 399334
rect 353293 399331 353359 399334
rect 353477 399394 353543 399397
rect 356145 399394 356211 399397
rect 357341 399396 357407 399397
rect 357341 399394 357388 399396
rect 353477 399392 356211 399394
rect 353477 399336 353482 399392
rect 353538 399336 356150 399392
rect 356206 399336 356211 399392
rect 353477 399334 356211 399336
rect 357296 399392 357388 399394
rect 357296 399336 357346 399392
rect 357296 399334 357388 399336
rect 353477 399331 353543 399334
rect 356145 399331 356211 399334
rect 357341 399332 357388 399334
rect 357452 399332 357458 399396
rect 358077 399394 358143 399397
rect 357942 399392 358143 399394
rect 357942 399336 358082 399392
rect 358138 399336 358143 399392
rect 357942 399334 358143 399336
rect 357341 399331 357407 399332
rect 357942 399261 358002 399334
rect 358077 399331 358143 399334
rect 364057 399394 364123 399397
rect 364609 399394 364675 399397
rect 364057 399392 364675 399394
rect 364057 399336 364062 399392
rect 364118 399336 364614 399392
rect 364670 399336 364675 399392
rect 364057 399334 364675 399336
rect 369810 399394 369870 399470
rect 370446 399468 370452 399532
rect 370516 399530 370522 399532
rect 371374 399530 371434 399841
rect 371550 399740 371556 399804
rect 371620 399802 371626 399804
rect 371926 399802 371986 399875
rect 372156 399805 372216 399875
rect 371620 399742 371986 399802
rect 372153 399800 372219 399805
rect 372383 399802 372449 399805
rect 372153 399744 372158 399800
rect 372214 399744 372219 399800
rect 371620 399740 371626 399742
rect 372153 399739 372219 399744
rect 372340 399800 372449 399802
rect 372340 399744 372388 399800
rect 372444 399744 372449 399800
rect 372340 399739 372449 399744
rect 372570 399802 372630 399875
rect 372838 399802 372844 399804
rect 372570 399742 372844 399802
rect 372838 399740 372844 399742
rect 372908 399740 372914 399804
rect 372340 399668 372400 399739
rect 372984 399669 373044 399875
rect 373947 399902 374013 399907
rect 373947 399846 373952 399902
rect 374008 399846 374013 399902
rect 373947 399841 374013 399846
rect 374131 399902 374197 399907
rect 374131 399846 374136 399902
rect 374192 399846 374197 399902
rect 374310 399876 374316 399940
rect 374380 399938 374386 399940
rect 375327 399938 375393 399941
rect 376247 399938 376313 399941
rect 374380 399936 375393 399938
rect 374380 399880 375332 399936
rect 375388 399880 375393 399936
rect 374380 399878 375393 399880
rect 374380 399876 374386 399878
rect 375327 399875 375393 399878
rect 375560 399936 376313 399938
rect 375560 399880 376252 399936
rect 376308 399880 376313 399936
rect 375560 399878 376313 399880
rect 374131 399841 374197 399846
rect 373395 399802 373461 399805
rect 373214 399800 373461 399802
rect 373214 399744 373400 399800
rect 373456 399744 373461 399800
rect 373214 399742 373461 399744
rect 372286 399604 372292 399668
rect 372356 399606 372400 399668
rect 372981 399664 373047 399669
rect 372981 399608 372986 399664
rect 373042 399608 373047 399664
rect 372356 399604 372362 399606
rect 372981 399603 373047 399608
rect 370516 399470 371434 399530
rect 372981 399530 373047 399533
rect 373214 399530 373274 399742
rect 373395 399739 373461 399742
rect 373349 399666 373415 399669
rect 373950 399666 374010 399841
rect 374134 399669 374194 399841
rect 374867 399804 374933 399805
rect 374862 399802 374868 399804
rect 374776 399742 374868 399802
rect 374862 399740 374868 399742
rect 374932 399740 374938 399804
rect 375560 399802 375620 399878
rect 376247 399875 376313 399878
rect 375054 399742 375620 399802
rect 374867 399739 374933 399740
rect 373349 399664 374010 399666
rect 373349 399608 373354 399664
rect 373410 399608 374010 399664
rect 373349 399606 374010 399608
rect 374085 399664 374194 399669
rect 374085 399608 374090 399664
rect 374146 399608 374194 399664
rect 374085 399606 374194 399608
rect 373349 399603 373415 399606
rect 374085 399603 374151 399606
rect 372981 399528 373274 399530
rect 372981 399472 372986 399528
rect 373042 399472 373274 399528
rect 372981 399470 373274 399472
rect 374821 399530 374887 399533
rect 375054 399530 375114 399742
rect 376710 399533 376770 400014
rect 377860 399941 377920 400014
rect 376983 399938 377049 399941
rect 374821 399528 375114 399530
rect 374821 399472 374826 399528
rect 374882 399472 375114 399528
rect 374821 399470 375114 399472
rect 376661 399528 376770 399533
rect 376661 399472 376666 399528
rect 376722 399472 376770 399528
rect 376661 399470 376770 399472
rect 376940 399936 377049 399938
rect 376940 399880 376988 399936
rect 377044 399880 377049 399936
rect 376940 399875 377049 399880
rect 377259 399936 377325 399941
rect 377627 399940 377693 399941
rect 377622 399938 377628 399940
rect 377259 399880 377264 399936
rect 377320 399880 377325 399936
rect 377259 399875 377325 399880
rect 377536 399878 377628 399938
rect 377622 399876 377628 399878
rect 377692 399876 377698 399940
rect 377860 399936 377969 399941
rect 377860 399880 377908 399936
rect 377964 399880 377969 399936
rect 377860 399878 377969 399880
rect 378228 399938 378288 400286
rect 387793 400283 387859 400286
rect 378358 400148 378364 400212
rect 378428 400210 378434 400212
rect 378428 400150 380588 400210
rect 378428 400148 378434 400150
rect 379278 400012 379284 400076
rect 379348 400074 379354 400076
rect 379348 400014 380266 400074
rect 379348 400012 379354 400014
rect 380206 399941 380266 400014
rect 378363 399938 378429 399941
rect 378823 399938 378889 399941
rect 378228 399936 378429 399938
rect 378228 399880 378368 399936
rect 378424 399880 378429 399936
rect 378228 399878 378429 399880
rect 377627 399875 377693 399876
rect 377903 399875 377969 399878
rect 378363 399875 378429 399878
rect 378780 399936 378889 399938
rect 378780 399880 378828 399936
rect 378884 399880 378889 399936
rect 378780 399875 378889 399880
rect 379094 399876 379100 399940
rect 379164 399938 379170 399940
rect 379283 399938 379349 399941
rect 379164 399936 379349 399938
rect 379164 399880 379288 399936
rect 379344 399880 379349 399936
rect 379164 399878 379349 399880
rect 379164 399876 379170 399878
rect 379283 399875 379349 399878
rect 379467 399936 379533 399941
rect 379927 399938 379993 399941
rect 379467 399880 379472 399936
rect 379528 399880 379533 399936
rect 379884 399936 379993 399938
rect 379467 399875 379533 399880
rect 379651 399902 379717 399907
rect 376940 399530 377000 399875
rect 377262 399666 377322 399875
rect 378174 399740 378180 399804
rect 378244 399802 378250 399804
rect 378780 399802 378840 399875
rect 378244 399742 378840 399802
rect 378244 399740 378250 399742
rect 377857 399666 377923 399669
rect 377262 399664 377923 399666
rect 377262 399608 377862 399664
rect 377918 399608 377923 399664
rect 377262 399606 377923 399608
rect 377857 399603 377923 399606
rect 378961 399666 379027 399669
rect 379470 399666 379530 399875
rect 379651 399846 379656 399902
rect 379712 399846 379717 399902
rect 379651 399841 379717 399846
rect 379884 399880 379932 399936
rect 379988 399880 379993 399936
rect 379884 399875 379993 399880
rect 380203 399936 380269 399941
rect 380203 399880 380208 399936
rect 380264 399880 380269 399936
rect 380203 399875 380269 399880
rect 380528 399938 380588 400150
rect 381670 400012 381676 400076
rect 381740 400074 381746 400076
rect 390001 400074 390067 400077
rect 381740 400014 384820 400074
rect 381740 400012 381746 400014
rect 381031 399938 381097 399941
rect 380528 399936 381097 399938
rect 380528 399880 381036 399936
rect 381092 399880 381097 399936
rect 380528 399878 381097 399880
rect 381031 399875 381097 399878
rect 381675 399936 381741 399941
rect 381675 399880 381680 399936
rect 381736 399880 381741 399936
rect 381675 399875 381741 399880
rect 382406 399876 382412 399940
rect 382476 399938 382482 399940
rect 382687 399938 382753 399941
rect 384343 399938 384409 399941
rect 382476 399936 382753 399938
rect 382476 399880 382692 399936
rect 382748 399880 382753 399936
rect 382476 399878 382753 399880
rect 382476 399876 382482 399878
rect 382687 399875 382753 399878
rect 383840 399936 384409 399938
rect 383840 399880 384348 399936
rect 384404 399880 384409 399936
rect 383840 399878 384409 399880
rect 384760 399938 384820 400014
rect 385358 400072 390067 400074
rect 385358 400016 390006 400072
rect 390062 400016 390067 400072
rect 385358 400014 390067 400016
rect 385358 399941 385418 400014
rect 390001 400011 390067 400014
rect 384895 399938 384961 399941
rect 384760 399936 384961 399938
rect 384760 399880 384900 399936
rect 384956 399880 384961 399936
rect 384760 399878 384961 399880
rect 378961 399664 379530 399666
rect 378961 399608 378966 399664
rect 379022 399608 379530 399664
rect 378961 399606 379530 399608
rect 378961 399603 379027 399606
rect 378225 399530 378291 399533
rect 378593 399532 378659 399533
rect 378542 399530 378548 399532
rect 376940 399528 378291 399530
rect 376940 399472 378230 399528
rect 378286 399472 378291 399528
rect 376940 399470 378291 399472
rect 378502 399470 378548 399530
rect 378612 399528 378659 399532
rect 378654 399472 378659 399528
rect 370516 399468 370522 399470
rect 372981 399467 373047 399470
rect 374821 399467 374887 399470
rect 376661 399467 376727 399470
rect 378225 399467 378291 399470
rect 378542 399468 378548 399470
rect 378612 399468 378659 399472
rect 379654 399530 379714 399841
rect 379884 399804 379944 399875
rect 379830 399740 379836 399804
rect 379900 399742 379944 399804
rect 380111 399802 380177 399805
rect 380111 399800 380312 399802
rect 380111 399744 380116 399800
rect 380172 399744 380312 399800
rect 380111 399742 380312 399744
rect 379900 399740 379906 399742
rect 380111 399739 380177 399742
rect 379973 399666 380039 399669
rect 380252 399666 380312 399742
rect 379973 399664 380312 399666
rect 379973 399608 379978 399664
rect 380034 399608 380312 399664
rect 379973 399606 380312 399608
rect 381169 399666 381235 399669
rect 381678 399666 381738 399875
rect 382963 399800 383029 399805
rect 382963 399744 382968 399800
rect 383024 399744 383029 399800
rect 382963 399739 383029 399744
rect 383147 399800 383213 399805
rect 383147 399744 383152 399800
rect 383208 399744 383213 399800
rect 383147 399739 383213 399744
rect 381169 399664 381738 399666
rect 381169 399608 381174 399664
rect 381230 399608 381738 399664
rect 381169 399606 381738 399608
rect 379973 399603 380039 399606
rect 381169 399603 381235 399606
rect 380157 399530 380223 399533
rect 379654 399528 380223 399530
rect 379654 399472 380162 399528
rect 380218 399472 380223 399528
rect 379654 399470 380223 399472
rect 378593 399467 378659 399468
rect 380157 399467 380223 399470
rect 382825 399530 382891 399533
rect 382966 399530 383026 399739
rect 383150 399533 383210 399739
rect 383840 399669 383900 399878
rect 384343 399875 384409 399878
rect 384895 399875 384961 399878
rect 385171 399936 385237 399941
rect 385171 399880 385176 399936
rect 385232 399880 385237 399936
rect 385171 399875 385237 399880
rect 385355 399936 385421 399941
rect 385355 399880 385360 399936
rect 385416 399880 385421 399936
rect 385355 399875 385421 399880
rect 386367 399938 386433 399941
rect 390829 399938 390895 399941
rect 386367 399936 390895 399938
rect 386367 399880 386372 399936
rect 386428 399880 390834 399936
rect 390890 399880 390895 399936
rect 386367 399878 390895 399880
rect 386367 399875 386433 399878
rect 390829 399875 390895 399878
rect 384619 399834 384685 399839
rect 383975 399802 384041 399805
rect 383975 399800 384498 399802
rect 383975 399744 383980 399800
rect 384036 399744 384498 399800
rect 384619 399778 384624 399834
rect 384680 399778 384685 399834
rect 384619 399773 384685 399778
rect 383975 399742 384498 399744
rect 383975 399739 384041 399742
rect 383837 399664 383903 399669
rect 383837 399608 383842 399664
rect 383898 399608 383903 399664
rect 383837 399603 383903 399608
rect 382825 399528 383026 399530
rect 382825 399472 382830 399528
rect 382886 399472 383026 399528
rect 382825 399470 383026 399472
rect 383101 399528 383210 399533
rect 383101 399472 383106 399528
rect 383162 399472 383210 399528
rect 383101 399470 383210 399472
rect 382825 399467 382891 399470
rect 383101 399467 383167 399470
rect 382222 399394 382228 399396
rect 369810 399334 382228 399394
rect 364057 399331 364123 399334
rect 364609 399331 364675 399334
rect 382222 399332 382228 399334
rect 382292 399332 382298 399396
rect 384438 399394 384498 399742
rect 384622 399669 384682 399773
rect 385174 399669 385234 399875
rect 385723 399834 385789 399839
rect 385723 399778 385728 399834
rect 385784 399778 385789 399834
rect 385723 399773 385789 399778
rect 386827 399800 386893 399805
rect 384622 399664 384731 399669
rect 384622 399608 384670 399664
rect 384726 399608 384731 399664
rect 384622 399606 384731 399608
rect 385174 399664 385283 399669
rect 385174 399608 385222 399664
rect 385278 399608 385283 399664
rect 385174 399606 385283 399608
rect 384665 399603 384731 399606
rect 385217 399603 385283 399606
rect 385726 399530 385786 399773
rect 386827 399744 386832 399800
rect 386888 399744 386893 399800
rect 386827 399739 386893 399744
rect 386830 399666 386890 399739
rect 387149 399666 387215 399669
rect 386830 399664 387215 399666
rect 386830 399608 387154 399664
rect 387210 399608 387215 399664
rect 386830 399606 387215 399608
rect 387149 399603 387215 399606
rect 388161 399530 388227 399533
rect 385726 399528 388227 399530
rect 385726 399472 388166 399528
rect 388222 399472 388227 399528
rect 385726 399470 388227 399472
rect 388161 399467 388227 399470
rect 392209 399394 392275 399397
rect 384438 399392 392275 399394
rect 384438 399336 392214 399392
rect 392270 399336 392275 399392
rect 384438 399334 392275 399336
rect 392209 399331 392275 399334
rect 347313 399258 347379 399261
rect 335310 399256 347379 399258
rect 335310 399200 347318 399256
rect 347374 399200 347379 399256
rect 335310 399198 347379 399200
rect 289118 398924 289124 398988
rect 289188 398986 289194 398988
rect 335310 398986 335370 399198
rect 347313 399195 347379 399198
rect 347773 399258 347839 399261
rect 349102 399258 349108 399260
rect 347773 399256 349108 399258
rect 347773 399200 347778 399256
rect 347834 399200 349108 399256
rect 347773 399198 349108 399200
rect 347773 399195 347839 399198
rect 349102 399196 349108 399198
rect 349172 399196 349178 399260
rect 353334 399196 353340 399260
rect 353404 399258 353410 399260
rect 354397 399258 354463 399261
rect 353404 399256 354463 399258
rect 353404 399200 354402 399256
rect 354458 399200 354463 399256
rect 353404 399198 354463 399200
rect 353404 399196 353410 399198
rect 354397 399195 354463 399198
rect 354581 399258 354647 399261
rect 354581 399256 356070 399258
rect 354581 399200 354586 399256
rect 354642 399200 356070 399256
rect 354581 399198 356070 399200
rect 354581 399195 354647 399198
rect 346761 399122 346827 399125
rect 348417 399122 348483 399125
rect 289188 398926 335370 398986
rect 340830 399062 346226 399122
rect 289188 398924 289194 398926
rect 310278 398788 310284 398852
rect 310348 398850 310354 398852
rect 340830 398850 340890 399062
rect 341425 398986 341491 398989
rect 346166 398986 346226 399062
rect 346761 399120 348483 399122
rect 346761 399064 346766 399120
rect 346822 399064 348422 399120
rect 348478 399064 348483 399120
rect 346761 399062 348483 399064
rect 346761 399059 346827 399062
rect 348417 399059 348483 399062
rect 348693 399122 348759 399125
rect 354029 399122 354095 399125
rect 348693 399120 354095 399122
rect 348693 399064 348698 399120
rect 348754 399064 354034 399120
rect 354090 399064 354095 399120
rect 348693 399062 354095 399064
rect 356010 399122 356070 399198
rect 357893 399256 358002 399261
rect 357893 399200 357898 399256
rect 357954 399200 358002 399256
rect 357893 399198 358002 399200
rect 357893 399195 357959 399198
rect 358118 399196 358124 399260
rect 358188 399258 358194 399260
rect 358261 399258 358327 399261
rect 364885 399258 364951 399261
rect 358188 399256 358327 399258
rect 358188 399200 358266 399256
rect 358322 399200 358327 399256
rect 358188 399198 358327 399200
rect 358188 399196 358194 399198
rect 358261 399195 358327 399198
rect 358448 399256 364951 399258
rect 358448 399200 364890 399256
rect 364946 399200 364951 399256
rect 358448 399198 364951 399200
rect 358448 399122 358508 399198
rect 364885 399195 364951 399198
rect 367553 399258 367619 399261
rect 373206 399258 373212 399260
rect 367553 399256 373212 399258
rect 367553 399200 367558 399256
rect 367614 399200 373212 399256
rect 367553 399198 373212 399200
rect 367553 399195 367619 399198
rect 373206 399196 373212 399198
rect 373276 399196 373282 399260
rect 373942 399196 373948 399260
rect 374012 399258 374018 399260
rect 374453 399258 374519 399261
rect 374012 399256 374519 399258
rect 374012 399200 374458 399256
rect 374514 399200 374519 399256
rect 374012 399198 374519 399200
rect 374012 399196 374018 399198
rect 374453 399195 374519 399198
rect 379237 399258 379303 399261
rect 380801 399258 380867 399261
rect 379237 399256 380867 399258
rect 379237 399200 379242 399256
rect 379298 399200 380806 399256
rect 380862 399200 380867 399256
rect 379237 399198 380867 399200
rect 379237 399195 379303 399198
rect 380801 399195 380867 399198
rect 368422 399122 368428 399124
rect 356010 399062 358508 399122
rect 360150 399062 368428 399122
rect 348693 399059 348759 399062
rect 354029 399059 354095 399062
rect 360150 398986 360210 399062
rect 368422 399060 368428 399062
rect 368492 399060 368498 399124
rect 370497 399122 370563 399125
rect 371734 399122 371740 399124
rect 370497 399120 371740 399122
rect 370497 399064 370502 399120
rect 370558 399064 371740 399120
rect 370497 399062 371740 399064
rect 370497 399059 370563 399062
rect 371734 399060 371740 399062
rect 371804 399060 371810 399124
rect 376937 399122 377003 399125
rect 377305 399122 377371 399125
rect 376937 399120 377371 399122
rect 376937 399064 376942 399120
rect 376998 399064 377310 399120
rect 377366 399064 377371 399120
rect 376937 399062 377371 399064
rect 376937 399059 377003 399062
rect 377305 399059 377371 399062
rect 364057 398986 364123 398989
rect 341425 398984 345858 398986
rect 341425 398928 341430 398984
rect 341486 398928 345858 398984
rect 341425 398926 345858 398928
rect 346166 398926 360210 398986
rect 361668 398984 364123 398986
rect 361668 398928 364062 398984
rect 364118 398928 364123 398984
rect 361668 398926 364123 398928
rect 341425 398923 341491 398926
rect 310348 398790 331230 398850
rect 310348 398788 310354 398790
rect 331170 398714 331230 398790
rect 340646 398790 340890 398850
rect 341885 398850 341951 398853
rect 345657 398850 345723 398853
rect 341885 398848 345723 398850
rect 341885 398792 341890 398848
rect 341946 398792 345662 398848
rect 345718 398792 345723 398848
rect 341885 398790 345723 398792
rect 340646 398714 340706 398790
rect 341885 398787 341951 398790
rect 345657 398787 345723 398790
rect 331170 398654 340706 398714
rect 343173 398714 343239 398717
rect 344737 398714 344803 398717
rect 343173 398712 344803 398714
rect 343173 398656 343178 398712
rect 343234 398656 344742 398712
rect 344798 398656 344803 398712
rect 343173 398654 344803 398656
rect 345798 398714 345858 398926
rect 347773 398850 347839 398853
rect 356329 398850 356395 398853
rect 347773 398848 356395 398850
rect 347773 398792 347778 398848
rect 347834 398792 356334 398848
rect 356390 398792 356395 398848
rect 347773 398790 356395 398792
rect 347773 398787 347839 398790
rect 356329 398787 356395 398790
rect 357157 398850 357223 398853
rect 361668 398850 361728 398926
rect 364057 398923 364123 398926
rect 371734 398924 371740 398988
rect 371804 398986 371810 398988
rect 375465 398986 375531 398989
rect 371804 398984 375531 398986
rect 371804 398928 375470 398984
rect 375526 398928 375531 398984
rect 371804 398926 375531 398928
rect 371804 398924 371810 398926
rect 375465 398923 375531 398926
rect 357157 398848 361728 398850
rect 357157 398792 357162 398848
rect 357218 398792 361728 398848
rect 357157 398790 361728 398792
rect 357157 398787 357223 398790
rect 355777 398714 355843 398717
rect 345798 398712 355843 398714
rect 345798 398656 355782 398712
rect 355838 398656 355843 398712
rect 345798 398654 355843 398656
rect 343173 398651 343239 398654
rect 344737 398651 344803 398654
rect 355777 398651 355843 398654
rect 365110 398652 365116 398716
rect 365180 398714 365186 398716
rect 370998 398714 371004 398716
rect 365180 398654 371004 398714
rect 365180 398652 365186 398654
rect 370998 398652 371004 398654
rect 371068 398652 371074 398716
rect 334157 398578 334223 398581
rect 344645 398578 344711 398581
rect 334157 398576 344711 398578
rect 334157 398520 334162 398576
rect 334218 398520 344650 398576
rect 344706 398520 344711 398576
rect 334157 398518 344711 398520
rect 334157 398515 334223 398518
rect 344645 398515 344711 398518
rect 350758 398516 350764 398580
rect 350828 398578 350834 398580
rect 351545 398578 351611 398581
rect 350828 398576 351611 398578
rect 350828 398520 351550 398576
rect 351606 398520 351611 398576
rect 350828 398518 351611 398520
rect 350828 398516 350834 398518
rect 351545 398515 351611 398518
rect 330937 398442 331003 398445
rect 371233 398442 371299 398445
rect 330937 398440 371299 398442
rect 330937 398384 330942 398440
rect 330998 398384 371238 398440
rect 371294 398384 371299 398440
rect 330937 398382 371299 398384
rect 330937 398379 331003 398382
rect 371233 398379 371299 398382
rect 264881 398306 264947 398309
rect 334157 398306 334223 398309
rect 264881 398304 334223 398306
rect 264881 398248 264886 398304
rect 264942 398248 334162 398304
rect 334218 398248 334223 398304
rect 264881 398246 334223 398248
rect 264881 398243 264947 398246
rect 334157 398243 334223 398246
rect 340229 398306 340295 398309
rect 348693 398306 348759 398309
rect 340229 398304 348759 398306
rect 340229 398248 340234 398304
rect 340290 398248 348698 398304
rect 348754 398248 348759 398304
rect 340229 398246 348759 398248
rect 340229 398243 340295 398246
rect 348693 398243 348759 398246
rect 352414 398244 352420 398308
rect 352484 398306 352490 398308
rect 369485 398306 369551 398309
rect 352484 398304 369551 398306
rect 352484 398248 369490 398304
rect 369546 398248 369551 398304
rect 352484 398246 369551 398248
rect 352484 398244 352490 398246
rect 369485 398243 369551 398246
rect 256601 398170 256667 398173
rect 343214 398170 343220 398172
rect 256601 398168 343220 398170
rect 256601 398112 256606 398168
rect 256662 398112 343220 398168
rect 256601 398110 343220 398112
rect 256601 398107 256667 398110
rect 343214 398108 343220 398110
rect 343284 398108 343290 398172
rect 344645 398170 344711 398173
rect 347998 398170 348004 398172
rect 344645 398168 348004 398170
rect 344645 398112 344650 398168
rect 344706 398112 348004 398168
rect 344645 398110 348004 398112
rect 344645 398107 344711 398110
rect 347998 398108 348004 398110
rect 348068 398108 348074 398172
rect 357566 398108 357572 398172
rect 357636 398170 357642 398172
rect 358445 398170 358511 398173
rect 357636 398168 358511 398170
rect 357636 398112 358450 398168
rect 358506 398112 358511 398168
rect 357636 398110 358511 398112
rect 357636 398108 357642 398110
rect 358445 398107 358511 398110
rect 384757 398170 384823 398173
rect 391933 398170 391999 398173
rect 384757 398168 391999 398170
rect 384757 398112 384762 398168
rect 384818 398112 391938 398168
rect 391994 398112 391999 398168
rect 384757 398110 391999 398112
rect 384757 398107 384823 398110
rect 391933 398107 391999 398110
rect 259361 398034 259427 398037
rect 345381 398034 345447 398037
rect 259361 398032 345447 398034
rect 259361 397976 259366 398032
rect 259422 397976 345386 398032
rect 345442 397976 345447 398032
rect 259361 397974 345447 397976
rect 259361 397971 259427 397974
rect 345381 397971 345447 397974
rect 355174 397972 355180 398036
rect 355244 398034 355250 398036
rect 357525 398034 357591 398037
rect 355244 398032 357591 398034
rect 355244 397976 357530 398032
rect 357586 397976 357591 398032
rect 355244 397974 357591 397976
rect 355244 397972 355250 397974
rect 357525 397971 357591 397974
rect 368974 397972 368980 398036
rect 369044 398034 369050 398036
rect 376293 398034 376359 398037
rect 369044 398032 376359 398034
rect 369044 397976 376298 398032
rect 376354 397976 376359 398032
rect 369044 397974 376359 397976
rect 369044 397972 369050 397974
rect 376293 397971 376359 397974
rect 357382 397836 357388 397900
rect 357452 397898 357458 397900
rect 358353 397898 358419 397901
rect 357452 397896 358419 397898
rect 357452 397840 358358 397896
rect 358414 397840 358419 397896
rect 357452 397838 358419 397840
rect 357452 397836 357458 397838
rect 358353 397835 358419 397838
rect 375966 397836 375972 397900
rect 376036 397898 376042 397900
rect 380709 397898 380775 397901
rect 376036 397896 380775 397898
rect 376036 397840 380714 397896
rect 380770 397840 380775 397896
rect 376036 397838 380775 397840
rect 376036 397836 376042 397838
rect 380709 397835 380775 397838
rect 360326 397700 360332 397764
rect 360396 397762 360402 397764
rect 361389 397762 361455 397765
rect 360396 397760 361455 397762
rect 360396 397704 361394 397760
rect 361450 397704 361455 397760
rect 360396 397702 361455 397704
rect 360396 397700 360402 397702
rect 361389 397699 361455 397702
rect 377254 397700 377260 397764
rect 377324 397762 377330 397764
rect 381813 397762 381879 397765
rect 377324 397760 381879 397762
rect 377324 397704 381818 397760
rect 381874 397704 381879 397760
rect 377324 397702 381879 397704
rect 377324 397700 377330 397702
rect 381813 397699 381879 397702
rect 336273 397626 336339 397629
rect 365621 397626 365687 397629
rect 372245 397628 372311 397629
rect 372245 397626 372292 397628
rect 336273 397624 365687 397626
rect -960 397490 480 397580
rect 336273 397568 336278 397624
rect 336334 397568 365626 397624
rect 365682 397568 365687 397624
rect 336273 397566 365687 397568
rect 372200 397624 372292 397626
rect 372200 397568 372250 397624
rect 372200 397566 372292 397568
rect 336273 397563 336339 397566
rect 365621 397563 365687 397566
rect 372245 397564 372292 397566
rect 372356 397564 372362 397628
rect 380934 397564 380940 397628
rect 381004 397626 381010 397628
rect 382089 397626 382155 397629
rect 381004 397624 382155 397626
rect 381004 397568 382094 397624
rect 382150 397568 382155 397624
rect 381004 397566 382155 397568
rect 381004 397564 381010 397566
rect 372245 397563 372311 397564
rect 382089 397563 382155 397566
rect 382222 397564 382228 397628
rect 382292 397626 382298 397628
rect 383469 397626 383535 397629
rect 382292 397624 383535 397626
rect 382292 397568 383474 397624
rect 383530 397568 383535 397624
rect 382292 397566 383535 397568
rect 382292 397564 382298 397566
rect 383469 397563 383535 397566
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 350390 397428 350396 397492
rect 350460 397490 350466 397492
rect 350533 397490 350599 397493
rect 350460 397488 350599 397490
rect 350460 397432 350538 397488
rect 350594 397432 350599 397488
rect 350460 397430 350599 397432
rect 350460 397428 350466 397430
rect 350533 397427 350599 397430
rect 352925 397490 352991 397493
rect 356513 397492 356579 397493
rect 353150 397490 353156 397492
rect 352925 397488 353156 397490
rect 352925 397432 352930 397488
rect 352986 397432 353156 397488
rect 352925 397430 353156 397432
rect 352925 397427 352991 397430
rect 353150 397428 353156 397430
rect 353220 397428 353226 397492
rect 356462 397490 356468 397492
rect 356422 397430 356468 397490
rect 356532 397488 356579 397492
rect 356574 397432 356579 397488
rect 356462 397428 356468 397430
rect 356532 397428 356579 397432
rect 356513 397427 356579 397428
rect 357433 397490 357499 397493
rect 358118 397490 358124 397492
rect 357433 397488 358124 397490
rect 357433 397432 357438 397488
rect 357494 397432 358124 397488
rect 357433 397430 358124 397432
rect 357433 397427 357499 397430
rect 358118 397428 358124 397430
rect 358188 397428 358194 397492
rect 359406 397428 359412 397492
rect 359476 397490 359482 397492
rect 372838 397490 372844 397492
rect 359476 397430 372844 397490
rect 359476 397428 359482 397430
rect 372838 397428 372844 397430
rect 372908 397428 372914 397492
rect 382038 397428 382044 397492
rect 382108 397490 382114 397492
rect 382273 397490 382339 397493
rect 382108 397488 382339 397490
rect 382108 397432 382278 397488
rect 382334 397432 382339 397488
rect 382108 397430 382339 397432
rect 382108 397428 382114 397430
rect 382273 397427 382339 397430
rect 337469 397354 337535 397357
rect 358077 397354 358143 397357
rect 337469 397352 358143 397354
rect 337469 397296 337474 397352
rect 337530 397296 358082 397352
rect 358138 397296 358143 397352
rect 337469 397294 358143 397296
rect 337469 397291 337535 397294
rect 358077 397291 358143 397294
rect 364374 397292 364380 397356
rect 364444 397354 364450 397356
rect 365253 397354 365319 397357
rect 367921 397356 367987 397357
rect 367870 397354 367876 397356
rect 364444 397352 365319 397354
rect 364444 397296 365258 397352
rect 365314 397296 365319 397352
rect 364444 397294 365319 397296
rect 367830 397294 367876 397354
rect 367940 397352 367987 397356
rect 367982 397296 367987 397352
rect 364444 397292 364450 397294
rect 365253 397291 365319 397294
rect 367870 397292 367876 397294
rect 367940 397292 367987 397296
rect 369158 397292 369164 397356
rect 369228 397354 369234 397356
rect 373073 397354 373139 397357
rect 369228 397352 373139 397354
rect 369228 397296 373078 397352
rect 373134 397296 373139 397352
rect 369228 397294 373139 397296
rect 369228 397292 369234 397294
rect 367921 397291 367987 397292
rect 373073 397291 373139 397294
rect 374913 397354 374979 397357
rect 382457 397356 382523 397357
rect 375414 397354 375420 397356
rect 374913 397352 375420 397354
rect 374913 397296 374918 397352
rect 374974 397296 375420 397352
rect 374913 397294 375420 397296
rect 374913 397291 374979 397294
rect 375414 397292 375420 397294
rect 375484 397292 375490 397356
rect 382406 397292 382412 397356
rect 382476 397354 382523 397356
rect 382476 397352 382568 397354
rect 382518 397296 382568 397352
rect 382476 397294 382568 397296
rect 382476 397292 382523 397294
rect 382774 397292 382780 397356
rect 382844 397354 382850 397356
rect 385401 397354 385467 397357
rect 382844 397352 385467 397354
rect 382844 397296 385406 397352
rect 385462 397296 385467 397352
rect 382844 397294 385467 397296
rect 382844 397292 382850 397294
rect 382457 397291 382523 397292
rect 385401 397291 385467 397294
rect 283414 397156 283420 397220
rect 283484 397218 283490 397220
rect 295333 397218 295399 397221
rect 283484 397216 295399 397218
rect 283484 397160 295338 397216
rect 295394 397160 295399 397216
rect 283484 397158 295399 397160
rect 283484 397156 283490 397158
rect 295333 397155 295399 397158
rect 333237 397218 333303 397221
rect 353477 397218 353543 397221
rect 333237 397216 353543 397218
rect 333237 397160 333242 397216
rect 333298 397160 353482 397216
rect 353538 397160 353543 397216
rect 333237 397158 353543 397160
rect 333237 397155 333303 397158
rect 353477 397155 353543 397158
rect 358118 397156 358124 397220
rect 358188 397218 358194 397220
rect 369025 397218 369091 397221
rect 372337 397220 372403 397221
rect 372286 397218 372292 397220
rect 358188 397216 369091 397218
rect 358188 397160 369030 397216
rect 369086 397160 369091 397216
rect 358188 397158 369091 397160
rect 372246 397158 372292 397218
rect 372356 397216 372403 397220
rect 372398 397160 372403 397216
rect 358188 397156 358194 397158
rect 369025 397155 369091 397158
rect 372286 397156 372292 397158
rect 372356 397156 372403 397160
rect 372337 397155 372403 397156
rect 274173 397082 274239 397085
rect 355542 397082 355548 397084
rect 274173 397080 355548 397082
rect 274173 397024 274178 397080
rect 274234 397024 355548 397080
rect 274173 397022 355548 397024
rect 274173 397019 274239 397022
rect 355542 397020 355548 397022
rect 355612 397020 355618 397084
rect 357014 397020 357020 397084
rect 357084 397082 357090 397084
rect 374310 397082 374316 397084
rect 357084 397022 374316 397082
rect 357084 397020 357090 397022
rect 374310 397020 374316 397022
rect 374380 397020 374386 397084
rect 270125 396946 270191 396949
rect 356973 396946 357039 396949
rect 358905 396948 358971 396949
rect 358854 396946 358860 396948
rect 270125 396944 357039 396946
rect 270125 396888 270130 396944
rect 270186 396888 356978 396944
rect 357034 396888 357039 396944
rect 270125 396886 357039 396888
rect 358814 396886 358860 396946
rect 358924 396944 358971 396948
rect 358966 396888 358971 396944
rect 270125 396883 270191 396886
rect 356973 396883 357039 396886
rect 358854 396884 358860 396886
rect 358924 396884 358971 396888
rect 362902 396884 362908 396948
rect 362972 396946 362978 396948
rect 363045 396946 363111 396949
rect 375373 396946 375439 396949
rect 362972 396944 363111 396946
rect 362972 396888 363050 396944
rect 363106 396888 363111 396944
rect 362972 396886 363111 396888
rect 362972 396884 362978 396886
rect 358905 396883 358971 396884
rect 363045 396883 363111 396886
rect 364290 396944 375439 396946
rect 364290 396888 375378 396944
rect 375434 396888 375439 396944
rect 364290 396886 375439 396888
rect 270033 396810 270099 396813
rect 352373 396810 352439 396813
rect 270033 396808 352439 396810
rect 270033 396752 270038 396808
rect 270094 396752 352378 396808
rect 352434 396752 352439 396808
rect 270033 396750 352439 396752
rect 270033 396747 270099 396750
rect 352373 396747 352439 396750
rect 353477 396810 353543 396813
rect 353477 396808 355610 396810
rect 353477 396752 353482 396808
rect 353538 396752 355610 396808
rect 353477 396750 355610 396752
rect 353477 396747 353543 396750
rect 270217 396674 270283 396677
rect 355550 396674 355610 396750
rect 356646 396748 356652 396812
rect 356716 396810 356722 396812
rect 364290 396810 364350 396886
rect 375373 396883 375439 396886
rect 356716 396750 364350 396810
rect 378041 396810 378107 396813
rect 378174 396810 378180 396812
rect 378041 396808 378180 396810
rect 378041 396752 378046 396808
rect 378102 396752 378180 396808
rect 378041 396750 378180 396752
rect 356716 396748 356722 396750
rect 378041 396747 378107 396750
rect 378174 396748 378180 396750
rect 378244 396748 378250 396812
rect 357382 396674 357388 396676
rect 270217 396672 355426 396674
rect 270217 396616 270222 396672
rect 270278 396616 355426 396672
rect 270217 396614 355426 396616
rect 355550 396614 357388 396674
rect 270217 396611 270283 396614
rect 340321 396538 340387 396541
rect 355174 396538 355180 396540
rect 340321 396536 355180 396538
rect 340321 396480 340326 396536
rect 340382 396480 355180 396536
rect 340321 396478 355180 396480
rect 340321 396475 340387 396478
rect 355174 396476 355180 396478
rect 355244 396476 355250 396540
rect 355366 396538 355426 396614
rect 357382 396612 357388 396614
rect 357452 396612 357458 396676
rect 358302 396612 358308 396676
rect 358372 396674 358378 396676
rect 362033 396674 362099 396677
rect 358372 396672 362099 396674
rect 358372 396616 362038 396672
rect 362094 396616 362099 396672
rect 358372 396614 362099 396616
rect 358372 396612 358378 396614
rect 362033 396611 362099 396614
rect 378174 396612 378180 396676
rect 378244 396674 378250 396676
rect 379329 396674 379395 396677
rect 378244 396672 379395 396674
rect 378244 396616 379334 396672
rect 379390 396616 379395 396672
rect 378244 396614 379395 396616
rect 378244 396612 378250 396614
rect 379329 396611 379395 396614
rect 379697 396674 379763 396677
rect 379830 396674 379836 396676
rect 379697 396672 379836 396674
rect 379697 396616 379702 396672
rect 379758 396616 379836 396672
rect 379697 396614 379836 396616
rect 379697 396611 379763 396614
rect 379830 396612 379836 396614
rect 379900 396612 379906 396676
rect 360285 396538 360351 396541
rect 355366 396536 360351 396538
rect 355366 396480 360290 396536
rect 360346 396480 360351 396536
rect 355366 396478 360351 396480
rect 360285 396475 360351 396478
rect 363454 396476 363460 396540
rect 363524 396538 363530 396540
rect 371049 396538 371115 396541
rect 363524 396536 371115 396538
rect 363524 396480 371054 396536
rect 371110 396480 371115 396536
rect 363524 396478 371115 396480
rect 363524 396476 363530 396478
rect 371049 396475 371115 396478
rect 377622 396476 377628 396540
rect 377692 396538 377698 396540
rect 381169 396538 381235 396541
rect 377692 396536 381235 396538
rect 377692 396480 381174 396536
rect 381230 396480 381235 396536
rect 377692 396478 381235 396480
rect 377692 396476 377698 396478
rect 381169 396475 381235 396478
rect 352373 396402 352439 396405
rect 359917 396402 359983 396405
rect 352373 396400 359983 396402
rect 352373 396344 352378 396400
rect 352434 396344 359922 396400
rect 359978 396344 359983 396400
rect 352373 396342 359983 396344
rect 352373 396339 352439 396342
rect 359917 396339 359983 396342
rect 361757 396402 361823 396405
rect 361757 396400 361866 396402
rect 361757 396344 361762 396400
rect 361818 396344 361866 396400
rect 361757 396339 361866 396344
rect 339861 396266 339927 396269
rect 354254 396266 354260 396268
rect 339861 396264 354260 396266
rect 339861 396208 339866 396264
rect 339922 396208 354260 396264
rect 339861 396206 354260 396208
rect 339861 396203 339927 396206
rect 354254 396204 354260 396206
rect 354324 396204 354330 396268
rect 361806 396130 361866 396339
rect 361941 396130 362007 396133
rect 361806 396128 362007 396130
rect 361806 396072 361946 396128
rect 362002 396072 362007 396128
rect 361806 396070 362007 396072
rect 361941 396067 362007 396070
rect 331949 395994 332015 395997
rect 350901 395994 350967 395997
rect 331949 395992 350967 395994
rect 331949 395936 331954 395992
rect 332010 395936 350906 395992
rect 350962 395936 350967 395992
rect 331949 395934 350967 395936
rect 331949 395931 332015 395934
rect 350901 395931 350967 395934
rect 354673 395994 354739 395997
rect 354806 395994 354812 395996
rect 354673 395992 354812 395994
rect 354673 395936 354678 395992
rect 354734 395936 354812 395992
rect 354673 395934 354812 395936
rect 354673 395931 354739 395934
rect 354806 395932 354812 395934
rect 354876 395932 354882 395996
rect 334801 395858 334867 395861
rect 367645 395858 367711 395861
rect 334801 395856 367711 395858
rect 334801 395800 334806 395856
rect 334862 395800 367650 395856
rect 367706 395800 367711 395856
rect 334801 395798 367711 395800
rect 334801 395795 334867 395798
rect 367645 395795 367711 395798
rect 341333 395722 341399 395725
rect 380249 395722 380315 395725
rect 341333 395720 380315 395722
rect 341333 395664 341338 395720
rect 341394 395664 380254 395720
rect 380310 395664 380315 395720
rect 341333 395662 380315 395664
rect 341333 395659 341399 395662
rect 380249 395659 380315 395662
rect 272885 395586 272951 395589
rect 342294 395586 342300 395588
rect 272885 395584 342300 395586
rect 272885 395528 272890 395584
rect 272946 395528 342300 395584
rect 272885 395526 342300 395528
rect 272885 395523 272951 395526
rect 342294 395524 342300 395526
rect 342364 395524 342370 395588
rect 368606 395524 368612 395588
rect 368676 395586 368682 395588
rect 368841 395586 368907 395589
rect 368676 395584 368907 395586
rect 368676 395528 368846 395584
rect 368902 395528 368907 395584
rect 368676 395526 368907 395528
rect 368676 395524 368682 395526
rect 368841 395523 368907 395526
rect 271781 395450 271847 395453
rect 352281 395450 352347 395453
rect 271781 395448 352347 395450
rect 271781 395392 271786 395448
rect 271842 395392 352286 395448
rect 352342 395392 352347 395448
rect 271781 395390 352347 395392
rect 271781 395387 271847 395390
rect 352281 395387 352347 395390
rect 373441 395450 373507 395453
rect 373758 395450 373764 395452
rect 373441 395448 373764 395450
rect 373441 395392 373446 395448
rect 373502 395392 373764 395448
rect 373441 395390 373764 395392
rect 373441 395387 373507 395390
rect 373758 395388 373764 395390
rect 373828 395388 373834 395452
rect 374126 395388 374132 395452
rect 374196 395450 374202 395452
rect 375189 395450 375255 395453
rect 374196 395448 375255 395450
rect 374196 395392 375194 395448
rect 375250 395392 375255 395448
rect 374196 395390 375255 395392
rect 374196 395388 374202 395390
rect 375189 395387 375255 395390
rect 271229 395314 271295 395317
rect 354622 395314 354628 395316
rect 271229 395312 354628 395314
rect 271229 395256 271234 395312
rect 271290 395256 354628 395312
rect 271229 395254 354628 395256
rect 271229 395251 271295 395254
rect 354622 395252 354628 395254
rect 354692 395252 354698 395316
rect 356830 395252 356836 395316
rect 356900 395314 356906 395316
rect 376937 395314 377003 395317
rect 356900 395312 377003 395314
rect 356900 395256 376942 395312
rect 376998 395256 377003 395312
rect 356900 395254 377003 395256
rect 356900 395252 356906 395254
rect 376937 395251 377003 395254
rect 379646 395252 379652 395316
rect 379716 395314 379722 395316
rect 380525 395314 380591 395317
rect 379716 395312 380591 395314
rect 379716 395256 380530 395312
rect 380586 395256 380591 395312
rect 379716 395254 380591 395256
rect 379716 395252 379722 395254
rect 380525 395251 380591 395254
rect 368381 395180 368447 395181
rect 368381 395176 368428 395180
rect 368492 395178 368498 395180
rect 378317 395178 378383 395181
rect 379094 395178 379100 395180
rect 368381 395120 368386 395176
rect 368381 395116 368428 395120
rect 368492 395118 368538 395178
rect 378317 395176 379100 395178
rect 378317 395120 378322 395176
rect 378378 395120 379100 395176
rect 378317 395118 379100 395120
rect 368492 395116 368498 395118
rect 368381 395115 368447 395116
rect 378317 395115 378383 395118
rect 379094 395116 379100 395118
rect 379164 395116 379170 395180
rect 338849 394770 338915 394773
rect 345422 394770 345428 394772
rect 338849 394768 345428 394770
rect 338849 394712 338854 394768
rect 338910 394712 345428 394768
rect 338849 394710 345428 394712
rect 338849 394707 338915 394710
rect 345422 394708 345428 394710
rect 345492 394708 345498 394772
rect 297214 394572 297220 394636
rect 297284 394634 297290 394636
rect 356421 394634 356487 394637
rect 297284 394632 356487 394634
rect 297284 394576 356426 394632
rect 356482 394576 356487 394632
rect 297284 394574 356487 394576
rect 297284 394572 297290 394574
rect 356421 394571 356487 394574
rect 368933 394634 368999 394637
rect 372286 394634 372292 394636
rect 368933 394632 372292 394634
rect 368933 394576 368938 394632
rect 368994 394576 372292 394632
rect 368933 394574 372292 394576
rect 368933 394571 368999 394574
rect 372286 394572 372292 394574
rect 372356 394572 372362 394636
rect 297950 394436 297956 394500
rect 298020 394498 298026 394500
rect 357566 394498 357572 394500
rect 298020 394438 357572 394498
rect 298020 394436 298026 394438
rect 357566 394436 357572 394438
rect 357636 394436 357642 394500
rect 296478 394300 296484 394364
rect 296548 394362 296554 394364
rect 355593 394362 355659 394365
rect 296548 394360 355659 394362
rect 296548 394304 355598 394360
rect 355654 394304 355659 394360
rect 296548 394302 355659 394304
rect 296548 394300 296554 394302
rect 355593 394299 355659 394302
rect 321318 394164 321324 394228
rect 321388 394226 321394 394228
rect 381537 394226 381603 394229
rect 321388 394224 381603 394226
rect 321388 394168 381542 394224
rect 381598 394168 381603 394224
rect 321388 394166 381603 394168
rect 321388 394164 321394 394166
rect 381537 394163 381603 394166
rect 270401 394090 270467 394093
rect 359917 394090 359983 394093
rect 270401 394088 359983 394090
rect 270401 394032 270406 394088
rect 270462 394032 359922 394088
rect 359978 394032 359983 394088
rect 270401 394030 359983 394032
rect 270401 394027 270467 394030
rect 359917 394027 359983 394030
rect 273713 393954 273779 393957
rect 366633 393954 366699 393957
rect 273713 393952 366699 393954
rect 273713 393896 273718 393952
rect 273774 393896 366638 393952
rect 366694 393896 366699 393952
rect 273713 393894 366699 393896
rect 273713 393891 273779 393894
rect 366633 393891 366699 393894
rect 372654 393892 372660 393956
rect 372724 393954 372730 393956
rect 373533 393954 373599 393957
rect 372724 393952 373599 393954
rect 372724 393896 373538 393952
rect 373594 393896 373599 393952
rect 372724 393894 373599 393896
rect 372724 393892 372730 393894
rect 373533 393891 373599 393894
rect 355593 393818 355659 393821
rect 374085 393818 374151 393821
rect 355593 393816 374151 393818
rect 355593 393760 355598 393816
rect 355654 393760 374090 393816
rect 374146 393760 374151 393816
rect 355593 393758 374151 393760
rect 355593 393755 355659 393758
rect 374085 393755 374151 393758
rect 343541 393546 343607 393549
rect 350022 393546 350028 393548
rect 343541 393544 350028 393546
rect 343541 393488 343546 393544
rect 343602 393488 350028 393544
rect 343541 393486 350028 393488
rect 343541 393483 343607 393486
rect 350022 393484 350028 393486
rect 350092 393484 350098 393548
rect 357934 393484 357940 393548
rect 358004 393546 358010 393548
rect 369577 393546 369643 393549
rect 358004 393544 369643 393546
rect 358004 393488 369582 393544
rect 369638 393488 369643 393544
rect 358004 393486 369643 393488
rect 358004 393484 358010 393486
rect 369577 393483 369643 393486
rect 378133 393546 378199 393549
rect 378358 393546 378364 393548
rect 378133 393544 378364 393546
rect 378133 393488 378138 393544
rect 378194 393488 378364 393544
rect 378133 393486 378364 393488
rect 378133 393483 378199 393486
rect 378358 393484 378364 393486
rect 378428 393484 378434 393548
rect 344093 393410 344159 393413
rect 344686 393410 344692 393412
rect 344093 393408 344692 393410
rect 344093 393352 344098 393408
rect 344154 393352 344692 393408
rect 344093 393350 344692 393352
rect 344093 393347 344159 393350
rect 344686 393348 344692 393350
rect 344756 393348 344762 393412
rect 347814 393348 347820 393412
rect 347884 393410 347890 393412
rect 348509 393410 348575 393413
rect 349337 393412 349403 393413
rect 349286 393410 349292 393412
rect 347884 393408 348575 393410
rect 347884 393352 348514 393408
rect 348570 393352 348575 393408
rect 347884 393350 348575 393352
rect 349246 393350 349292 393410
rect 349356 393408 349403 393412
rect 349398 393352 349403 393408
rect 347884 393348 347890 393350
rect 348509 393347 348575 393350
rect 349286 393348 349292 393350
rect 349356 393348 349403 393352
rect 362534 393348 362540 393412
rect 362604 393410 362610 393412
rect 369710 393410 369716 393412
rect 362604 393350 369716 393410
rect 362604 393348 362610 393350
rect 369710 393348 369716 393350
rect 369780 393348 369786 393412
rect 349337 393347 349403 393348
rect 299238 393212 299244 393276
rect 299308 393274 299314 393276
rect 357893 393274 357959 393277
rect 299308 393272 357959 393274
rect 299308 393216 357898 393272
rect 357954 393216 357959 393272
rect 299308 393214 357959 393216
rect 299308 393212 299314 393214
rect 357893 393211 357959 393214
rect 360469 393274 360535 393277
rect 360878 393274 360884 393276
rect 360469 393272 360884 393274
rect 360469 393216 360474 393272
rect 360530 393216 360884 393272
rect 360469 393214 360884 393216
rect 360469 393211 360535 393214
rect 360878 393212 360884 393214
rect 360948 393212 360954 393276
rect 364926 393212 364932 393276
rect 364996 393274 365002 393276
rect 367277 393274 367343 393277
rect 364996 393272 367343 393274
rect 364996 393216 367282 393272
rect 367338 393216 367343 393272
rect 364996 393214 367343 393216
rect 364996 393212 365002 393214
rect 367277 393211 367343 393214
rect 367870 393212 367876 393276
rect 367940 393274 367946 393276
rect 368013 393274 368079 393277
rect 367940 393272 368079 393274
rect 367940 393216 368018 393272
rect 368074 393216 368079 393272
rect 367940 393214 368079 393216
rect 367940 393212 367946 393214
rect 368013 393211 368079 393214
rect 306230 393076 306236 393140
rect 306300 393138 306306 393140
rect 364190 393138 364196 393140
rect 306300 393078 364196 393138
rect 306300 393076 306306 393078
rect 364190 393076 364196 393078
rect 364260 393076 364266 393140
rect 365897 393138 365963 393141
rect 366766 393138 366772 393140
rect 365897 393136 366772 393138
rect 365897 393080 365902 393136
rect 365958 393080 366772 393136
rect 365897 393078 366772 393080
rect 365897 393075 365963 393078
rect 366766 393076 366772 393078
rect 366836 393076 366842 393140
rect 367686 393076 367692 393140
rect 367756 393138 367762 393140
rect 370129 393138 370195 393141
rect 367756 393136 370195 393138
rect 367756 393080 370134 393136
rect 370190 393080 370195 393136
rect 367756 393078 370195 393080
rect 367756 393076 367762 393078
rect 370129 393075 370195 393078
rect 304758 392940 304764 393004
rect 304828 393002 304834 393004
rect 361297 393002 361363 393005
rect 304828 393000 361363 393002
rect 304828 392944 361302 393000
rect 361358 392944 361363 393000
rect 304828 392942 361363 392944
rect 304828 392940 304834 392942
rect 361297 392939 361363 392942
rect 366214 392940 366220 393004
rect 366284 393002 366290 393004
rect 367645 393002 367711 393005
rect 366284 393000 367711 393002
rect 366284 392944 367650 393000
rect 367706 392944 367711 393000
rect 366284 392942 367711 392944
rect 366284 392940 366290 392942
rect 367645 392939 367711 392942
rect 300710 392804 300716 392868
rect 300780 392866 300786 392868
rect 360561 392866 360627 392869
rect 300780 392864 360627 392866
rect 300780 392808 360566 392864
rect 360622 392808 360627 392864
rect 300780 392806 360627 392808
rect 300780 392804 300786 392806
rect 360561 392803 360627 392806
rect 367277 392866 367343 392869
rect 368054 392866 368060 392868
rect 367277 392864 368060 392866
rect 367277 392808 367282 392864
rect 367338 392808 368060 392864
rect 367277 392806 368060 392808
rect 367277 392803 367343 392806
rect 368054 392804 368060 392806
rect 368124 392804 368130 392868
rect 304574 392668 304580 392732
rect 304644 392730 304650 392732
rect 362861 392730 362927 392733
rect 304644 392728 362927 392730
rect 304644 392672 362866 392728
rect 362922 392672 362927 392728
rect 304644 392670 362927 392672
rect 304644 392668 304650 392670
rect 362861 392667 362927 392670
rect 293166 392532 293172 392596
rect 293236 392594 293242 392596
rect 352230 392594 352236 392596
rect 293236 392534 352236 392594
rect 293236 392532 293242 392534
rect 352230 392532 352236 392534
rect 352300 392532 352306 392596
rect 358077 392594 358143 392597
rect 358670 392594 358676 392596
rect 358077 392592 358676 392594
rect 358077 392536 358082 392592
rect 358138 392536 358676 392592
rect 358077 392534 358676 392536
rect 358077 392531 358143 392534
rect 358670 392532 358676 392534
rect 358740 392532 358746 392596
rect 303470 392396 303476 392460
rect 303540 392458 303546 392460
rect 362769 392458 362835 392461
rect 303540 392456 362835 392458
rect 303540 392400 362774 392456
rect 362830 392400 362835 392456
rect 303540 392398 362835 392400
rect 303540 392396 303546 392398
rect 362769 392395 362835 392398
rect 282913 392052 282979 392053
rect 282862 392050 282868 392052
rect 282822 391990 282868 392050
rect 282932 392048 282979 392052
rect 282974 391992 282979 392048
rect 282862 391988 282868 391990
rect 282932 391988 282979 391992
rect 341006 391988 341012 392052
rect 341076 392050 341082 392052
rect 341793 392050 341859 392053
rect 341076 392048 341859 392050
rect 341076 391992 341798 392048
rect 341854 391992 341859 392048
rect 341076 391990 341859 391992
rect 341076 391988 341082 391990
rect 282913 391987 282979 391988
rect 341793 391987 341859 391990
rect 311750 391716 311756 391780
rect 311820 391778 311826 391780
rect 371182 391778 371188 391780
rect 311820 391718 371188 391778
rect 311820 391716 311826 391718
rect 371182 391716 371188 391718
rect 371252 391716 371258 391780
rect 295006 391580 295012 391644
rect 295076 391642 295082 391644
rect 353702 391642 353708 391644
rect 295076 391582 353708 391642
rect 295076 391580 295082 391582
rect 353702 391580 353708 391582
rect 353772 391580 353778 391644
rect 583520 391628 584960 391868
rect 269021 391506 269087 391509
rect 340965 391506 341031 391509
rect 269021 391504 341031 391506
rect 269021 391448 269026 391504
rect 269082 391448 340970 391504
rect 341026 391448 341031 391504
rect 269021 391446 341031 391448
rect 269021 391443 269087 391446
rect 340965 391443 341031 391446
rect 263501 391370 263567 391373
rect 344737 391370 344803 391373
rect 263501 391368 344803 391370
rect 263501 391312 263506 391368
rect 263562 391312 344742 391368
rect 344798 391312 344803 391368
rect 263501 391310 344803 391312
rect 263501 391307 263567 391310
rect 344737 391307 344803 391310
rect 262029 391234 262095 391237
rect 346301 391234 346367 391237
rect 262029 391232 346367 391234
rect 262029 391176 262034 391232
rect 262090 391176 346306 391232
rect 346362 391176 346367 391232
rect 262029 391174 346367 391176
rect 262029 391171 262095 391174
rect 346301 391171 346367 391174
rect 295190 391036 295196 391100
rect 295260 391098 295266 391100
rect 353017 391098 353083 391101
rect 295260 391096 353083 391098
rect 295260 391040 353022 391096
rect 353078 391040 353083 391096
rect 295260 391038 353083 391040
rect 295260 391036 295266 391038
rect 353017 391035 353083 391038
rect 314142 390900 314148 390964
rect 314212 390962 314218 390964
rect 373901 390962 373967 390965
rect 314212 390960 373967 390962
rect 314212 390904 373906 390960
rect 373962 390904 373967 390960
rect 314212 390902 373967 390904
rect 314212 390900 314218 390902
rect 373901 390899 373967 390902
rect 294638 390492 294644 390556
rect 294708 390554 294714 390556
rect 341149 390554 341215 390557
rect 294708 390552 341215 390554
rect 294708 390496 341154 390552
rect 341210 390496 341215 390552
rect 294708 390494 341215 390496
rect 294708 390492 294714 390494
rect 341149 390491 341215 390494
rect 317270 390356 317276 390420
rect 317340 390418 317346 390420
rect 377581 390418 377647 390421
rect 317340 390416 377647 390418
rect 317340 390360 377586 390416
rect 377642 390360 377647 390416
rect 317340 390358 377647 390360
rect 317340 390356 317346 390358
rect 377581 390355 377647 390358
rect 278037 390282 278103 390285
rect 351085 390282 351151 390285
rect 278037 390280 351151 390282
rect 278037 390224 278042 390280
rect 278098 390224 351090 390280
rect 351146 390224 351151 390280
rect 278037 390222 351151 390224
rect 278037 390219 278103 390222
rect 351085 390219 351151 390222
rect 268653 390146 268719 390149
rect 350165 390146 350231 390149
rect 268653 390144 350231 390146
rect 268653 390088 268658 390144
rect 268714 390088 350170 390144
rect 350226 390088 350231 390144
rect 268653 390086 350231 390088
rect 268653 390083 268719 390086
rect 350165 390083 350231 390086
rect 266169 390010 266235 390013
rect 345841 390010 345907 390013
rect 266169 390008 345907 390010
rect 266169 389952 266174 390008
rect 266230 389952 345846 390008
rect 345902 389952 345907 390008
rect 266169 389950 345907 389952
rect 266169 389947 266235 389950
rect 345841 389947 345907 389950
rect 260649 389874 260715 389877
rect 344553 389874 344619 389877
rect 260649 389872 344619 389874
rect 260649 389816 260654 389872
rect 260710 389816 344558 389872
rect 344614 389816 344619 389872
rect 260649 389814 344619 389816
rect 260649 389811 260715 389814
rect 344553 389811 344619 389814
rect 345054 389812 345060 389876
rect 345124 389874 345130 389876
rect 345933 389874 345999 389877
rect 345124 389872 345999 389874
rect 345124 389816 345938 389872
rect 345994 389816 345999 389872
rect 345124 389814 345999 389816
rect 345124 389812 345130 389814
rect 345933 389811 345999 389814
rect 316718 389676 316724 389740
rect 316788 389738 316794 389740
rect 372429 389738 372495 389741
rect 316788 389736 372495 389738
rect 316788 389680 372434 389736
rect 372490 389680 372495 389736
rect 316788 389678 372495 389680
rect 316788 389676 316794 389678
rect 372429 389675 372495 389678
rect 378133 389330 378199 389333
rect 378542 389330 378548 389332
rect 378133 389328 378548 389330
rect 378133 389272 378138 389328
rect 378194 389272 378548 389328
rect 378133 389270 378548 389272
rect 378133 389267 378199 389270
rect 378542 389268 378548 389270
rect 378612 389268 378618 389332
rect 373901 389196 373967 389197
rect 373901 389194 373948 389196
rect 373856 389192 373948 389194
rect 373856 389136 373906 389192
rect 373856 389134 373948 389136
rect 373901 389132 373948 389134
rect 374012 389132 374018 389196
rect 373901 389131 373967 389132
rect 291694 388996 291700 389060
rect 291764 389058 291770 389060
rect 345013 389058 345079 389061
rect 291764 389056 345079 389058
rect 291764 389000 345018 389056
rect 345074 389000 345079 389056
rect 291764 388998 345079 389000
rect 291764 388996 291770 388998
rect 345013 388995 345079 388998
rect 288014 388860 288020 388924
rect 288084 388922 288090 388924
rect 347865 388922 347931 388925
rect 288084 388920 347931 388922
rect 288084 388864 347870 388920
rect 347926 388864 347931 388920
rect 288084 388862 347931 388864
rect 288084 388860 288090 388862
rect 347865 388859 347931 388862
rect 287462 388724 287468 388788
rect 287532 388786 287538 388788
rect 348366 388786 348372 388788
rect 287532 388726 348372 388786
rect 287532 388724 287538 388726
rect 348366 388724 348372 388726
rect 348436 388724 348442 388788
rect 289486 388588 289492 388652
rect 289556 388650 289562 388652
rect 348550 388650 348556 388652
rect 289556 388590 348556 388650
rect 289556 388588 289562 388590
rect 348550 388588 348556 388590
rect 348620 388588 348626 388652
rect 268837 388514 268903 388517
rect 344870 388514 344876 388516
rect 268837 388512 344876 388514
rect 268837 388456 268842 388512
rect 268898 388456 344876 388512
rect 268837 388454 344876 388456
rect 268837 388451 268903 388454
rect 344870 388452 344876 388454
rect 344940 388452 344946 388516
rect 347497 388514 347563 388517
rect 383694 388514 383700 388516
rect 347497 388512 383700 388514
rect 347497 388456 347502 388512
rect 347558 388456 383700 388512
rect 347497 388454 383700 388456
rect 347497 388451 347563 388454
rect 383694 388452 383700 388454
rect 383764 388452 383770 388516
rect 260465 388378 260531 388381
rect 345238 388378 345244 388380
rect 260465 388376 345244 388378
rect 260465 388320 260470 388376
rect 260526 388320 345244 388376
rect 260465 388318 345244 388320
rect 260465 388315 260531 388318
rect 345238 388316 345244 388318
rect 345308 388316 345314 388380
rect 345565 388378 345631 388381
rect 384982 388378 384988 388380
rect 345565 388376 384988 388378
rect 345565 388320 345570 388376
rect 345626 388320 384988 388376
rect 345565 388318 384988 388320
rect 345565 388315 345631 388318
rect 384982 388316 384988 388318
rect 385052 388316 385058 388380
rect 286726 388180 286732 388244
rect 286796 388242 286802 388244
rect 346209 388242 346275 388245
rect 286796 388240 346275 388242
rect 286796 388184 346214 388240
rect 346270 388184 346275 388240
rect 286796 388182 346275 388184
rect 286796 388180 286802 388182
rect 346209 388179 346275 388182
rect 307518 387636 307524 387700
rect 307588 387698 307594 387700
rect 366582 387698 366588 387700
rect 307588 387638 366588 387698
rect 307588 387636 307594 387638
rect 366582 387636 366588 387638
rect 366652 387636 366658 387700
rect 287830 387500 287836 387564
rect 287900 387562 287906 387564
rect 346393 387562 346459 387565
rect 287900 387560 346459 387562
rect 287900 387504 346398 387560
rect 346454 387504 346459 387560
rect 287900 387502 346459 387504
rect 287900 387500 287906 387502
rect 346393 387499 346459 387502
rect 297582 387364 297588 387428
rect 297652 387426 297658 387428
rect 357617 387426 357683 387429
rect 297652 387424 357683 387426
rect 297652 387368 357622 387424
rect 357678 387368 357683 387424
rect 297652 387366 357683 387368
rect 297652 387364 297658 387366
rect 357617 387363 357683 387366
rect 273897 387290 273963 387293
rect 344185 387290 344251 387293
rect 273897 387288 344251 387290
rect 273897 387232 273902 387288
rect 273958 387232 344190 387288
rect 344246 387232 344251 387288
rect 273897 387230 344251 387232
rect 273897 387227 273963 387230
rect 344185 387227 344251 387230
rect 281390 387092 281396 387156
rect 281460 387154 281466 387156
rect 357014 387154 357020 387156
rect 281460 387094 357020 387154
rect 281460 387092 281466 387094
rect 357014 387092 357020 387094
rect 357084 387092 357090 387156
rect 260557 387018 260623 387021
rect 347262 387018 347268 387020
rect 260557 387016 347268 387018
rect 260557 386960 260562 387016
rect 260618 386960 347268 387016
rect 260557 386958 347268 386960
rect 260557 386955 260623 386958
rect 347262 386956 347268 386958
rect 347332 386956 347338 387020
rect 301998 385868 302004 385932
rect 302068 385930 302074 385932
rect 360469 385930 360535 385933
rect 302068 385928 360535 385930
rect 302068 385872 360474 385928
rect 360530 385872 360535 385928
rect 302068 385870 360535 385872
rect 302068 385868 302074 385870
rect 360469 385867 360535 385870
rect 317689 385794 317755 385797
rect 376886 385794 376892 385796
rect 317689 385792 376892 385794
rect 317689 385736 317694 385792
rect 317750 385736 376892 385792
rect 317689 385734 376892 385736
rect 317689 385731 317755 385734
rect 376886 385732 376892 385734
rect 376956 385732 376962 385796
rect 268745 385658 268811 385661
rect 360326 385658 360332 385660
rect 268745 385656 360332 385658
rect 268745 385600 268750 385656
rect 268806 385600 360332 385656
rect 268745 385598 360332 385600
rect 268745 385595 268811 385598
rect 360326 385596 360332 385598
rect 360396 385596 360402 385660
rect -960 384284 480 384524
rect 298870 384372 298876 384436
rect 298940 384434 298946 384436
rect 357525 384434 357591 384437
rect 298940 384432 357591 384434
rect 298940 384376 357530 384432
rect 357586 384376 357591 384432
rect 298940 384374 357591 384376
rect 298940 384372 298946 384374
rect 357525 384371 357591 384374
rect 303613 384298 303679 384301
rect 363270 384298 363276 384300
rect 303613 384296 363276 384298
rect 303613 384240 303618 384296
rect 303674 384240 363276 384296
rect 303613 384238 363276 384240
rect 303613 384235 303679 384238
rect 363270 384236 363276 384238
rect 363340 384236 363346 384300
rect 373942 383828 373948 383892
rect 374012 383828 374018 383892
rect 373950 383757 374010 383828
rect 373901 383754 374010 383757
rect 373856 383752 374010 383754
rect 373856 383696 373906 383752
rect 373962 383696 374010 383752
rect 373856 383694 374010 383696
rect 373901 383691 373967 383694
rect 373901 383618 373967 383621
rect 373856 383616 374010 383618
rect 373856 383560 373906 383616
rect 373962 383560 374010 383616
rect 373856 383558 374010 383560
rect 373901 383555 374010 383558
rect 373950 383484 374010 383555
rect 373942 383420 373948 383484
rect 374012 383420 374018 383484
rect 349981 382122 350047 382125
rect 366398 382122 366404 382124
rect 349981 382120 366404 382122
rect 349981 382064 349986 382120
rect 350042 382064 366404 382120
rect 349981 382062 366404 382064
rect 349981 382059 350047 382062
rect 366398 382060 366404 382062
rect 366468 382060 366474 382124
rect 344369 381986 344435 381989
rect 364374 381986 364380 381988
rect 344369 381984 364380 381986
rect 344369 381928 344374 381984
rect 344430 381928 364380 381984
rect 344369 381926 364380 381928
rect 344369 381923 344435 381926
rect 364374 381924 364380 381926
rect 364444 381924 364450 381988
rect 351545 381850 351611 381853
rect 371734 381850 371740 381852
rect 351545 381848 371740 381850
rect 351545 381792 351550 381848
rect 351606 381792 371740 381848
rect 351545 381790 371740 381792
rect 351545 381787 351611 381790
rect 371734 381788 371740 381790
rect 371804 381788 371810 381852
rect 286358 381652 286364 381716
rect 286428 381714 286434 381716
rect 343817 381714 343883 381717
rect 286428 381712 343883 381714
rect 286428 381656 343822 381712
rect 343878 381656 343883 381712
rect 286428 381654 343883 381656
rect 286428 381652 286434 381654
rect 343817 381651 343883 381654
rect 347221 381714 347287 381717
rect 368606 381714 368612 381716
rect 347221 381712 368612 381714
rect 347221 381656 347226 381712
rect 347282 381656 368612 381712
rect 347221 381654 368612 381656
rect 347221 381651 347287 381654
rect 368606 381652 368612 381654
rect 368676 381652 368682 381716
rect 292982 381516 292988 381580
rect 293052 381578 293058 381580
rect 353569 381578 353635 381581
rect 293052 381576 353635 381578
rect 293052 381520 353574 381576
rect 353630 381520 353635 381576
rect 293052 381518 353635 381520
rect 293052 381516 293058 381518
rect 353569 381515 353635 381518
rect 291878 379340 291884 379404
rect 291948 379402 291954 379404
rect 350901 379402 350967 379405
rect 291948 379400 350967 379402
rect 291948 379344 350906 379400
rect 350962 379344 350967 379400
rect 291948 379342 350967 379344
rect 291948 379340 291954 379342
rect 350901 379339 350967 379342
rect 290958 379204 290964 379268
rect 291028 379266 291034 379268
rect 349521 379266 349587 379269
rect 291028 379264 349587 379266
rect 291028 379208 349526 379264
rect 349582 379208 349587 379264
rect 291028 379206 349587 379208
rect 291028 379204 291034 379206
rect 349521 379203 349587 379206
rect 291326 379068 291332 379132
rect 291396 379130 291402 379132
rect 350993 379130 351059 379133
rect 291396 379128 351059 379130
rect 291396 379072 350998 379128
rect 351054 379072 351059 379128
rect 291396 379070 351059 379072
rect 291396 379068 291402 379070
rect 350993 379067 351059 379070
rect 292246 378932 292252 378996
rect 292316 378994 292322 378996
rect 352281 378994 352347 378997
rect 292316 378992 352347 378994
rect 292316 378936 352286 378992
rect 352342 378936 352347 378992
rect 292316 378934 352347 378936
rect 292316 378932 292322 378934
rect 352281 378931 352347 378934
rect 290774 378796 290780 378860
rect 290844 378858 290850 378860
rect 350809 378858 350875 378861
rect 290844 378856 350875 378858
rect 290844 378800 350814 378856
rect 350870 378800 350875 378856
rect 290844 378798 350875 378800
rect 290844 378796 290850 378798
rect 350809 378795 350875 378798
rect 288750 378660 288756 378724
rect 288820 378722 288826 378724
rect 349429 378722 349495 378725
rect 288820 378720 349495 378722
rect 288820 378664 349434 378720
rect 349490 378664 349495 378720
rect 288820 378662 349495 378664
rect 288820 378660 288826 378662
rect 349429 378659 349495 378662
rect 289302 378524 289308 378588
rect 289372 378586 289378 378588
rect 344921 378586 344987 378589
rect 289372 378584 344987 378586
rect 289372 378528 344926 378584
rect 344982 378528 344987 378584
rect 289372 378526 344987 378528
rect 289372 378524 289378 378526
rect 344921 378523 344987 378526
rect 580257 378450 580323 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 583520 378300 584960 378390
rect 350073 378042 350139 378045
rect 354806 378042 354812 378044
rect 350073 378040 354812 378042
rect 350073 377984 350078 378040
rect 350134 377984 354812 378040
rect 350073 377982 354812 377984
rect 350073 377979 350139 377982
rect 354806 377980 354812 377982
rect 354876 377980 354882 378044
rect 348877 377906 348943 377909
rect 353334 377906 353340 377908
rect 348877 377904 353340 377906
rect 348877 377848 348882 377904
rect 348938 377848 353340 377904
rect 348877 377846 353340 377848
rect 348877 377843 348943 377846
rect 353334 377844 353340 377846
rect 353404 377844 353410 377908
rect 308990 377436 308996 377500
rect 309060 377498 309066 377500
rect 367277 377498 367343 377501
rect 309060 377496 367343 377498
rect 309060 377440 367282 377496
rect 367338 377440 367343 377496
rect 309060 377438 367343 377440
rect 309060 377436 309066 377438
rect 367277 377435 367343 377438
rect 314694 377300 314700 377364
rect 314764 377362 314770 377364
rect 374729 377362 374795 377365
rect 314764 377360 374795 377362
rect 314764 377304 374734 377360
rect 374790 377304 374795 377360
rect 314764 377302 374795 377304
rect 314764 377300 314770 377302
rect 374729 377299 374795 377302
rect 285070 376756 285076 376820
rect 285140 376818 285146 376820
rect 289077 376818 289143 376821
rect 285140 376816 289143 376818
rect 285140 376760 289082 376816
rect 289138 376760 289143 376816
rect 285140 376758 289143 376760
rect 285140 376756 285146 376758
rect 289077 376755 289143 376758
rect 296294 375940 296300 376004
rect 296364 376002 296370 376004
rect 356329 376002 356395 376005
rect 296364 376000 356395 376002
rect 296364 375944 356334 376000
rect 356390 375944 356395 376000
rect 296364 375942 356395 375944
rect 296364 375940 296370 375942
rect 356329 375939 356395 375942
rect 279366 375396 279372 375460
rect 279436 375458 279442 375460
rect 309593 375458 309659 375461
rect 310053 375458 310119 375461
rect 279436 375456 310119 375458
rect 279436 375400 309598 375456
rect 309654 375400 310058 375456
rect 310114 375400 310119 375456
rect 279436 375398 310119 375400
rect 279436 375396 279442 375398
rect 309593 375395 309659 375398
rect 310053 375395 310119 375398
rect 292798 374716 292804 374780
rect 292868 374778 292874 374780
rect 347957 374778 348023 374781
rect 292868 374776 348023 374778
rect 292868 374720 347962 374776
rect 348018 374720 348023 374776
rect 292868 374718 348023 374720
rect 292868 374716 292874 374718
rect 347957 374715 348023 374718
rect 297398 374580 297404 374644
rect 297468 374642 297474 374644
rect 356237 374642 356303 374645
rect 297468 374640 356303 374642
rect 297468 374584 356242 374640
rect 356298 374584 356303 374640
rect 297468 374582 356303 374584
rect 297468 374580 297474 374582
rect 356237 374579 356303 374582
rect 287145 374506 287211 374509
rect 287697 374506 287763 374509
rect 287145 374504 287763 374506
rect 287145 374448 287150 374504
rect 287206 374448 287702 374504
rect 287758 374448 287763 374504
rect 287145 374446 287763 374448
rect 287145 374443 287211 374446
rect 287697 374443 287763 374446
rect 222101 374098 222167 374101
rect 287145 374098 287211 374101
rect 373901 374100 373967 374101
rect 373901 374098 373948 374100
rect 222101 374096 287211 374098
rect 222101 374040 222106 374096
rect 222162 374040 287150 374096
rect 287206 374040 287211 374096
rect 222101 374038 287211 374040
rect 373856 374096 373948 374098
rect 374012 374098 374018 374100
rect 373856 374040 373906 374096
rect 373856 374038 373948 374040
rect 222101 374035 222167 374038
rect 287145 374035 287211 374038
rect 373901 374036 373948 374038
rect 374012 374038 374094 374098
rect 374012 374036 374018 374038
rect 373901 374035 373967 374036
rect 280797 373962 280863 373965
rect 284109 373962 284175 373965
rect 373901 373962 373967 373965
rect 280797 373960 284175 373962
rect 280797 373904 280802 373960
rect 280858 373904 284114 373960
rect 284170 373904 284175 373960
rect 280797 373902 284175 373904
rect 373856 373960 374010 373962
rect 373856 373904 373906 373960
rect 373962 373904 374010 373960
rect 373856 373902 374010 373904
rect 280797 373899 280863 373902
rect 284109 373899 284175 373902
rect 373901 373899 374010 373902
rect 373950 373828 374010 373899
rect 373942 373764 373948 373828
rect 374012 373764 374018 373828
rect 220670 373356 220676 373420
rect 220740 373418 220746 373420
rect 278313 373418 278379 373421
rect 220740 373416 278379 373418
rect 220740 373360 278318 373416
rect 278374 373360 278379 373416
rect 220740 373358 278379 373360
rect 220740 373356 220746 373358
rect 278313 373355 278379 373358
rect 220445 373282 220511 373285
rect 280889 373282 280955 373285
rect 284201 373282 284267 373285
rect 220445 373280 284267 373282
rect 220445 373224 220450 373280
rect 220506 373224 280894 373280
rect 280950 373224 284206 373280
rect 284262 373224 284267 373280
rect 220445 373222 284267 373224
rect 220445 373219 220511 373222
rect 280889 373219 280955 373222
rect 284201 373219 284267 373222
rect 280470 372948 280476 373012
rect 280540 373010 280546 373012
rect 280797 373010 280863 373013
rect 280540 373008 280863 373010
rect 280540 372952 280802 373008
rect 280858 372952 280863 373008
rect 280540 372950 280863 372952
rect 280540 372948 280546 372950
rect 280797 372947 280863 372950
rect 279918 372676 279924 372740
rect 279988 372738 279994 372740
rect 286041 372738 286107 372741
rect 279988 372736 286107 372738
rect 279988 372680 286046 372736
rect 286102 372680 286107 372736
rect 279988 372678 286107 372680
rect 279988 372676 279994 372678
rect 286041 372675 286107 372678
rect 310513 372602 310579 372605
rect 311341 372602 311407 372605
rect 292530 372600 311407 372602
rect 292530 372544 310518 372600
rect 310574 372544 311346 372600
rect 311402 372544 311407 372600
rect 292530 372542 311407 372544
rect 280654 372268 280660 372332
rect 280724 372330 280730 372332
rect 292530 372330 292590 372542
rect 310513 372539 310579 372542
rect 311341 372539 311407 372542
rect 280724 372270 292590 372330
rect 280724 372268 280730 372270
rect 277894 372132 277900 372196
rect 277964 372194 277970 372196
rect 289721 372194 289787 372197
rect 277964 372192 289787 372194
rect 277964 372136 289726 372192
rect 289782 372136 289787 372192
rect 277964 372134 289787 372136
rect 277964 372132 277970 372134
rect 289721 372131 289787 372134
rect 276606 371996 276612 372060
rect 276676 372058 276682 372060
rect 280613 372058 280679 372061
rect 276676 372056 280679 372058
rect 276676 372000 280618 372056
rect 280674 372000 280679 372056
rect 276676 371998 280679 372000
rect 276676 371996 276682 371998
rect 280613 371995 280679 371998
rect 280061 371922 280127 371925
rect 287789 371922 287855 371925
rect 280061 371920 287855 371922
rect 280061 371864 280066 371920
rect 280122 371864 287794 371920
rect 287850 371864 287855 371920
rect 280061 371862 287855 371864
rect 280061 371859 280127 371862
rect 287789 371859 287855 371862
rect 314326 371860 314332 371924
rect 314396 371922 314402 371924
rect 372654 371922 372660 371924
rect 314396 371862 372660 371922
rect 314396 371860 314402 371862
rect 372654 371860 372660 371862
rect 372724 371860 372730 371924
rect 277761 371786 277827 371789
rect 278313 371786 278379 371789
rect 289997 371786 290063 371789
rect 310237 371786 310303 371789
rect 277761 371784 290063 371786
rect 277761 371728 277766 371784
rect 277822 371728 278318 371784
rect 278374 371728 290002 371784
rect 290058 371728 290063 371784
rect 277761 371726 290063 371728
rect 277761 371723 277827 371726
rect 278313 371723 278379 371726
rect 289997 371723 290063 371726
rect 292530 371784 310303 371786
rect 292530 371728 310242 371784
rect 310298 371728 310303 371784
rect 292530 371726 310303 371728
rect 284109 371650 284175 371653
rect 292530 371650 292590 371726
rect 310237 371723 310303 371726
rect 284109 371648 292590 371650
rect 284109 371592 284114 371648
rect 284170 371592 292590 371648
rect 284109 371590 292590 371592
rect 284109 371587 284175 371590
rect -960 371378 480 371468
rect 279550 371452 279556 371516
rect 279620 371514 279626 371516
rect 288249 371514 288315 371517
rect 279620 371512 288315 371514
rect 279620 371456 288254 371512
rect 288310 371456 288315 371512
rect 279620 371454 288315 371456
rect 279620 371452 279626 371454
rect 288249 371451 288315 371454
rect 307702 371452 307708 371516
rect 307772 371514 307778 371516
rect 308765 371514 308831 371517
rect 307772 371512 308831 371514
rect 307772 371456 308770 371512
rect 308826 371456 308831 371512
rect 307772 371454 308831 371456
rect 307772 371452 307778 371454
rect 308765 371451 308831 371454
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 282678 371316 282684 371380
rect 282748 371378 282754 371380
rect 282821 371378 282887 371381
rect 282748 371376 282887 371378
rect 282748 371320 282826 371376
rect 282882 371320 282887 371376
rect 282748 371318 282887 371320
rect 282748 371316 282754 371318
rect 282821 371315 282887 371318
rect 289721 371378 289787 371381
rect 323158 371378 323164 371380
rect 289721 371376 323164 371378
rect 289721 371320 289726 371376
rect 289782 371320 323164 371376
rect 289721 371318 323164 371320
rect 289721 371315 289787 371318
rect 323158 371316 323164 371318
rect 323228 371316 323234 371380
rect 316902 370500 316908 370564
rect 316972 370562 316978 370564
rect 376017 370562 376083 370565
rect 316972 370560 376083 370562
rect 316972 370504 376022 370560
rect 376078 370504 376083 370560
rect 316972 370502 376083 370504
rect 316972 370500 316978 370502
rect 376017 370499 376083 370502
rect 311850 370230 321570 370290
rect 286409 370154 286475 370157
rect 285814 370152 286475 370154
rect 285814 370096 286414 370152
rect 286470 370096 286475 370152
rect 285814 370094 286475 370096
rect 222009 369882 222075 369885
rect 285075 369882 285141 369885
rect 285254 369882 285260 369884
rect 222009 369880 285260 369882
rect 222009 369824 222014 369880
rect 222070 369824 285080 369880
rect 285136 369824 285260 369880
rect 222009 369822 285260 369824
rect 222009 369819 222075 369822
rect 285075 369819 285141 369822
rect 285254 369820 285260 369822
rect 285324 369820 285330 369884
rect 285814 369882 285874 370094
rect 286409 370091 286475 370094
rect 285949 370018 286015 370021
rect 287053 370018 287119 370021
rect 311850 370018 311910 370230
rect 312486 370092 312492 370156
rect 312556 370154 312562 370156
rect 313181 370154 313247 370157
rect 312556 370152 313247 370154
rect 312556 370096 313186 370152
rect 313242 370096 313247 370152
rect 312556 370094 313247 370096
rect 312556 370092 312562 370094
rect 313181 370091 313247 370094
rect 315254 370094 319960 370154
rect 285949 370016 311910 370018
rect 285949 369960 285954 370016
rect 286010 369960 287058 370016
rect 287114 369960 311910 370016
rect 285949 369958 311910 369960
rect 285949 369955 286015 369958
rect 287053 369955 287119 369958
rect 315254 369882 315314 370094
rect 285814 369822 315314 369882
rect 286182 369749 286242 369822
rect 315614 369820 315620 369884
rect 315684 369882 315690 369884
rect 315849 369882 315915 369885
rect 315684 369880 315915 369882
rect 315684 369824 315854 369880
rect 315910 369824 315915 369880
rect 315684 369822 315915 369824
rect 315684 369820 315690 369822
rect 315849 369819 315915 369822
rect 319437 369882 319503 369885
rect 319662 369882 319668 369884
rect 319437 369880 319668 369882
rect 319437 369824 319442 369880
rect 319498 369824 319668 369880
rect 319437 369822 319668 369824
rect 319437 369819 319503 369822
rect 319662 369820 319668 369822
rect 319732 369820 319738 369884
rect 319900 369882 319960 370094
rect 321510 370018 321570 370230
rect 331806 370018 331812 370020
rect 321510 369958 331812 370018
rect 331806 369956 331812 369958
rect 331876 369956 331882 370020
rect 335854 369882 335860 369884
rect 319900 369822 335860 369882
rect 335854 369820 335860 369822
rect 335924 369820 335930 369884
rect 282126 369684 282132 369748
rect 282196 369746 282202 369748
rect 286179 369746 286245 369749
rect 282196 369744 286245 369746
rect 282196 369688 286184 369744
rect 286240 369688 286245 369744
rect 282196 369686 286245 369688
rect 282196 369684 282202 369686
rect 286179 369683 286245 369686
rect 286915 369746 286981 369749
rect 287053 369746 287119 369749
rect 286915 369744 287119 369746
rect 286915 369688 286920 369744
rect 286976 369688 287058 369744
rect 287114 369688 287119 369744
rect 286915 369686 287119 369688
rect 286915 369683 286981 369686
rect 287053 369683 287119 369686
rect 303475 369746 303541 369749
rect 303981 369746 304047 369749
rect 303475 369744 304047 369746
rect 303475 369688 303480 369744
rect 303536 369688 303986 369744
rect 304042 369688 304047 369744
rect 303475 369686 304047 369688
rect 303475 369683 303541 369686
rect 303981 369683 304047 369686
rect 286918 369610 286978 369683
rect 277350 369550 286978 369610
rect 227069 369202 227135 369205
rect 277350 369202 277410 369550
rect 319294 369548 319300 369612
rect 319364 369610 319370 369612
rect 319805 369610 319871 369613
rect 319364 369608 319871 369610
rect 319364 369552 319810 369608
rect 319866 369552 319871 369608
rect 319364 369550 319871 369552
rect 319364 369548 319370 369550
rect 319805 369547 319871 369550
rect 281574 369412 281580 369476
rect 281644 369474 281650 369476
rect 282678 369474 282684 369476
rect 281644 369414 282684 369474
rect 281644 369412 281650 369414
rect 282678 369412 282684 369414
rect 282748 369474 282754 369476
rect 284477 369474 284543 369477
rect 282748 369472 284543 369474
rect 282748 369416 284482 369472
rect 284538 369416 284543 369472
rect 282748 369414 284543 369416
rect 282748 369412 282754 369414
rect 284477 369411 284543 369414
rect 286542 369412 286548 369476
rect 286612 369474 286618 369476
rect 286777 369474 286843 369477
rect 287283 369476 287349 369477
rect 287278 369474 287284 369476
rect 286612 369472 286843 369474
rect 286612 369416 286782 369472
rect 286838 369416 286843 369472
rect 286612 369414 286843 369416
rect 287192 369414 287284 369474
rect 286612 369412 286618 369414
rect 286777 369411 286843 369414
rect 287278 369412 287284 369414
rect 287348 369412 287354 369476
rect 304942 369412 304948 369476
rect 305012 369474 305018 369476
rect 306281 369474 306347 369477
rect 305012 369472 306347 369474
rect 305012 369416 306286 369472
rect 306342 369416 306347 369472
rect 305012 369414 306347 369416
rect 305012 369412 305018 369414
rect 287283 369411 287349 369412
rect 306281 369411 306347 369414
rect 306966 369412 306972 369476
rect 307036 369474 307042 369476
rect 307661 369474 307727 369477
rect 307036 369472 307727 369474
rect 307036 369416 307666 369472
rect 307722 369416 307727 369472
rect 307036 369414 307727 369416
rect 307036 369412 307042 369414
rect 307661 369411 307727 369414
rect 311014 369412 311020 369476
rect 311084 369474 311090 369476
rect 311801 369474 311867 369477
rect 311084 369472 311867 369474
rect 311084 369416 311806 369472
rect 311862 369416 311867 369472
rect 311084 369414 311867 369416
rect 311084 369412 311090 369414
rect 311801 369411 311867 369414
rect 312307 369472 312373 369477
rect 312307 369416 312312 369472
rect 312368 369416 312373 369472
rect 312307 369411 312373 369416
rect 313774 369412 313780 369476
rect 313844 369474 313850 369476
rect 314377 369474 314443 369477
rect 313844 369472 314443 369474
rect 313844 369416 314382 369472
rect 314438 369416 314443 369472
rect 313844 369414 314443 369416
rect 313844 369412 313850 369414
rect 314377 369411 314443 369414
rect 318006 369412 318012 369476
rect 318076 369474 318082 369476
rect 318425 369474 318491 369477
rect 319897 369476 319963 369477
rect 319846 369474 319852 369476
rect 318076 369472 318491 369474
rect 318076 369416 318430 369472
rect 318486 369416 318491 369472
rect 318076 369414 318491 369416
rect 319806 369414 319852 369474
rect 319916 369472 319963 369476
rect 319958 369416 319963 369472
rect 318076 369412 318082 369414
rect 318425 369411 318491 369414
rect 319846 369412 319852 369414
rect 319916 369412 319963 369416
rect 320766 369412 320772 369476
rect 320836 369474 320842 369476
rect 321369 369474 321435 369477
rect 320836 369472 321435 369474
rect 320836 369416 321374 369472
rect 321430 369416 321435 369472
rect 320836 369414 321435 369416
rect 320836 369412 320842 369414
rect 319897 369411 319963 369412
rect 321369 369411 321435 369414
rect 322054 369412 322060 369476
rect 322124 369474 322130 369476
rect 322841 369474 322907 369477
rect 322124 369472 322907 369474
rect 322124 369416 322846 369472
rect 322902 369416 322907 369472
rect 322124 369414 322907 369416
rect 322124 369412 322130 369414
rect 322841 369411 322907 369414
rect 312310 369341 312370 369411
rect 278630 369276 278636 369340
rect 278700 369338 278706 369340
rect 288019 369338 288085 369341
rect 278700 369336 288085 369338
rect 278700 369280 288024 369336
rect 288080 369280 288085 369336
rect 278700 369278 288085 369280
rect 278700 369276 278706 369278
rect 288019 369275 288085 369278
rect 288934 369276 288940 369340
rect 289004 369338 289010 369340
rect 289123 369338 289189 369341
rect 312307 369338 312373 369341
rect 289004 369336 289189 369338
rect 289004 369280 289128 369336
rect 289184 369280 289189 369336
rect 289004 369278 289189 369280
rect 289004 369276 289010 369278
rect 289123 369275 289189 369278
rect 292530 369336 312373 369338
rect 292530 369280 312312 369336
rect 312368 369280 312373 369336
rect 292530 369278 312373 369280
rect 227069 369200 277410 369202
rect 227069 369144 227074 369200
rect 227130 369144 277410 369200
rect 227069 369142 277410 369144
rect 227069 369139 227135 369142
rect 251817 369066 251883 369069
rect 292530 369066 292590 369278
rect 312307 369275 312373 369278
rect 251817 369064 292590 369066
rect 251817 369008 251822 369064
rect 251878 369008 292590 369064
rect 251817 369006 292590 369008
rect 251817 369003 251883 369006
rect 315430 369004 315436 369068
rect 315500 369066 315506 369068
rect 375925 369066 375991 369069
rect 315500 369064 375991 369066
rect 315500 369008 375930 369064
rect 375986 369008 375991 369064
rect 315500 369006 375991 369008
rect 315500 369004 315506 369006
rect 375925 369003 375991 369006
rect 229737 368930 229803 368933
rect 229737 368928 282194 368930
rect 229737 368872 229742 368928
rect 229798 368872 282194 368928
rect 229737 368870 282194 368872
rect 229737 368867 229803 368870
rect 276013 368658 276079 368661
rect 276473 368658 276539 368661
rect 278630 368658 278636 368660
rect 276013 368656 278636 368658
rect 276013 368600 276018 368656
rect 276074 368600 276478 368656
rect 276534 368600 278636 368656
rect 276013 368598 278636 368600
rect 276013 368595 276079 368598
rect 276473 368595 276539 368598
rect 278630 368596 278636 368598
rect 278700 368596 278706 368660
rect 282134 368658 282194 368870
rect 285254 368732 285260 368796
rect 285324 368794 285330 368796
rect 333881 368794 333947 368797
rect 285324 368792 333947 368794
rect 285324 368736 333886 368792
rect 333942 368736 333947 368792
rect 285324 368734 333947 368736
rect 285324 368732 285330 368734
rect 333881 368731 333947 368734
rect 288934 368658 288940 368660
rect 282134 368598 288940 368658
rect 288934 368596 288940 368598
rect 289004 368658 289010 368660
rect 338757 368658 338823 368661
rect 289004 368656 338823 368658
rect 289004 368600 338762 368656
rect 338818 368600 338823 368656
rect 289004 368598 338823 368600
rect 289004 368596 289010 368598
rect 338757 368595 338823 368598
rect 287278 368460 287284 368524
rect 287348 368522 287354 368524
rect 337377 368522 337443 368525
rect 287348 368520 337443 368522
rect 287348 368464 337382 368520
rect 337438 368464 337443 368520
rect 287348 368462 337443 368464
rect 287348 368460 287354 368462
rect 337377 368459 337443 368462
rect 248413 367706 248479 367709
rect 307702 367706 307708 367708
rect 248413 367704 307708 367706
rect 248413 367648 248418 367704
rect 248474 367648 307708 367704
rect 248413 367646 307708 367648
rect 248413 367643 248479 367646
rect 307702 367644 307708 367646
rect 307772 367644 307778 367708
rect 321134 367644 321140 367708
rect 321204 367706 321210 367708
rect 379646 367706 379652 367708
rect 321204 367646 379652 367706
rect 321204 367644 321210 367646
rect 379646 367644 379652 367646
rect 379716 367644 379722 367708
rect 250621 366346 250687 366349
rect 280470 366346 280476 366348
rect 250621 366344 280476 366346
rect 250621 366288 250626 366344
rect 250682 366288 280476 366344
rect 250621 366286 280476 366288
rect 250621 366283 250687 366286
rect 280470 366284 280476 366286
rect 280540 366284 280546 366348
rect 323158 366284 323164 366348
rect 323228 366346 323234 366348
rect 580441 366346 580507 366349
rect 323228 366344 580507 366346
rect 323228 366288 580446 366344
rect 580502 366288 580507 366344
rect 323228 366286 580507 366288
rect 323228 366284 323234 366286
rect 580441 366283 580507 366286
rect 328361 365666 328427 365669
rect 340045 365666 340111 365669
rect 328361 365664 340111 365666
rect 328361 365608 328366 365664
rect 328422 365608 340050 365664
rect 340106 365608 340111 365664
rect 328361 365606 340111 365608
rect 328361 365603 328427 365606
rect 340045 365603 340111 365606
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 340045 364986 340111 364989
rect 340781 364986 340847 364989
rect 580257 364986 580323 364989
rect 340045 364984 580323 364986
rect 340045 364928 340050 364984
rect 340106 364928 340786 364984
rect 340842 364928 580262 364984
rect 580318 364928 580323 364984
rect 583520 364972 584960 365062
rect 340045 364926 580323 364928
rect 340045 364923 340111 364926
rect 340781 364923 340847 364926
rect 580257 364923 580323 364926
rect 373901 364444 373967 364445
rect 373901 364442 373948 364444
rect 373856 364440 373948 364442
rect 374012 364442 374018 364444
rect 373856 364384 373906 364440
rect 373856 364382 373948 364384
rect 373901 364380 373948 364382
rect 374012 364382 374094 364442
rect 374012 364380 374018 364382
rect 373901 364379 373967 364380
rect 373901 364306 373967 364309
rect 373856 364304 374010 364306
rect 373856 364248 373906 364304
rect 373962 364248 374010 364304
rect 373856 364246 374010 364248
rect 373901 364243 374010 364246
rect 373950 364172 374010 364243
rect 373942 364108 373948 364172
rect 374012 364108 374018 364172
rect 247677 363626 247743 363629
rect 281993 363626 282059 363629
rect 247677 363624 282059 363626
rect 247677 363568 247682 363624
rect 247738 363568 281998 363624
rect 282054 363568 282059 363624
rect 247677 363566 282059 363568
rect 247677 363563 247743 363566
rect 281993 363563 282059 363566
rect 279877 361858 279943 361861
rect 281574 361858 281580 361860
rect 279877 361856 281580 361858
rect 279877 361800 279882 361856
rect 279938 361800 281580 361856
rect 279877 361798 281580 361800
rect 279877 361795 279943 361798
rect 281574 361796 281580 361798
rect 281644 361796 281650 361860
rect 278037 361722 278103 361725
rect 282177 361722 282243 361725
rect 278037 361720 282243 361722
rect 278037 361664 278042 361720
rect 278098 361664 282182 361720
rect 282238 361664 282243 361720
rect 278037 361662 282243 361664
rect 278037 361659 278103 361662
rect 282177 361659 282243 361662
rect 251909 361042 251975 361045
rect 280654 361042 280660 361044
rect 251909 361040 280660 361042
rect 251909 360984 251914 361040
rect 251970 360984 280660 361040
rect 251909 360982 280660 360984
rect 251909 360979 251975 360982
rect 280654 360980 280660 360982
rect 280724 360980 280730 361044
rect 225597 360906 225663 360909
rect 282126 360906 282132 360908
rect 225597 360904 282132 360906
rect 225597 360848 225602 360904
rect 225658 360848 282132 360904
rect 225597 360846 282132 360848
rect 225597 360843 225663 360846
rect 282126 360844 282132 360846
rect 282196 360844 282202 360908
rect 327717 360906 327783 360909
rect 580533 360906 580599 360909
rect 327717 360904 580599 360906
rect 327717 360848 327722 360904
rect 327778 360848 580538 360904
rect 580594 360848 580599 360904
rect 327717 360846 580599 360848
rect 327717 360843 327783 360846
rect 580533 360843 580599 360846
rect 225689 359410 225755 359413
rect 279918 359410 279924 359412
rect 225689 359408 279924 359410
rect 225689 359352 225694 359408
rect 225750 359352 279924 359408
rect 225689 359350 279924 359352
rect 225689 359347 225755 359350
rect 279918 359348 279924 359350
rect 279988 359410 279994 359412
rect 280654 359410 280660 359412
rect 279988 359350 280660 359410
rect 279988 359348 279994 359350
rect 280654 359348 280660 359350
rect 280724 359348 280730 359412
rect 327717 359410 327783 359413
rect 350717 359410 350783 359413
rect 327717 359408 350783 359410
rect 327717 359352 327722 359408
rect 327778 359352 350722 359408
rect 350778 359352 350783 359408
rect 327717 359350 350783 359352
rect 327717 359347 327783 359350
rect 350717 359347 350783 359350
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 327809 358050 327875 358053
rect 349337 358050 349403 358053
rect 327809 358048 349403 358050
rect 327809 357992 327814 358048
rect 327870 357992 349342 358048
rect 349398 357992 349403 358048
rect 327809 357990 349403 357992
rect 327809 357987 327875 357990
rect 349337 357987 349403 357990
rect 327441 355330 327507 355333
rect 386965 355330 387031 355333
rect 327441 355328 387031 355330
rect 327441 355272 327446 355328
rect 327502 355272 386970 355328
rect 387026 355272 387031 355328
rect 327441 355270 387031 355272
rect 327441 355267 327507 355270
rect 386965 355267 387031 355270
rect 373901 354788 373967 354789
rect 373901 354786 373948 354788
rect 373856 354784 373948 354786
rect 374012 354786 374018 354788
rect 373856 354728 373906 354784
rect 373856 354726 373948 354728
rect 373901 354724 373948 354726
rect 374012 354726 374094 354786
rect 374012 354724 374018 354726
rect 373901 354723 373967 354724
rect 373901 354650 373967 354653
rect 373856 354648 374010 354650
rect 373856 354592 373906 354648
rect 373962 354592 374010 354648
rect 373856 354590 374010 354592
rect 373901 354587 374010 354590
rect 373950 354516 374010 354587
rect 373942 354452 373948 354516
rect 374012 354452 374018 354516
rect 247769 352610 247835 352613
rect 282453 352610 282519 352613
rect 247769 352608 282519 352610
rect 247769 352552 247774 352608
rect 247830 352552 282458 352608
rect 282514 352552 282519 352608
rect 247769 352550 282519 352552
rect 247769 352547 247835 352550
rect 282453 352547 282519 352550
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect 327901 351114 327967 351117
rect 374177 351114 374243 351117
rect 327901 351112 374243 351114
rect 327901 351056 327906 351112
rect 327962 351056 374182 351112
rect 374238 351056 374243 351112
rect 327901 351054 374243 351056
rect 327901 351051 327967 351054
rect 374177 351051 374243 351054
rect 325366 345612 325372 345676
rect 325436 345674 325442 345676
rect 381670 345674 381676 345676
rect 325436 345614 381676 345674
rect 325436 345612 325442 345614
rect 381670 345612 381676 345614
rect 381740 345612 381746 345676
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 373901 345132 373967 345133
rect 373901 345130 373948 345132
rect 373856 345128 373948 345130
rect 374012 345130 374018 345132
rect 373856 345072 373906 345128
rect 373856 345070 373948 345072
rect 373901 345068 373948 345070
rect 374012 345070 374094 345130
rect 374012 345068 374018 345070
rect 373901 345067 373967 345068
rect 373901 344996 373967 344997
rect 373901 344994 373948 344996
rect 373856 344992 373948 344994
rect 374012 344994 374018 344996
rect 373856 344936 373906 344992
rect 373856 344934 373948 344936
rect 373901 344932 373948 344934
rect 374012 344934 374094 344994
rect 374012 344932 374018 344934
rect 373901 344931 373967 344932
rect 324262 342892 324268 342956
rect 324332 342954 324338 342956
rect 382774 342954 382780 342956
rect 324332 342894 382780 342954
rect 324332 342892 324338 342894
rect 382774 342892 382780 342894
rect 382844 342892 382850 342956
rect 373901 340780 373967 340781
rect 373901 340776 373948 340780
rect 374012 340778 374018 340780
rect 373901 340720 373906 340776
rect 373901 340716 373948 340720
rect 374012 340718 374058 340778
rect 374012 340716 374018 340718
rect 373901 340715 373967 340716
rect 583520 338452 584960 338692
rect 340689 337378 340755 337381
rect 379278 337378 379284 337380
rect 340689 337376 379284 337378
rect 340689 337320 340694 337376
rect 340750 337320 379284 337376
rect 340689 337318 379284 337320
rect 340689 337315 340755 337318
rect 379278 337316 379284 337318
rect 379348 337316 379354 337380
rect -960 332196 480 332436
rect 373901 331260 373967 331261
rect 373901 331258 373948 331260
rect 373856 331256 373948 331258
rect 373856 331200 373906 331256
rect 373856 331198 373948 331200
rect 373901 331196 373948 331198
rect 374012 331196 374018 331260
rect 373901 331195 373967 331196
rect 225781 330442 225847 330445
rect 276606 330442 276612 330444
rect 225781 330440 276612 330442
rect 225781 330384 225786 330440
rect 225842 330384 276612 330440
rect 225781 330382 276612 330384
rect 225781 330379 225847 330382
rect 276606 330380 276612 330382
rect 276676 330380 276682 330444
rect 327533 330442 327599 330445
rect 386781 330442 386847 330445
rect 327533 330440 386847 330442
rect 327533 330384 327538 330440
rect 327594 330384 386786 330440
rect 386842 330384 386847 330440
rect 327533 330382 386847 330384
rect 327533 330379 327599 330382
rect 386781 330379 386847 330382
rect 382038 329898 382044 329900
rect 380942 329838 382044 329898
rect 380942 329762 381002 329838
rect 382038 329836 382044 329838
rect 382108 329898 382114 329900
rect 513373 329898 513439 329901
rect 382108 329896 513439 329898
rect 382108 329840 513378 329896
rect 513434 329840 513439 329896
rect 382108 329838 513439 329840
rect 382108 329836 382114 329838
rect 513373 329835 513439 329838
rect 373950 329702 381002 329762
rect 341977 329354 342043 329357
rect 368422 329354 368428 329356
rect 341977 329352 368428 329354
rect 341977 329296 341982 329352
rect 342038 329296 368428 329352
rect 341977 329294 368428 329296
rect 341977 329291 342043 329294
rect 368422 329292 368428 329294
rect 368492 329292 368498 329356
rect 335261 329218 335327 329221
rect 373950 329218 374010 329702
rect 335261 329216 374010 329218
rect 335261 329160 335266 329216
rect 335322 329160 374010 329216
rect 335261 329158 374010 329160
rect 335261 329155 335327 329158
rect 338246 329082 338252 329084
rect 335310 329022 338252 329082
rect 326838 328476 326844 328540
rect 326908 328538 326914 328540
rect 335310 328538 335370 329022
rect 338246 329020 338252 329022
rect 338316 329082 338322 329084
rect 386965 329082 387031 329085
rect 338316 329080 387031 329082
rect 338316 329024 386970 329080
rect 387026 329024 387031 329080
rect 338316 329022 387031 329024
rect 338316 329020 338322 329022
rect 386965 329019 387031 329022
rect 326908 328478 335370 328538
rect 326908 328476 326914 328478
rect 375230 328476 375236 328540
rect 375300 328538 375306 328540
rect 416773 328538 416839 328541
rect 375300 328536 416839 328538
rect 375300 328480 416778 328536
rect 416834 328480 416839 328536
rect 375300 328478 416839 328480
rect 375300 328476 375306 328478
rect 416773 328475 416839 328478
rect 337929 327722 337995 327725
rect 375230 327722 375236 327724
rect 337929 327720 375236 327722
rect 337929 327664 337934 327720
rect 337990 327664 375236 327720
rect 337929 327662 375236 327664
rect 337929 327659 337995 327662
rect 375230 327660 375236 327662
rect 375300 327660 375306 327724
rect 346301 326634 346367 326637
rect 378174 326634 378180 326636
rect 346301 326632 378180 326634
rect 346301 326576 346306 326632
rect 346362 326576 378180 326632
rect 346301 326574 378180 326576
rect 346301 326571 346367 326574
rect 378174 326572 378180 326574
rect 378244 326572 378250 326636
rect 336457 326498 336523 326501
rect 374126 326498 374132 326500
rect 336457 326496 374132 326498
rect 336457 326440 336462 326496
rect 336518 326440 374132 326496
rect 336457 326438 374132 326440
rect 336457 326435 336523 326438
rect 374126 326436 374132 326438
rect 374196 326436 374202 326500
rect 327574 326300 327580 326364
rect 327644 326362 327650 326364
rect 386689 326362 386755 326365
rect 327644 326360 386755 326362
rect 327644 326304 386694 326360
rect 386750 326304 386755 326360
rect 327644 326302 386755 326304
rect 327644 326300 327650 326302
rect 386689 326299 386755 326302
rect 373942 325892 373948 325956
rect 374012 325892 374018 325956
rect 373950 325821 374010 325892
rect 323342 325756 323348 325820
rect 323412 325818 323418 325820
rect 345013 325818 345079 325821
rect 346301 325818 346367 325821
rect 373901 325818 374010 325821
rect 323412 325816 346367 325818
rect 323412 325760 345018 325816
rect 345074 325760 346306 325816
rect 346362 325760 346367 325816
rect 323412 325758 346367 325760
rect 373856 325816 374010 325818
rect 373856 325760 373906 325816
rect 373962 325760 374010 325816
rect 373856 325758 374010 325760
rect 323412 325756 323418 325758
rect 345013 325755 345079 325758
rect 346301 325755 346367 325758
rect 373901 325755 373967 325758
rect 344921 325410 344987 325413
rect 371366 325410 371372 325412
rect 344921 325408 371372 325410
rect 344921 325352 344926 325408
rect 344982 325352 371372 325408
rect 344921 325350 371372 325352
rect 344921 325347 344987 325350
rect 371366 325348 371372 325350
rect 371436 325348 371442 325412
rect 338113 325274 338179 325277
rect 374126 325274 374132 325276
rect 338113 325272 374132 325274
rect 338113 325216 338118 325272
rect 338174 325216 374132 325272
rect 338113 325214 374132 325216
rect 338113 325211 338179 325214
rect 374126 325212 374132 325214
rect 374196 325212 374202 325276
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 330334 325076 330340 325140
rect 330404 325138 330410 325140
rect 385309 325138 385375 325141
rect 330404 325136 385375 325138
rect 330404 325080 385314 325136
rect 385370 325080 385375 325136
rect 583520 325124 584960 325214
rect 330404 325078 385375 325080
rect 330404 325076 330410 325078
rect 385309 325075 385375 325078
rect 323526 324940 323532 325004
rect 323596 325002 323602 325004
rect 382222 325002 382228 325004
rect 323596 324942 382228 325002
rect 323596 324940 323602 324942
rect 382222 324940 382228 324942
rect 382292 324940 382298 325004
rect 327758 324396 327764 324460
rect 327828 324458 327834 324460
rect 330334 324458 330340 324460
rect 327828 324398 330340 324458
rect 327828 324396 327834 324398
rect 330334 324396 330340 324398
rect 330404 324396 330410 324460
rect 373758 324396 373764 324460
rect 373828 324458 373834 324460
rect 398925 324458 398991 324461
rect 373828 324456 398991 324458
rect 373828 324400 398930 324456
rect 398986 324400 398991 324456
rect 373828 324398 398991 324400
rect 373828 324396 373834 324398
rect 340965 323778 341031 323781
rect 373950 323778 374010 324398
rect 398925 324395 398991 324398
rect 340965 323776 374010 323778
rect 340965 323720 340970 323776
rect 341026 323720 374010 323776
rect 340965 323718 374010 323720
rect 340965 323715 341031 323718
rect 229921 323642 229987 323645
rect 277894 323642 277900 323644
rect 229921 323640 277900 323642
rect 229921 323584 229926 323640
rect 229982 323584 277900 323640
rect 229921 323582 277900 323584
rect 229921 323579 229987 323582
rect 277894 323580 277900 323582
rect 277964 323580 277970 323644
rect 328177 323642 328243 323645
rect 377765 323642 377831 323645
rect 328177 323640 377831 323642
rect 328177 323584 328182 323640
rect 328238 323584 377770 323640
rect 377826 323584 377831 323640
rect 328177 323582 377831 323584
rect 328177 323579 328243 323582
rect 377765 323579 377831 323582
rect 260465 322962 260531 322965
rect 282085 322962 282151 322965
rect 260465 322960 282151 322962
rect 260465 322904 260470 322960
rect 260526 322904 282090 322960
rect 282146 322904 282151 322960
rect 260465 322902 282151 322904
rect 260465 322899 260531 322902
rect 282085 322899 282151 322902
rect 323710 322900 323716 322964
rect 323780 322962 323786 322964
rect 331213 322962 331279 322965
rect 323780 322960 331279 322962
rect 323780 322904 331218 322960
rect 331274 322904 331279 322960
rect 323780 322902 331279 322904
rect 323780 322900 323786 322902
rect 331213 322899 331279 322902
rect 228541 322282 228607 322285
rect 279550 322282 279556 322284
rect 228541 322280 279556 322282
rect 228541 322224 228546 322280
rect 228602 322224 279556 322280
rect 228541 322222 279556 322224
rect 228541 322219 228607 322222
rect 279550 322220 279556 322222
rect 279620 322220 279626 322284
rect 204161 322146 204227 322149
rect 276657 322146 276723 322149
rect 281901 322146 281967 322149
rect 331305 322146 331371 322149
rect 204161 322144 281967 322146
rect 204161 322088 204166 322144
rect 204222 322088 276662 322144
rect 276718 322088 281906 322144
rect 281962 322088 281967 322144
rect 204161 322086 281967 322088
rect 204161 322083 204227 322086
rect 276657 322083 276723 322086
rect 281901 322083 281967 322086
rect 323166 322144 331371 322146
rect 323166 322088 331310 322144
rect 331366 322088 331371 322144
rect 323166 322086 331371 322088
rect 288934 321948 288940 322012
rect 289004 322010 289010 322012
rect 293350 322010 293356 322012
rect 289004 321950 293356 322010
rect 289004 321948 289010 321950
rect 293350 321948 293356 321950
rect 293420 321948 293426 322012
rect 321686 321948 321692 322012
rect 321756 322010 321762 322012
rect 323166 322010 323226 322086
rect 331305 322083 331371 322086
rect 321756 321950 323226 322010
rect 321756 321948 321762 321950
rect 325182 321948 325188 322012
rect 325252 322010 325258 322012
rect 332685 322010 332751 322013
rect 325252 322008 332751 322010
rect 325252 321952 332690 322008
rect 332746 321952 332751 322008
rect 325252 321950 332751 321952
rect 325252 321948 325258 321950
rect 332685 321947 332751 321950
rect 279233 321874 279299 321877
rect 282678 321874 282684 321876
rect 279233 321872 282684 321874
rect 279233 321816 279238 321872
rect 279294 321816 282684 321872
rect 279233 321814 282684 321816
rect 279233 321811 279299 321814
rect 282678 321812 282684 321814
rect 282748 321874 282754 321876
rect 284334 321874 284340 321876
rect 282748 321814 284340 321874
rect 282748 321812 282754 321814
rect 284334 321812 284340 321814
rect 284404 321812 284410 321876
rect 288566 321812 288572 321876
rect 288636 321874 288642 321876
rect 298318 321874 298324 321876
rect 288636 321814 298324 321874
rect 288636 321812 288642 321814
rect 298318 321812 298324 321814
rect 298388 321812 298394 321876
rect 324078 321812 324084 321876
rect 324148 321874 324154 321876
rect 330385 321874 330451 321877
rect 330702 321874 330708 321876
rect 324148 321872 330708 321874
rect 324148 321816 330390 321872
rect 330446 321816 330708 321872
rect 324148 321814 330708 321816
rect 324148 321812 324154 321814
rect 330385 321811 330451 321814
rect 330702 321812 330708 321814
rect 330772 321812 330778 321876
rect 219341 321738 219407 321741
rect 281993 321738 282059 321741
rect 301262 321738 301268 321740
rect 219341 321736 279434 321738
rect 219341 321680 219346 321736
rect 219402 321680 279434 321736
rect 219341 321678 279434 321680
rect 219341 321675 219407 321678
rect 205541 321602 205607 321605
rect 279233 321602 279299 321605
rect 205541 321600 279299 321602
rect 205541 321544 205546 321600
rect 205602 321544 279238 321600
rect 279294 321544 279299 321600
rect 205541 321542 279299 321544
rect 279374 321602 279434 321678
rect 281993 321736 301268 321738
rect 281993 321680 281998 321736
rect 282054 321680 301268 321736
rect 281993 321678 301268 321680
rect 281993 321675 282059 321678
rect 301262 321676 301268 321678
rect 301332 321676 301338 321740
rect 321502 321676 321508 321740
rect 321572 321738 321578 321740
rect 338205 321738 338271 321741
rect 378041 321738 378107 321741
rect 321572 321736 378107 321738
rect 321572 321680 338210 321736
rect 338266 321680 378046 321736
rect 378102 321680 378107 321736
rect 321572 321678 378107 321680
rect 321572 321676 321578 321678
rect 338205 321675 338271 321678
rect 378041 321675 378107 321678
rect 282361 321602 282427 321605
rect 282678 321602 282684 321604
rect 279374 321600 282684 321602
rect 279374 321544 282366 321600
rect 282422 321544 282684 321600
rect 279374 321542 282684 321544
rect 205541 321539 205607 321542
rect 279233 321539 279299 321542
rect 282361 321539 282427 321542
rect 282678 321540 282684 321542
rect 282748 321540 282754 321604
rect 284518 321540 284524 321604
rect 284588 321602 284594 321604
rect 286358 321602 286364 321604
rect 284588 321542 286364 321602
rect 284588 321540 284594 321542
rect 286358 321540 286364 321542
rect 286428 321540 286434 321604
rect 290590 321540 290596 321604
rect 290660 321602 290666 321604
rect 299054 321602 299060 321604
rect 290660 321542 299060 321602
rect 290660 321540 290666 321542
rect 299054 321540 299060 321542
rect 299124 321540 299130 321604
rect 326654 321540 326660 321604
rect 326724 321602 326730 321604
rect 330518 321602 330524 321604
rect 326724 321542 330524 321602
rect 326724 321540 326730 321542
rect 330518 321540 330524 321542
rect 330588 321602 330594 321604
rect 386597 321602 386663 321605
rect 387057 321602 387123 321605
rect 330588 321600 387123 321602
rect 330588 321544 386602 321600
rect 386658 321544 387062 321600
rect 387118 321544 387123 321600
rect 330588 321542 387123 321544
rect 330588 321540 330594 321542
rect 386597 321539 386663 321542
rect 387057 321539 387123 321542
rect 282453 321466 282519 321469
rect 282453 321464 291026 321466
rect 282453 321408 282458 321464
rect 282514 321408 291026 321464
rect 282453 321406 291026 321408
rect 282453 321403 282519 321406
rect 279509 321330 279575 321333
rect 288934 321330 288940 321332
rect 279509 321328 288940 321330
rect 279509 321272 279514 321328
rect 279570 321272 288940 321328
rect 279509 321270 288940 321272
rect 279509 321267 279575 321270
rect 288934 321268 288940 321270
rect 289004 321268 289010 321332
rect 290966 321330 291026 321406
rect 291142 321404 291148 321468
rect 291212 321466 291218 321468
rect 291212 321406 316786 321466
rect 291212 321404 291218 321406
rect 292614 321330 292620 321332
rect 290966 321270 292620 321330
rect 292614 321268 292620 321270
rect 292684 321268 292690 321332
rect 293350 321268 293356 321332
rect 293420 321330 293426 321332
rect 314510 321330 314516 321332
rect 293420 321270 314516 321330
rect 293420 321268 293426 321270
rect 314510 321268 314516 321270
rect 314580 321268 314586 321332
rect 316726 321330 316786 321406
rect 320214 321404 320220 321468
rect 320284 321466 320290 321468
rect 328361 321466 328427 321469
rect 320284 321464 328427 321466
rect 320284 321408 328366 321464
rect 328422 321408 328427 321464
rect 320284 321406 328427 321408
rect 320284 321404 320290 321406
rect 328361 321403 328427 321406
rect 335813 321330 335879 321333
rect 350758 321330 350764 321332
rect 316726 321270 321570 321330
rect 281993 321194 282059 321197
rect 290958 321194 290964 321196
rect 281993 321192 289600 321194
rect 281993 321136 281998 321192
rect 282054 321136 289600 321192
rect 281993 321134 289600 321136
rect 281993 321131 282059 321134
rect 276749 321058 276815 321061
rect 282453 321058 282519 321061
rect 276749 321056 282519 321058
rect 276749 321000 276754 321056
rect 276810 321000 282458 321056
rect 282514 321000 282519 321056
rect 276749 320998 282519 321000
rect 276749 320995 276815 320998
rect 282453 320995 282519 320998
rect 283230 320996 283236 321060
rect 283300 321058 283306 321060
rect 288566 321058 288572 321060
rect 283300 320998 288572 321058
rect 283300 320996 283306 320998
rect 288566 320996 288572 320998
rect 288636 320996 288642 321060
rect 277853 320922 277919 320925
rect 288382 320922 288388 320924
rect 277853 320920 288388 320922
rect 277853 320864 277858 320920
rect 277914 320864 288388 320920
rect 277853 320862 288388 320864
rect 277853 320859 277919 320862
rect 285538 320789 285598 320862
rect 288382 320860 288388 320862
rect 288452 320860 288458 320924
rect 275093 320786 275159 320789
rect 275369 320786 275435 320789
rect 280153 320786 280219 320789
rect 282683 320788 282749 320789
rect 283971 320788 284037 320789
rect 282678 320786 282684 320788
rect 275093 320784 278514 320786
rect 275093 320728 275098 320784
rect 275154 320728 275374 320784
rect 275430 320728 278514 320784
rect 275093 320726 278514 320728
rect 275093 320723 275159 320726
rect 275369 320723 275435 320726
rect 273897 320650 273963 320653
rect 278221 320650 278287 320653
rect 273897 320648 278287 320650
rect 273897 320592 273902 320648
rect 273958 320592 278226 320648
rect 278282 320592 278287 320648
rect 273897 320590 278287 320592
rect 278454 320650 278514 320726
rect 280153 320784 282516 320786
rect 280153 320728 280158 320784
rect 280214 320728 282516 320784
rect 280153 320726 282516 320728
rect 282592 320726 282684 320786
rect 280153 320723 280219 320726
rect 281993 320650 282059 320653
rect 278454 320648 282059 320650
rect 278454 320592 281998 320648
rect 282054 320592 282059 320648
rect 278454 320590 282059 320592
rect 282456 320650 282516 320726
rect 282678 320724 282684 320726
rect 282748 320724 282754 320788
rect 283966 320786 283972 320788
rect 283880 320726 283972 320786
rect 283966 320724 283972 320726
rect 284036 320724 284042 320788
rect 284339 320786 284405 320789
rect 285070 320786 285076 320788
rect 284339 320784 285076 320786
rect 284339 320728 284344 320784
rect 284400 320728 285076 320784
rect 284339 320726 285076 320728
rect 282683 320723 282749 320724
rect 283971 320723 284037 320724
rect 284339 320723 284405 320726
rect 285070 320724 285076 320726
rect 285140 320724 285146 320788
rect 285535 320784 285601 320789
rect 285535 320728 285540 320784
rect 285596 320728 285601 320784
rect 285535 320723 285601 320728
rect 287462 320724 287468 320788
rect 287532 320786 287538 320788
rect 288198 320786 288204 320788
rect 287532 320726 288204 320786
rect 287532 320724 287538 320726
rect 288198 320724 288204 320726
rect 288268 320786 288274 320788
rect 288387 320786 288453 320789
rect 288268 320784 288453 320786
rect 288268 320728 288392 320784
rect 288448 320728 288453 320784
rect 288268 320726 288453 320728
rect 288268 320724 288274 320726
rect 288387 320723 288453 320726
rect 288566 320724 288572 320788
rect 288636 320786 288642 320788
rect 289123 320786 289189 320789
rect 289307 320788 289373 320789
rect 288636 320784 289189 320786
rect 288636 320728 289128 320784
rect 289184 320728 289189 320784
rect 288636 320726 289189 320728
rect 288636 320724 288642 320726
rect 289123 320723 289189 320726
rect 289302 320724 289308 320788
rect 289372 320786 289378 320788
rect 289372 320726 289464 320786
rect 289372 320724 289378 320726
rect 289307 320723 289373 320724
rect 284707 320652 284773 320653
rect 284702 320650 284708 320652
rect 282456 320590 284708 320650
rect 273897 320587 273963 320590
rect 278221 320587 278287 320590
rect 281993 320587 282059 320590
rect 284702 320588 284708 320590
rect 284772 320588 284778 320652
rect 284886 320588 284892 320652
rect 284956 320650 284962 320652
rect 285075 320650 285141 320653
rect 284956 320648 285141 320650
rect 284956 320592 285080 320648
rect 285136 320592 285141 320648
rect 284956 320590 285141 320592
rect 284956 320588 284962 320590
rect 284707 320587 284773 320588
rect 285075 320587 285141 320590
rect 287462 320588 287468 320652
rect 287532 320650 287538 320652
rect 288295 320650 288361 320653
rect 287532 320648 288361 320650
rect 287532 320592 288300 320648
rect 288356 320592 288361 320648
rect 287532 320590 288361 320592
rect 289540 320650 289600 321134
rect 289862 321134 290964 321194
rect 289862 320789 289922 321134
rect 290958 321132 290964 321134
rect 291028 321132 291034 321196
rect 294270 321132 294276 321196
rect 294340 321194 294346 321196
rect 295006 321194 295012 321196
rect 294340 321134 295012 321194
rect 294340 321132 294346 321134
rect 295006 321132 295012 321134
rect 295076 321132 295082 321196
rect 321510 321194 321570 321270
rect 335813 321328 350764 321330
rect 335813 321272 335818 321328
rect 335874 321272 350764 321328
rect 335813 321270 350764 321272
rect 335813 321267 335879 321270
rect 350758 321268 350764 321270
rect 350828 321268 350834 321332
rect 346117 321194 346183 321197
rect 321510 321192 346183 321194
rect 321510 321136 346122 321192
rect 346178 321136 346183 321192
rect 321510 321134 346183 321136
rect 346117 321131 346183 321134
rect 298318 320996 298324 321060
rect 298388 321058 298394 321060
rect 343449 321058 343515 321061
rect 298388 321056 343515 321058
rect 298388 321000 343454 321056
rect 343510 321000 343515 321056
rect 298388 320998 343515 321000
rect 298388 320996 298394 320998
rect 343449 320995 343515 320998
rect 321502 320922 321508 320924
rect 290966 320862 299490 320922
rect 289859 320784 289925 320789
rect 289859 320728 289864 320784
rect 289920 320728 289925 320784
rect 289859 320723 289925 320728
rect 290966 320650 291026 320862
rect 291423 320786 291489 320789
rect 291878 320786 291884 320788
rect 291423 320784 291884 320786
rect 291423 320728 291428 320784
rect 291484 320728 291884 320784
rect 291423 320726 291884 320728
rect 291423 320723 291489 320726
rect 291878 320724 291884 320726
rect 291948 320724 291954 320788
rect 292614 320724 292620 320788
rect 292684 320786 292690 320788
rect 295379 320786 295445 320789
rect 292684 320784 295445 320786
rect 292684 320728 295384 320784
rect 295440 320728 295445 320784
rect 292684 320726 295445 320728
rect 292684 320724 292690 320726
rect 295379 320723 295445 320726
rect 297035 320786 297101 320789
rect 297214 320786 297220 320788
rect 297035 320784 297220 320786
rect 297035 320728 297040 320784
rect 297096 320728 297220 320784
rect 297035 320726 297220 320728
rect 297035 320723 297101 320726
rect 297214 320724 297220 320726
rect 297284 320724 297290 320788
rect 299238 320786 299244 320788
rect 298326 320726 299244 320786
rect 289540 320590 291026 320650
rect 292159 320650 292225 320653
rect 292430 320650 292436 320652
rect 292159 320648 292436 320650
rect 287532 320588 287538 320590
rect 288295 320587 288361 320590
rect 291334 320556 292038 320616
rect 292159 320592 292164 320648
rect 292220 320592 292436 320648
rect 292159 320590 292436 320592
rect 292159 320587 292225 320590
rect 292430 320588 292436 320590
rect 292500 320588 292506 320652
rect 293166 320588 293172 320652
rect 293236 320650 293242 320652
rect 293447 320650 293513 320653
rect 293236 320648 293513 320650
rect 293236 320592 293452 320648
rect 293508 320592 293513 320648
rect 293236 320590 293513 320592
rect 293236 320588 293242 320590
rect 293447 320587 293513 320590
rect 294091 320650 294157 320653
rect 295558 320650 295564 320652
rect 294091 320648 295564 320650
rect 294091 320592 294096 320648
rect 294152 320592 295564 320648
rect 294091 320590 295564 320592
rect 294091 320587 294157 320590
rect 295558 320588 295564 320590
rect 295628 320588 295634 320652
rect 298139 320650 298205 320653
rect 298326 320652 298386 320726
rect 299238 320724 299244 320726
rect 299308 320724 299314 320788
rect 298507 320652 298573 320653
rect 299243 320652 299309 320653
rect 298318 320650 298324 320652
rect 298139 320648 298324 320650
rect 298139 320592 298144 320648
rect 298200 320592 298324 320648
rect 298139 320590 298324 320592
rect 298139 320587 298205 320590
rect 298318 320588 298324 320590
rect 298388 320588 298394 320652
rect 298502 320588 298508 320652
rect 298572 320650 298578 320652
rect 299238 320650 299244 320652
rect 298572 320590 298664 320650
rect 299152 320590 299244 320650
rect 298572 320588 298578 320590
rect 299238 320588 299244 320590
rect 299308 320588 299314 320652
rect 299430 320650 299490 320862
rect 302190 320862 304090 320922
rect 301267 320788 301333 320789
rect 301262 320786 301268 320788
rect 301176 320726 301268 320786
rect 301262 320724 301268 320726
rect 301332 320724 301338 320788
rect 301267 320723 301333 320724
rect 302190 320650 302250 320862
rect 304030 320789 304090 320862
rect 320038 320862 321508 320922
rect 304027 320784 304093 320789
rect 304763 320788 304829 320789
rect 304758 320786 304764 320788
rect 304027 320728 304032 320784
rect 304088 320728 304093 320784
rect 304027 320723 304093 320728
rect 304672 320726 304764 320786
rect 304758 320724 304764 320726
rect 304828 320724 304834 320788
rect 306414 320724 306420 320788
rect 306484 320786 306490 320788
rect 306966 320786 306972 320788
rect 306484 320726 306972 320786
rect 306484 320724 306490 320726
rect 306966 320724 306972 320726
rect 307036 320786 307042 320788
rect 307523 320786 307589 320789
rect 307036 320784 307589 320786
rect 307036 320728 307528 320784
rect 307584 320728 307589 320784
rect 307036 320726 307589 320728
rect 307036 320724 307042 320726
rect 304763 320723 304829 320724
rect 307523 320723 307589 320726
rect 310646 320724 310652 320788
rect 310716 320786 310722 320788
rect 311111 320786 311177 320789
rect 311750 320786 311756 320788
rect 310716 320784 311756 320786
rect 310716 320728 311116 320784
rect 311172 320728 311756 320784
rect 310716 320726 311756 320728
rect 310716 320724 310722 320726
rect 311111 320723 311177 320726
rect 311750 320724 311756 320726
rect 311820 320724 311826 320788
rect 314510 320724 314516 320788
rect 314580 320786 314586 320788
rect 314791 320786 314857 320789
rect 314580 320784 314857 320786
rect 314580 320728 314796 320784
rect 314852 320728 314857 320784
rect 314580 320726 314857 320728
rect 314580 320724 314586 320726
rect 314791 320723 314857 320726
rect 315430 320724 315436 320788
rect 315500 320786 315506 320788
rect 315803 320786 315869 320789
rect 315500 320784 315869 320786
rect 315500 320728 315808 320784
rect 315864 320728 315869 320784
rect 315500 320726 315869 320728
rect 315500 320724 315506 320726
rect 315803 320723 315869 320726
rect 318471 320786 318537 320789
rect 320038 320786 320098 320862
rect 321502 320860 321508 320862
rect 321572 320860 321578 320924
rect 325550 320922 325556 320924
rect 324638 320862 325556 320922
rect 324638 320789 324698 320862
rect 325550 320860 325556 320862
rect 325620 320922 325626 320924
rect 383929 320922 383995 320925
rect 325620 320920 383995 320922
rect 325620 320864 383934 320920
rect 383990 320864 383995 320920
rect 325620 320862 383995 320864
rect 325620 320860 325626 320862
rect 383929 320859 383995 320862
rect 321691 320788 321757 320789
rect 321686 320786 321692 320788
rect 318471 320784 320098 320786
rect 318471 320728 318476 320784
rect 318532 320728 320098 320784
rect 318471 320726 320098 320728
rect 321600 320726 321692 320786
rect 318471 320723 318537 320726
rect 321686 320724 321692 320726
rect 321756 320724 321762 320788
rect 322054 320724 322060 320788
rect 322124 320786 322130 320788
rect 322427 320786 322493 320789
rect 324083 320788 324149 320789
rect 324078 320786 324084 320788
rect 322124 320784 322493 320786
rect 322124 320728 322432 320784
rect 322488 320728 322493 320784
rect 322124 320726 322493 320728
rect 323992 320726 324084 320786
rect 322124 320724 322130 320726
rect 321691 320723 321757 320724
rect 322427 320723 322493 320726
rect 324078 320724 324084 320726
rect 324148 320724 324154 320788
rect 324635 320784 324701 320789
rect 325187 320788 325253 320789
rect 325182 320786 325188 320788
rect 324635 320728 324640 320784
rect 324696 320728 324701 320784
rect 324083 320723 324149 320724
rect 324635 320723 324701 320728
rect 325096 320726 325188 320786
rect 325182 320724 325188 320726
rect 325252 320724 325258 320788
rect 326475 320786 326541 320789
rect 327395 320788 327461 320789
rect 326654 320786 326660 320788
rect 326475 320784 326660 320786
rect 326475 320728 326480 320784
rect 326536 320728 326660 320784
rect 326475 320726 326660 320728
rect 325187 320723 325253 320724
rect 326475 320723 326541 320726
rect 326654 320724 326660 320726
rect 326724 320724 326730 320788
rect 327390 320786 327396 320788
rect 327268 320726 327396 320786
rect 327460 320786 327466 320788
rect 327625 320786 327691 320789
rect 388161 320786 388227 320789
rect 327460 320784 327691 320786
rect 327460 320728 327630 320784
rect 327686 320728 327691 320784
rect 327390 320724 327396 320726
rect 327460 320726 327691 320728
rect 327460 320724 327466 320726
rect 327395 320723 327461 320724
rect 327625 320723 327691 320726
rect 335310 320784 388227 320786
rect 335310 320728 388166 320784
rect 388222 320728 388227 320784
rect 335310 320726 388227 320728
rect 299430 320590 302250 320650
rect 304022 320588 304028 320652
rect 304092 320650 304098 320652
rect 304487 320650 304553 320653
rect 304092 320648 304553 320650
rect 304092 320592 304492 320648
rect 304548 320592 304553 320648
rect 304092 320590 304553 320592
rect 304092 320588 304098 320590
rect 298507 320587 298573 320588
rect 299243 320587 299309 320588
rect 304487 320587 304553 320590
rect 305315 320650 305381 320653
rect 305862 320650 305868 320652
rect 305315 320648 305868 320650
rect 305315 320592 305320 320648
rect 305376 320592 305868 320648
rect 305315 320590 305868 320592
rect 305315 320587 305381 320590
rect 305862 320588 305868 320590
rect 305932 320588 305938 320652
rect 307615 320648 307681 320653
rect 307615 320592 307620 320648
rect 307676 320592 307681 320648
rect 307615 320587 307681 320592
rect 313590 320588 313596 320652
rect 313660 320650 313666 320652
rect 313779 320650 313845 320653
rect 313660 320648 313845 320650
rect 313660 320592 313784 320648
rect 313840 320592 313845 320648
rect 313660 320590 313845 320592
rect 313660 320588 313666 320590
rect 313779 320587 313845 320590
rect 317827 320650 317893 320653
rect 320214 320650 320220 320652
rect 317827 320648 320220 320650
rect 317827 320592 317832 320648
rect 317888 320592 320220 320648
rect 317827 320590 320220 320592
rect 317827 320587 317893 320590
rect 320214 320588 320220 320590
rect 320284 320588 320290 320652
rect 324814 320588 324820 320652
rect 324884 320650 324890 320652
rect 326751 320650 326817 320653
rect 324884 320590 325066 320650
rect 324884 320588 324890 320590
rect 269481 320514 269547 320517
rect 270033 320514 270099 320517
rect 291334 320514 291394 320556
rect 269481 320512 288818 320514
rect 269481 320456 269486 320512
rect 269542 320456 270038 320512
rect 270094 320456 288818 320512
rect 269481 320454 288818 320456
rect 269481 320451 269547 320454
rect 270033 320451 270099 320454
rect 271137 320378 271203 320381
rect 288758 320378 288818 320454
rect 289494 320454 291394 320514
rect 291978 320514 292038 320556
rect 299979 320514 300045 320517
rect 291978 320512 300045 320514
rect 291978 320456 299984 320512
rect 300040 320456 300045 320512
rect 291978 320454 300045 320456
rect 289494 320378 289554 320454
rect 299979 320451 300045 320454
rect 300342 320452 300348 320516
rect 300412 320514 300418 320516
rect 300531 320514 300597 320517
rect 300412 320512 300597 320514
rect 300412 320456 300536 320512
rect 300592 320456 300597 320512
rect 300412 320454 300597 320456
rect 300412 320452 300418 320454
rect 300531 320451 300597 320454
rect 301630 320452 301636 320516
rect 301700 320514 301706 320516
rect 302095 320514 302161 320517
rect 301700 320512 302161 320514
rect 301700 320456 302100 320512
rect 302156 320456 302161 320512
rect 301700 320454 302161 320456
rect 301700 320452 301706 320454
rect 302095 320451 302161 320454
rect 305499 320514 305565 320517
rect 305678 320514 305684 320516
rect 305499 320512 305684 320514
rect 305499 320456 305504 320512
rect 305560 320456 305684 320512
rect 305499 320454 305684 320456
rect 305499 320451 305565 320454
rect 305678 320452 305684 320454
rect 305748 320452 305754 320516
rect 307618 320378 307678 320587
rect 325006 320517 325066 320590
rect 326708 320648 326817 320650
rect 326708 320592 326756 320648
rect 326812 320592 326817 320648
rect 326708 320587 326817 320592
rect 327303 320650 327369 320653
rect 327574 320650 327580 320652
rect 327303 320648 327580 320650
rect 327303 320592 327308 320648
rect 327364 320592 327580 320648
rect 327303 320590 327580 320592
rect 327303 320587 327369 320590
rect 327574 320588 327580 320590
rect 327644 320588 327650 320652
rect 327717 320650 327783 320653
rect 335310 320650 335370 320726
rect 388161 320723 388227 320726
rect 327717 320648 335370 320650
rect 327717 320592 327722 320648
rect 327778 320592 335370 320648
rect 327717 320590 335370 320592
rect 327717 320587 327783 320590
rect 312302 320452 312308 320516
rect 312372 320514 312378 320516
rect 312583 320514 312649 320517
rect 312372 320512 312649 320514
rect 312372 320456 312588 320512
rect 312644 320456 312649 320512
rect 312372 320454 312649 320456
rect 312372 320452 312378 320454
rect 312583 320451 312649 320454
rect 313503 320514 313569 320517
rect 313958 320514 313964 320516
rect 313503 320512 313964 320514
rect 313503 320456 313508 320512
rect 313564 320456 313964 320512
rect 313503 320454 313964 320456
rect 313503 320451 313569 320454
rect 313958 320452 313964 320454
rect 314028 320452 314034 320516
rect 318926 320452 318932 320516
rect 318996 320514 319002 320516
rect 319667 320514 319733 320517
rect 319846 320514 319852 320516
rect 318996 320512 319852 320514
rect 318996 320456 319672 320512
rect 319728 320456 319852 320512
rect 318996 320454 319852 320456
rect 318996 320452 319002 320454
rect 319667 320451 319733 320454
rect 319846 320452 319852 320454
rect 319916 320452 319922 320516
rect 322979 320514 323045 320517
rect 323158 320514 323164 320516
rect 322979 320512 323164 320514
rect 322979 320456 322984 320512
rect 323040 320456 323164 320512
rect 322979 320454 323164 320456
rect 322979 320451 323045 320454
rect 323158 320452 323164 320454
rect 323228 320452 323234 320516
rect 324359 320514 324425 320517
rect 324630 320514 324636 320516
rect 324359 320512 324636 320514
rect 324359 320456 324364 320512
rect 324420 320456 324636 320512
rect 324359 320454 324636 320456
rect 324359 320451 324425 320454
rect 324630 320452 324636 320454
rect 324700 320452 324706 320516
rect 325003 320512 325069 320517
rect 325003 320456 325008 320512
rect 325064 320456 325069 320512
rect 325003 320451 325069 320456
rect 326708 320514 326768 320587
rect 327717 320516 327783 320517
rect 326838 320514 326844 320516
rect 326708 320454 326844 320514
rect 326838 320452 326844 320454
rect 326908 320452 326914 320516
rect 327717 320514 327764 320516
rect 327672 320512 327764 320514
rect 327672 320456 327722 320512
rect 327672 320454 327764 320456
rect 327717 320452 327764 320454
rect 327828 320452 327834 320516
rect 328361 320514 328427 320517
rect 336825 320514 336891 320517
rect 337193 320514 337259 320517
rect 328361 320512 337259 320514
rect 328361 320456 328366 320512
rect 328422 320456 336830 320512
rect 336886 320456 337198 320512
rect 337254 320456 337259 320512
rect 328361 320454 337259 320456
rect 327717 320451 327783 320452
rect 328361 320451 328427 320454
rect 336825 320451 336891 320454
rect 337193 320451 337259 320454
rect 271137 320376 288634 320378
rect 271137 320320 271142 320376
rect 271198 320320 288634 320376
rect 271137 320318 288634 320320
rect 288758 320318 289554 320378
rect 289770 320344 291394 320378
rect 291518 320344 307678 320378
rect 289770 320318 307678 320344
rect 271137 320315 271203 320318
rect 217869 320242 217935 320245
rect 277853 320242 277919 320245
rect 217869 320240 277919 320242
rect 217869 320184 217874 320240
rect 217930 320184 277858 320240
rect 277914 320184 277919 320240
rect 217869 320182 277919 320184
rect 217869 320179 217935 320182
rect 277853 320179 277919 320182
rect 278221 320242 278287 320245
rect 284523 320242 284589 320245
rect 278221 320240 284589 320242
rect 278221 320184 278226 320240
rect 278282 320184 284528 320240
rect 284584 320184 284589 320240
rect 278221 320182 284589 320184
rect 278221 320179 278287 320182
rect 284523 320179 284589 320182
rect 284891 320240 284957 320245
rect 285443 320242 285509 320245
rect 284891 320184 284896 320240
rect 284952 320184 284957 320240
rect 284891 320179 284957 320184
rect 285262 320240 285509 320242
rect 285262 320184 285448 320240
rect 285504 320184 285509 320240
rect 285262 320182 285509 320184
rect 282867 320104 282933 320109
rect 282867 320048 282872 320104
rect 282928 320048 282933 320104
rect 282867 320043 282933 320048
rect 283327 320104 283393 320109
rect 283327 320048 283332 320104
rect 283388 320048 283393 320104
rect 283327 320043 283393 320048
rect 283603 320106 283669 320109
rect 283782 320106 283788 320108
rect 283603 320104 283788 320106
rect 283603 320048 283608 320104
rect 283664 320048 283788 320104
rect 283603 320046 283788 320048
rect 283603 320043 283669 320046
rect 283782 320044 283788 320046
rect 283852 320044 283858 320108
rect 284063 320106 284129 320109
rect 284020 320104 284129 320106
rect 284020 320048 284068 320104
rect 284124 320048 284129 320104
rect 284020 320043 284129 320048
rect 284518 320044 284524 320108
rect 284588 320106 284594 320108
rect 284894 320106 284954 320179
rect 284588 320046 284954 320106
rect 284588 320044 284594 320046
rect 281625 319970 281691 319973
rect 282870 319970 282930 320043
rect 281625 319968 282930 319970
rect 281625 319912 281630 319968
rect 281686 319912 282930 319968
rect 281625 319910 282930 319912
rect 283330 319970 283390 320043
rect 283598 319970 283604 319972
rect 283330 319910 283604 319970
rect 281625 319907 281691 319910
rect 283598 319908 283604 319910
rect 283668 319908 283674 319972
rect 283787 319934 283853 319939
rect 283787 319878 283792 319934
rect 283848 319878 283853 319934
rect 283787 319873 283853 319878
rect 282499 319832 282565 319837
rect 282499 319776 282504 319832
rect 282560 319776 282565 319832
rect 282499 319771 282565 319776
rect 215201 319698 215267 319701
rect 281809 319698 281875 319701
rect 282502 319698 282562 319771
rect 215201 319696 282562 319698
rect 215201 319640 215206 319696
rect 215262 319640 281814 319696
rect 281870 319640 282562 319696
rect 215201 319638 282562 319640
rect 283097 319698 283163 319701
rect 283790 319698 283850 319873
rect 284020 319701 284080 320043
rect 284334 319970 284340 319972
rect 284296 319939 284340 319970
rect 284247 319934 284340 319939
rect 284247 319878 284252 319934
rect 284308 319908 284340 319934
rect 284404 319908 284410 319972
rect 284308 319878 284356 319908
rect 284247 319876 284356 319878
rect 284247 319873 284313 319876
rect 285262 319834 285322 320182
rect 285443 320179 285509 320182
rect 286542 320180 286548 320244
rect 286612 320242 286618 320244
rect 286823 320242 286889 320245
rect 287283 320244 287349 320245
rect 287278 320242 287284 320244
rect 286612 320240 286889 320242
rect 286612 320184 286828 320240
rect 286884 320184 286889 320240
rect 286612 320182 286889 320184
rect 287192 320182 287284 320242
rect 286612 320180 286618 320182
rect 286823 320179 286889 320182
rect 287278 320180 287284 320182
rect 287348 320180 287354 320244
rect 288019 320242 288085 320245
rect 288382 320242 288388 320244
rect 288019 320240 288388 320242
rect 288019 320184 288024 320240
rect 288080 320184 288388 320240
rect 288019 320182 288388 320184
rect 287283 320179 287349 320180
rect 288019 320179 288085 320182
rect 288382 320180 288388 320182
rect 288452 320180 288458 320244
rect 288574 320242 288634 320318
rect 289770 320242 289830 320318
rect 291334 320284 291578 320318
rect 308254 320316 308260 320380
rect 308324 320378 308330 320380
rect 308719 320378 308785 320381
rect 308324 320376 308785 320378
rect 308324 320320 308724 320376
rect 308780 320320 308785 320376
rect 308324 320318 308785 320320
rect 308324 320316 308330 320318
rect 308719 320315 308785 320318
rect 309174 320316 309180 320380
rect 309244 320378 309250 320380
rect 309455 320378 309521 320381
rect 310278 320378 310284 320380
rect 309244 320376 310284 320378
rect 309244 320320 309460 320376
rect 309516 320320 310284 320376
rect 309244 320318 310284 320320
rect 309244 320316 309250 320318
rect 309455 320315 309521 320318
rect 310278 320316 310284 320318
rect 310348 320316 310354 320380
rect 310927 320378 310993 320381
rect 311198 320378 311204 320380
rect 310927 320376 311204 320378
rect 310927 320320 310932 320376
rect 310988 320320 311204 320376
rect 310927 320318 311204 320320
rect 310927 320315 310993 320318
rect 311198 320316 311204 320318
rect 311268 320316 311274 320380
rect 311479 320378 311545 320381
rect 323531 320380 323597 320381
rect 311479 320376 321570 320378
rect 311479 320320 311484 320376
rect 311540 320320 321570 320376
rect 311479 320318 321570 320320
rect 311479 320315 311545 320318
rect 290319 320242 290385 320245
rect 291142 320242 291148 320244
rect 288574 320182 289830 320242
rect 290046 320240 291148 320242
rect 290046 320184 290324 320240
rect 290380 320184 291148 320240
rect 290046 320182 291148 320184
rect 285627 320108 285693 320109
rect 285622 320106 285628 320108
rect 285536 320046 285628 320106
rect 285622 320044 285628 320046
rect 285692 320044 285698 320108
rect 286271 320106 286337 320109
rect 286915 320108 286981 320109
rect 286726 320106 286732 320108
rect 286271 320104 286732 320106
rect 286271 320048 286276 320104
rect 286332 320048 286732 320104
rect 286271 320046 286732 320048
rect 285627 320043 285693 320044
rect 286271 320043 286337 320046
rect 286726 320044 286732 320046
rect 286796 320044 286802 320108
rect 286910 320044 286916 320108
rect 286980 320106 286986 320108
rect 287191 320106 287257 320109
rect 286980 320046 287072 320106
rect 287191 320104 287300 320106
rect 287191 320048 287196 320104
rect 287252 320048 287300 320104
rect 286980 320044 286986 320046
rect 286915 320043 286981 320044
rect 287191 320043 287300 320048
rect 287467 320104 287533 320109
rect 287467 320048 287472 320104
rect 287528 320048 287533 320104
rect 287467 320043 287533 320048
rect 287646 320044 287652 320108
rect 287716 320106 287722 320108
rect 287835 320106 287901 320109
rect 288111 320106 288177 320109
rect 288479 320106 288545 320109
rect 287716 320104 287901 320106
rect 287716 320048 287840 320104
rect 287896 320048 287901 320104
rect 287716 320046 287901 320048
rect 287716 320044 287722 320046
rect 287835 320043 287901 320046
rect 287976 320104 288177 320106
rect 287976 320048 288116 320104
rect 288172 320048 288177 320104
rect 287976 320046 288177 320048
rect 286455 319936 286521 319939
rect 286455 319934 286564 319936
rect 286455 319878 286460 319934
rect 286516 319878 286564 319934
rect 286455 319873 286564 319878
rect 285581 319834 285647 319837
rect 285262 319832 285647 319834
rect 285262 319776 285586 319832
rect 285642 319776 285647 319832
rect 285262 319774 285647 319776
rect 285581 319771 285647 319774
rect 285765 319834 285831 319837
rect 286179 319834 286245 319837
rect 285765 319832 286245 319834
rect 285765 319776 285770 319832
rect 285826 319776 286184 319832
rect 286240 319776 286245 319832
rect 285765 319774 286245 319776
rect 285765 319771 285831 319774
rect 286179 319771 286245 319774
rect 283097 319696 283850 319698
rect 283097 319640 283102 319696
rect 283158 319640 283850 319696
rect 283097 319638 283850 319640
rect 284017 319696 284083 319701
rect 284017 319640 284022 319696
rect 284078 319640 284083 319696
rect 215201 319635 215267 319638
rect 281809 319635 281875 319638
rect 283097 319635 283163 319638
rect 284017 319635 284083 319640
rect 284293 319698 284359 319701
rect 285070 319698 285076 319700
rect 284293 319696 285076 319698
rect 284293 319640 284298 319696
rect 284354 319640 285076 319696
rect 284293 319638 285076 319640
rect 284293 319635 284359 319638
rect 285070 319636 285076 319638
rect 285140 319636 285146 319700
rect 286504 319698 286564 319873
rect 287240 319837 287300 320043
rect 287470 319970 287530 320043
rect 287976 319970 288036 320046
rect 288111 320043 288177 320046
rect 288344 320104 288545 320106
rect 288344 320048 288484 320104
rect 288540 320048 288545 320104
rect 288344 320046 288545 320048
rect 287470 319910 287668 319970
rect 287976 319910 288266 319970
rect 287237 319832 287303 319837
rect 287237 319776 287242 319832
rect 287298 319776 287303 319832
rect 287237 319771 287303 319776
rect 287608 319701 287668 319910
rect 287927 319834 287993 319837
rect 287927 319832 288036 319834
rect 287927 319776 287932 319832
rect 287988 319776 288036 319832
rect 287927 319771 288036 319776
rect 287976 319701 288036 319771
rect 286777 319698 286843 319701
rect 287421 319700 287487 319701
rect 287421 319698 287468 319700
rect 286504 319696 286843 319698
rect 286504 319640 286782 319696
rect 286838 319640 286843 319696
rect 286504 319638 286843 319640
rect 287376 319696 287468 319698
rect 287376 319640 287426 319696
rect 287376 319638 287468 319640
rect 286777 319635 286843 319638
rect 287421 319636 287468 319638
rect 287532 319636 287538 319700
rect 287605 319696 287671 319701
rect 287973 319700 288039 319701
rect 287973 319698 288020 319700
rect 287605 319640 287610 319696
rect 287666 319640 287671 319696
rect 287421 319635 287487 319636
rect 287605 319635 287671 319640
rect 287928 319696 288020 319698
rect 287928 319640 287978 319696
rect 287928 319638 288020 319640
rect 287973 319636 288020 319638
rect 288084 319636 288090 319700
rect 288206 319698 288266 319910
rect 288344 319834 288404 320046
rect 288479 320043 288545 320046
rect 288663 320106 288729 320109
rect 288934 320106 288940 320108
rect 288663 320104 288940 320106
rect 288663 320048 288668 320104
rect 288724 320048 288940 320104
rect 288663 320046 288940 320048
rect 288663 320043 288729 320046
rect 288934 320044 288940 320046
rect 289004 320044 289010 320108
rect 289215 320106 289281 320109
rect 289486 320106 289492 320108
rect 289172 320104 289492 320106
rect 289172 320048 289220 320104
rect 289276 320048 289492 320104
rect 289172 320046 289492 320048
rect 289172 320043 289281 320046
rect 289486 320044 289492 320046
rect 289556 320044 289562 320108
rect 289767 320104 289833 320109
rect 289767 320048 289772 320104
rect 289828 320048 289833 320104
rect 289767 320043 289833 320048
rect 288566 319908 288572 319972
rect 288636 319970 288642 319972
rect 288636 319939 289002 319970
rect 288636 319934 289005 319939
rect 288636 319910 288944 319934
rect 288636 319908 288642 319910
rect 288939 319878 288944 319910
rect 289000 319878 289005 319934
rect 288939 319873 289005 319878
rect 289172 319837 289232 320043
rect 289770 319970 289830 320043
rect 289678 319910 289830 319970
rect 288617 319834 288683 319837
rect 288344 319832 288683 319834
rect 288344 319776 288622 319832
rect 288678 319776 288683 319832
rect 288344 319774 288683 319776
rect 288617 319771 288683 319774
rect 289169 319832 289235 319837
rect 289169 319776 289174 319832
rect 289230 319776 289235 319832
rect 289169 319771 289235 319776
rect 288525 319698 288591 319701
rect 288206 319696 288591 319698
rect 288206 319640 288530 319696
rect 288586 319640 288591 319696
rect 288206 319638 288591 319640
rect 287973 319635 288039 319636
rect 288525 319635 288591 319638
rect 288750 319636 288756 319700
rect 288820 319698 288826 319700
rect 289678 319698 289738 319910
rect 289813 319834 289879 319837
rect 290046 319834 290106 320182
rect 290319 320179 290385 320182
rect 291142 320180 291148 320182
rect 291212 320180 291218 320244
rect 291975 320242 292041 320245
rect 292246 320242 292252 320244
rect 291975 320240 292252 320242
rect 291975 320184 291980 320240
rect 292036 320184 292252 320240
rect 291975 320182 292252 320184
rect 291975 320179 292041 320182
rect 292246 320180 292252 320182
rect 292316 320180 292322 320244
rect 292435 320240 292501 320245
rect 292435 320184 292440 320240
rect 292496 320184 292501 320240
rect 292435 320179 292501 320184
rect 292982 320180 292988 320244
rect 293052 320242 293058 320244
rect 293350 320242 293356 320244
rect 293052 320182 293356 320242
rect 293052 320180 293058 320182
rect 293350 320180 293356 320182
rect 293420 320242 293426 320244
rect 293723 320242 293789 320245
rect 293420 320240 293789 320242
rect 293420 320184 293728 320240
rect 293784 320184 293789 320240
rect 293420 320182 293789 320184
rect 293420 320180 293426 320182
rect 293723 320179 293789 320182
rect 294275 320242 294341 320245
rect 294643 320242 294709 320245
rect 295011 320244 295077 320245
rect 294822 320242 294828 320244
rect 294275 320240 294522 320242
rect 294275 320184 294280 320240
rect 294336 320184 294522 320240
rect 294275 320182 294522 320184
rect 294275 320179 294341 320182
rect 290411 320104 290477 320109
rect 290687 320106 290753 320109
rect 290411 320048 290416 320104
rect 290472 320048 290477 320104
rect 290411 320043 290477 320048
rect 290552 320104 290753 320106
rect 290552 320048 290692 320104
rect 290748 320048 290753 320104
rect 290552 320046 290753 320048
rect 290414 319970 290474 320043
rect 289813 319832 290106 319834
rect 289813 319776 289818 319832
rect 289874 319776 290106 319832
rect 289813 319774 290106 319776
rect 290322 319910 290474 319970
rect 290552 319970 290612 320046
rect 290687 320043 290753 320046
rect 290963 320104 291029 320109
rect 290963 320048 290968 320104
rect 291024 320048 291029 320104
rect 290963 320043 291029 320048
rect 291147 320104 291213 320109
rect 291147 320048 291152 320104
rect 291208 320048 291213 320104
rect 291147 320043 291213 320048
rect 291326 320044 291332 320108
rect 291396 320106 291402 320108
rect 291699 320106 291765 320109
rect 291396 320104 291765 320106
rect 291396 320048 291704 320104
rect 291760 320048 291765 320104
rect 291396 320046 291765 320048
rect 291396 320044 291402 320046
rect 291699 320043 291765 320046
rect 292062 320044 292068 320108
rect 292132 320106 292138 320108
rect 292438 320106 292498 320179
rect 292132 320046 292498 320106
rect 292132 320044 292138 320046
rect 292614 320044 292620 320108
rect 292684 320106 292690 320108
rect 292803 320106 292869 320109
rect 292684 320104 292869 320106
rect 292684 320048 292808 320104
rect 292864 320048 292869 320104
rect 292684 320046 292869 320048
rect 292684 320044 292690 320046
rect 292803 320043 292869 320046
rect 293079 320106 293145 320109
rect 293999 320106 294065 320109
rect 294462 320108 294522 320182
rect 294643 320240 294828 320242
rect 294643 320184 294648 320240
rect 294704 320184 294828 320240
rect 294643 320182 294828 320184
rect 294643 320179 294709 320182
rect 294822 320180 294828 320182
rect 294892 320180 294898 320244
rect 295006 320180 295012 320244
rect 295076 320242 295082 320244
rect 295076 320182 295168 320242
rect 295076 320180 295082 320182
rect 295742 320180 295748 320244
rect 295812 320242 295818 320244
rect 296023 320242 296089 320245
rect 295812 320240 296089 320242
rect 295812 320184 296028 320240
rect 296084 320184 296089 320240
rect 295812 320182 296089 320184
rect 295812 320180 295818 320182
rect 295011 320179 295077 320180
rect 296023 320179 296089 320182
rect 296294 320180 296300 320244
rect 296364 320242 296370 320244
rect 296483 320242 296549 320245
rect 296943 320242 297009 320245
rect 298691 320244 298757 320245
rect 298686 320242 298692 320244
rect 296364 320240 296549 320242
rect 296364 320184 296488 320240
rect 296544 320184 296549 320240
rect 296364 320182 296549 320184
rect 296364 320180 296370 320182
rect 296483 320179 296549 320182
rect 296670 320240 297009 320242
rect 296670 320184 296948 320240
rect 297004 320184 297009 320240
rect 296670 320182 297009 320184
rect 298600 320182 298692 320242
rect 294270 320106 294276 320108
rect 293079 320104 293188 320106
rect 293079 320048 293084 320104
rect 293140 320048 293188 320104
rect 293079 320043 293188 320048
rect 293999 320104 294276 320106
rect 293999 320048 294004 320104
rect 294060 320048 294276 320104
rect 293999 320046 294276 320048
rect 293999 320043 294065 320046
rect 294270 320044 294276 320046
rect 294340 320044 294346 320108
rect 294454 320044 294460 320108
rect 294524 320106 294530 320108
rect 295190 320106 295196 320108
rect 294524 320046 295196 320106
rect 294524 320044 294530 320046
rect 295190 320044 295196 320046
rect 295260 320044 295266 320108
rect 295374 320044 295380 320108
rect 295444 320106 295450 320108
rect 295839 320106 295905 320109
rect 295444 320104 295905 320106
rect 295444 320048 295844 320104
rect 295900 320048 295905 320104
rect 295444 320046 295905 320048
rect 295444 320044 295450 320046
rect 295839 320043 295905 320046
rect 296207 320106 296273 320109
rect 296478 320106 296484 320108
rect 296207 320104 296484 320106
rect 296207 320048 296212 320104
rect 296268 320048 296484 320104
rect 296207 320046 296484 320048
rect 296207 320043 296273 320046
rect 296478 320044 296484 320046
rect 296548 320044 296554 320108
rect 290774 319970 290780 319972
rect 290552 319910 290780 319970
rect 289813 319771 289879 319774
rect 288820 319638 289738 319698
rect 290322 319701 290382 319910
rect 290774 319908 290780 319910
rect 290844 319908 290850 319972
rect 290595 319834 290661 319837
rect 290774 319834 290780 319836
rect 290595 319832 290780 319834
rect 290595 319776 290600 319832
rect 290656 319776 290780 319832
rect 290595 319774 290780 319776
rect 290595 319771 290661 319774
rect 290774 319772 290780 319774
rect 290844 319772 290850 319836
rect 290322 319696 290431 319701
rect 290322 319640 290370 319696
rect 290426 319640 290431 319696
rect 290322 319638 290431 319640
rect 288820 319636 288826 319638
rect 290365 319635 290431 319638
rect 290733 319698 290799 319701
rect 290966 319698 291026 320043
rect 291150 319837 291210 320043
rect 292982 319908 292988 319972
rect 293052 319970 293058 319972
rect 293128 319970 293188 320043
rect 296670 319970 296730 320182
rect 296943 320179 297009 320182
rect 298686 320180 298692 320182
rect 298756 320180 298762 320244
rect 299151 320242 299217 320245
rect 300163 320244 300229 320245
rect 302739 320244 302805 320245
rect 299422 320242 299428 320244
rect 299151 320240 299428 320242
rect 299151 320184 299156 320240
rect 299212 320184 299428 320240
rect 299151 320182 299428 320184
rect 298691 320179 298757 320180
rect 299151 320179 299217 320182
rect 299422 320180 299428 320182
rect 299492 320180 299498 320244
rect 300158 320242 300164 320244
rect 300036 320182 300164 320242
rect 300228 320242 300234 320244
rect 302734 320242 302740 320244
rect 300158 320180 300164 320182
rect 300228 320182 302434 320242
rect 302648 320182 302740 320242
rect 300228 320180 300234 320182
rect 300163 320179 300229 320180
rect 296846 320044 296852 320108
rect 296916 320106 296922 320108
rect 297219 320106 297285 320109
rect 297587 320108 297653 320109
rect 297771 320108 297837 320109
rect 297582 320106 297588 320108
rect 296916 320104 297285 320106
rect 296916 320048 297224 320104
rect 297280 320048 297285 320104
rect 296916 320046 297285 320048
rect 297496 320046 297588 320106
rect 296916 320044 296922 320046
rect 297219 320043 297285 320046
rect 297582 320044 297588 320046
rect 297652 320044 297658 320108
rect 297766 320044 297772 320108
rect 297836 320106 297842 320108
rect 297836 320046 297928 320106
rect 297836 320044 297842 320046
rect 298134 320044 298140 320108
rect 298204 320106 298210 320108
rect 298415 320106 298481 320109
rect 299059 320108 299125 320109
rect 298870 320106 298876 320108
rect 298204 320104 298876 320106
rect 298204 320048 298420 320104
rect 298476 320048 298876 320104
rect 298204 320046 298876 320048
rect 298204 320044 298210 320046
rect 297587 320043 297653 320044
rect 297771 320043 297837 320044
rect 298415 320043 298481 320046
rect 298870 320044 298876 320046
rect 298940 320044 298946 320108
rect 299054 320044 299060 320108
rect 299124 320106 299130 320108
rect 299124 320046 299216 320106
rect 299427 320104 299493 320109
rect 299427 320048 299432 320104
rect 299488 320048 299493 320104
rect 299124 320044 299130 320046
rect 299059 320043 299125 320044
rect 299427 320043 299493 320048
rect 299790 320044 299796 320108
rect 299860 320106 299866 320108
rect 300071 320106 300137 320109
rect 299860 320104 300137 320106
rect 299860 320048 300076 320104
rect 300132 320048 300137 320104
rect 299860 320046 300137 320048
rect 299860 320044 299866 320046
rect 300071 320043 300137 320046
rect 300255 320106 300321 320109
rect 300899 320108 300965 320109
rect 300526 320106 300532 320108
rect 300255 320104 300532 320106
rect 300255 320048 300260 320104
rect 300316 320048 300532 320104
rect 300255 320046 300532 320048
rect 300255 320043 300321 320046
rect 300526 320044 300532 320046
rect 300596 320044 300602 320108
rect 300894 320106 300900 320108
rect 300808 320046 300900 320106
rect 300964 320106 300970 320108
rect 301998 320106 302004 320108
rect 300894 320044 300900 320046
rect 300964 320046 302004 320106
rect 300964 320044 300970 320046
rect 301998 320044 302004 320046
rect 302068 320044 302074 320108
rect 300899 320043 300965 320044
rect 293052 319910 293188 319970
rect 294232 319910 296730 319970
rect 293052 319908 293058 319910
rect 294232 319837 294292 319910
rect 298870 319908 298876 319972
rect 298940 319970 298946 319972
rect 299430 319970 299490 320043
rect 298940 319910 299490 319970
rect 302374 319970 302434 320182
rect 302734 320180 302740 320182
rect 302804 320180 302810 320244
rect 304758 320180 304764 320244
rect 304828 320242 304834 320244
rect 305131 320242 305197 320245
rect 304828 320240 305197 320242
rect 304828 320184 305136 320240
rect 305192 320184 305197 320240
rect 304828 320182 305197 320184
rect 304828 320180 304834 320182
rect 302739 320179 302805 320180
rect 305131 320179 305197 320182
rect 305494 320180 305500 320244
rect 305564 320242 305570 320244
rect 306235 320242 306301 320245
rect 305564 320240 306301 320242
rect 305564 320184 306240 320240
rect 306296 320184 306301 320240
rect 305564 320182 306301 320184
rect 305564 320180 305570 320182
rect 306235 320179 306301 320182
rect 306782 320180 306788 320244
rect 306852 320242 306858 320244
rect 307063 320242 307129 320245
rect 308443 320244 308509 320245
rect 308627 320244 308693 320245
rect 308438 320242 308444 320244
rect 306852 320240 307129 320242
rect 306852 320184 307068 320240
rect 307124 320184 307129 320240
rect 306852 320182 307129 320184
rect 308352 320182 308444 320242
rect 306852 320180 306858 320182
rect 307063 320179 307129 320182
rect 308438 320180 308444 320182
rect 308508 320180 308514 320244
rect 308622 320180 308628 320244
rect 308692 320242 308698 320244
rect 308692 320182 308784 320242
rect 308692 320180 308698 320182
rect 309358 320180 309364 320244
rect 309428 320242 309434 320244
rect 309639 320242 309705 320245
rect 309428 320240 309705 320242
rect 309428 320184 309644 320240
rect 309700 320184 309705 320240
rect 309428 320182 309705 320184
rect 309428 320180 309434 320182
rect 308443 320179 308509 320180
rect 308627 320179 308693 320180
rect 309639 320179 309705 320182
rect 312491 320242 312557 320245
rect 312670 320242 312676 320244
rect 312491 320240 312676 320242
rect 312491 320184 312496 320240
rect 312552 320184 312676 320240
rect 312491 320182 312676 320184
rect 312491 320179 312557 320182
rect 312670 320180 312676 320182
rect 312740 320180 312746 320244
rect 313774 320180 313780 320244
rect 313844 320242 313850 320244
rect 314147 320242 314213 320245
rect 313844 320240 314213 320242
rect 313844 320184 314152 320240
rect 314208 320184 314213 320240
rect 313844 320182 314213 320184
rect 313844 320180 313850 320182
rect 314147 320179 314213 320182
rect 314975 320242 315041 320245
rect 315614 320242 315620 320244
rect 314975 320240 315620 320242
rect 314975 320184 314980 320240
rect 315036 320184 315620 320240
rect 314975 320182 315620 320184
rect 314975 320179 315041 320182
rect 315614 320180 315620 320182
rect 315684 320180 315690 320244
rect 316350 320180 316356 320244
rect 316420 320242 316426 320244
rect 316907 320242 316973 320245
rect 316420 320240 316973 320242
rect 316420 320184 316912 320240
rect 316968 320184 316973 320240
rect 316420 320182 316973 320184
rect 316420 320180 316426 320182
rect 316907 320179 316973 320182
rect 319115 320242 319181 320245
rect 319851 320244 319917 320245
rect 320587 320244 320653 320245
rect 319662 320242 319668 320244
rect 319115 320240 319668 320242
rect 319115 320184 319120 320240
rect 319176 320184 319668 320240
rect 319115 320182 319668 320184
rect 319115 320179 319181 320182
rect 319662 320180 319668 320182
rect 319732 320180 319738 320244
rect 319846 320180 319852 320244
rect 319916 320242 319922 320244
rect 320582 320242 320588 320244
rect 319916 320182 320008 320242
rect 320496 320182 320588 320242
rect 319916 320180 319922 320182
rect 320582 320180 320588 320182
rect 320652 320180 320658 320244
rect 321510 320242 321570 320318
rect 322974 320316 322980 320380
rect 323044 320378 323050 320380
rect 323526 320378 323532 320380
rect 323044 320318 323532 320378
rect 323044 320316 323050 320318
rect 323526 320316 323532 320318
rect 323596 320316 323602 320380
rect 324262 320316 324268 320380
rect 324332 320378 324338 320380
rect 325182 320378 325188 320380
rect 324332 320318 325188 320378
rect 324332 320316 324338 320318
rect 325182 320316 325188 320318
rect 325252 320378 325258 320380
rect 325463 320378 325529 320381
rect 325252 320376 325529 320378
rect 325252 320320 325468 320376
rect 325524 320320 325529 320376
rect 325252 320318 325529 320320
rect 325252 320316 325258 320318
rect 323531 320315 323597 320316
rect 325463 320315 325529 320318
rect 326291 320378 326357 320381
rect 342253 320378 342319 320381
rect 326291 320376 342319 320378
rect 326291 320320 326296 320376
rect 326352 320320 342258 320376
rect 342314 320320 342319 320376
rect 326291 320318 342319 320320
rect 326291 320315 326357 320318
rect 342253 320315 342319 320318
rect 335445 320242 335511 320245
rect 335813 320242 335879 320245
rect 321510 320240 335879 320242
rect 321510 320184 335450 320240
rect 335506 320184 335818 320240
rect 335874 320184 335879 320240
rect 321510 320182 335879 320184
rect 319851 320179 319917 320180
rect 320587 320179 320653 320180
rect 335445 320179 335511 320182
rect 335813 320179 335879 320182
rect 302550 320044 302556 320108
rect 302620 320106 302626 320108
rect 302831 320106 302897 320109
rect 303659 320108 303725 320109
rect 303286 320106 303292 320108
rect 302620 320104 303292 320106
rect 302620 320048 302836 320104
rect 302892 320048 303292 320104
rect 302620 320046 303292 320048
rect 302620 320044 302626 320046
rect 302831 320043 302897 320046
rect 303286 320044 303292 320046
rect 303356 320044 303362 320108
rect 303654 320106 303660 320108
rect 303568 320046 303660 320106
rect 303654 320044 303660 320046
rect 303724 320044 303730 320108
rect 305126 320044 305132 320108
rect 305196 320106 305202 320108
rect 305867 320106 305933 320109
rect 306971 320108 307037 320109
rect 307339 320108 307405 320109
rect 308075 320108 308141 320109
rect 306230 320106 306236 320108
rect 305196 320104 306236 320106
rect 305196 320048 305872 320104
rect 305928 320048 306236 320104
rect 305196 320046 306236 320048
rect 305196 320044 305202 320046
rect 303659 320043 303725 320044
rect 305867 320043 305933 320046
rect 306230 320044 306236 320046
rect 306300 320044 306306 320108
rect 306966 320106 306972 320108
rect 306880 320046 306972 320106
rect 306966 320044 306972 320046
rect 307036 320044 307042 320108
rect 307334 320106 307340 320108
rect 307248 320046 307340 320106
rect 307334 320044 307340 320046
rect 307404 320044 307410 320108
rect 308070 320106 308076 320108
rect 307984 320046 308076 320106
rect 308140 320106 308146 320108
rect 308990 320106 308996 320108
rect 308070 320044 308076 320046
rect 308140 320046 308996 320106
rect 308140 320044 308146 320046
rect 308990 320044 308996 320046
rect 309060 320044 309066 320108
rect 309542 320044 309548 320108
rect 309612 320106 309618 320108
rect 309823 320106 309889 320109
rect 309612 320104 309889 320106
rect 309612 320048 309828 320104
rect 309884 320048 309889 320104
rect 309612 320046 309889 320048
rect 309612 320044 309618 320046
rect 306971 320043 307037 320044
rect 307339 320043 307405 320044
rect 308075 320043 308141 320044
rect 309823 320043 309889 320046
rect 310094 320044 310100 320108
rect 310164 320106 310170 320108
rect 310283 320106 310349 320109
rect 310164 320104 310349 320106
rect 310164 320048 310288 320104
rect 310344 320048 310349 320104
rect 310164 320046 310349 320048
rect 310164 320044 310170 320046
rect 310283 320043 310349 320046
rect 310830 320044 310836 320108
rect 310900 320106 310906 320108
rect 311663 320106 311729 320109
rect 312123 320108 312189 320109
rect 312118 320106 312124 320108
rect 310900 320104 311729 320106
rect 310900 320048 311668 320104
rect 311724 320048 311729 320104
rect 310900 320046 311729 320048
rect 312032 320046 312124 320106
rect 310900 320044 310906 320046
rect 311663 320043 311729 320046
rect 312118 320044 312124 320046
rect 312188 320044 312194 320108
rect 312486 320044 312492 320108
rect 312556 320106 312562 320108
rect 312767 320106 312833 320109
rect 312556 320104 312833 320106
rect 312556 320048 312772 320104
rect 312828 320048 312833 320104
rect 312556 320046 312833 320048
rect 312556 320044 312562 320046
rect 312123 320043 312189 320044
rect 312767 320043 312833 320046
rect 313871 320106 313937 320109
rect 314142 320106 314148 320108
rect 313871 320104 314148 320106
rect 313871 320048 313876 320104
rect 313932 320048 314148 320104
rect 313871 320046 314148 320048
rect 313871 320043 313937 320046
rect 314142 320044 314148 320046
rect 314212 320044 314218 320108
rect 314694 320044 314700 320108
rect 314764 320106 314770 320108
rect 315527 320106 315593 320109
rect 314764 320104 315593 320106
rect 314764 320048 315532 320104
rect 315588 320048 315593 320104
rect 314764 320046 315593 320048
rect 314764 320044 314770 320046
rect 315527 320043 315593 320046
rect 316631 320106 316697 320109
rect 316902 320106 316908 320108
rect 316631 320104 316908 320106
rect 316631 320048 316636 320104
rect 316692 320048 316908 320104
rect 316631 320046 316908 320048
rect 316631 320043 316697 320046
rect 316902 320044 316908 320046
rect 316972 320044 316978 320108
rect 317638 320044 317644 320108
rect 317708 320106 317714 320108
rect 318287 320106 318353 320109
rect 317708 320104 318353 320106
rect 317708 320048 318292 320104
rect 318348 320048 318353 320104
rect 317708 320046 318353 320048
rect 317708 320044 317714 320046
rect 318287 320043 318353 320046
rect 318839 320106 318905 320109
rect 319483 320108 319549 320109
rect 320035 320108 320101 320109
rect 319294 320106 319300 320108
rect 318839 320104 319300 320106
rect 318839 320048 318844 320104
rect 318900 320048 319300 320104
rect 318839 320046 319300 320048
rect 318839 320043 318905 320046
rect 319294 320044 319300 320046
rect 319364 320044 319370 320108
rect 319478 320044 319484 320108
rect 319548 320106 319554 320108
rect 320030 320106 320036 320108
rect 319548 320046 319640 320106
rect 319944 320046 320036 320106
rect 319548 320044 319554 320046
rect 320030 320044 320036 320046
rect 320100 320044 320106 320108
rect 320495 320106 320561 320109
rect 321323 320108 321389 320109
rect 322795 320108 322861 320109
rect 320950 320106 320956 320108
rect 320495 320104 320956 320106
rect 320495 320048 320500 320104
rect 320556 320048 320956 320104
rect 320495 320046 320956 320048
rect 319483 320043 319549 320044
rect 320035 320043 320101 320044
rect 320495 320043 320561 320046
rect 320950 320044 320956 320046
rect 321020 320044 321026 320108
rect 321318 320106 321324 320108
rect 321232 320046 321324 320106
rect 321318 320044 321324 320046
rect 321388 320044 321394 320108
rect 322790 320106 322796 320108
rect 322704 320046 322796 320106
rect 322790 320044 322796 320046
rect 322860 320044 322866 320108
rect 323347 320106 323413 320109
rect 323526 320106 323532 320108
rect 323347 320104 323532 320106
rect 323347 320048 323352 320104
rect 323408 320048 323532 320104
rect 323347 320046 323532 320048
rect 321323 320043 321389 320044
rect 322795 320043 322861 320044
rect 323347 320043 323413 320046
rect 323526 320044 323532 320046
rect 323596 320044 323602 320108
rect 324175 320106 324241 320109
rect 324451 320108 324517 320109
rect 324446 320106 324452 320108
rect 324132 320104 324241 320106
rect 324132 320048 324180 320104
rect 324236 320048 324241 320104
rect 324132 320043 324241 320048
rect 324360 320046 324452 320106
rect 324446 320044 324452 320046
rect 324516 320044 324522 320108
rect 324911 320106 324977 320109
rect 325366 320106 325372 320108
rect 324911 320104 325372 320106
rect 324911 320048 324916 320104
rect 324972 320048 325372 320104
rect 324911 320046 325372 320048
rect 324451 320043 324517 320044
rect 324911 320043 324977 320046
rect 325366 320044 325372 320046
rect 325436 320044 325442 320108
rect 325555 320104 325621 320109
rect 326567 320106 326633 320109
rect 326935 320106 327001 320109
rect 327206 320106 327212 320108
rect 325555 320048 325560 320104
rect 325616 320048 325621 320104
rect 325555 320043 325621 320048
rect 325742 320046 326170 320106
rect 306046 319970 306052 319972
rect 302374 319910 306052 319970
rect 298940 319908 298946 319910
rect 306046 319908 306052 319910
rect 306116 319908 306122 319972
rect 324132 319970 324192 320043
rect 324998 319970 325004 319972
rect 324132 319910 325004 319970
rect 324998 319908 325004 319910
rect 325068 319908 325074 319972
rect 325366 319908 325372 319972
rect 325436 319970 325442 319972
rect 325558 319970 325618 320043
rect 325436 319910 325618 319970
rect 325436 319908 325442 319910
rect 291101 319832 291210 319837
rect 291101 319776 291106 319832
rect 291162 319776 291210 319832
rect 291101 319774 291210 319776
rect 292297 319834 292363 319837
rect 292527 319834 292593 319837
rect 292297 319832 292593 319834
rect 292297 319776 292302 319832
rect 292358 319776 292532 319832
rect 292588 319776 292593 319832
rect 292297 319774 292593 319776
rect 291101 319771 291167 319774
rect 292297 319771 292363 319774
rect 292527 319771 292593 319774
rect 292760 319774 293188 319834
rect 292760 319698 292820 319774
rect 290733 319696 291026 319698
rect 290733 319640 290738 319696
rect 290794 319640 291026 319696
rect 290733 319638 291026 319640
rect 291840 319638 292820 319698
rect 290733 319635 290799 319638
rect 211061 319562 211127 319565
rect 278313 319562 278379 319565
rect 291840 319562 291900 319638
rect 292573 319562 292639 319565
rect 211061 319560 258090 319562
rect 211061 319504 211066 319560
rect 211122 319504 258090 319560
rect 211061 319502 258090 319504
rect 211061 319499 211127 319502
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect 258030 319290 258090 319502
rect 278313 319560 291900 319562
rect 278313 319504 278318 319560
rect 278374 319504 291900 319560
rect 278313 319502 291900 319504
rect 291978 319560 292639 319562
rect 291978 319504 292578 319560
rect 292634 319504 292639 319560
rect 291978 319502 292639 319504
rect 293128 319562 293188 319774
rect 294229 319832 294295 319837
rect 294229 319776 294234 319832
rect 294290 319776 294295 319832
rect 294229 319771 294295 319776
rect 295190 319772 295196 319836
rect 295260 319834 295266 319836
rect 325742 319834 325802 320046
rect 295260 319774 325802 319834
rect 326110 319834 326170 320046
rect 326567 320104 326768 320106
rect 326567 320048 326572 320104
rect 326628 320048 326768 320104
rect 326567 320046 326768 320048
rect 326567 320043 326633 320046
rect 326708 319972 326768 320046
rect 326935 320104 327212 320106
rect 326935 320048 326940 320104
rect 326996 320048 327212 320104
rect 326935 320046 327212 320048
rect 326935 320043 327001 320046
rect 327206 320044 327212 320046
rect 327276 320044 327282 320108
rect 326654 319908 326660 319972
rect 326724 319910 326768 319972
rect 327533 319972 327599 319973
rect 327533 319970 327580 319972
rect 327488 319968 327580 319970
rect 327488 319912 327538 319968
rect 327488 319910 327580 319912
rect 326724 319908 326730 319910
rect 327533 319908 327580 319910
rect 327644 319908 327650 319972
rect 327717 319970 327783 319973
rect 333973 319970 334039 319973
rect 327717 319968 334039 319970
rect 327717 319912 327722 319968
rect 327778 319912 333978 319968
rect 334034 319912 334039 319968
rect 327717 319910 334039 319912
rect 327533 319907 327599 319908
rect 327717 319907 327783 319910
rect 333973 319907 334039 319910
rect 346761 319834 346827 319837
rect 326110 319832 346827 319834
rect 326110 319776 346766 319832
rect 346822 319776 346827 319832
rect 326110 319774 346827 319776
rect 295260 319772 295266 319774
rect 346761 319771 346827 319774
rect 294965 319698 295031 319701
rect 344001 319698 344067 319701
rect 294965 319696 325802 319698
rect 294965 319640 294970 319696
rect 295026 319664 325802 319696
rect 326110 319696 344067 319698
rect 326110 319664 344006 319696
rect 295026 319640 344006 319664
rect 344062 319640 344067 319696
rect 294965 319638 344067 319640
rect 294965 319635 295031 319638
rect 325742 319604 326170 319638
rect 344001 319635 344067 319638
rect 305177 319562 305243 319565
rect 305494 319562 305500 319564
rect 293128 319502 302250 319562
rect 278313 319499 278379 319502
rect 283649 319426 283715 319429
rect 283782 319426 283788 319428
rect 283649 319424 283788 319426
rect 283649 319368 283654 319424
rect 283710 319368 283788 319424
rect 283649 319366 283788 319368
rect 283649 319363 283715 319366
rect 283782 319364 283788 319366
rect 283852 319364 283858 319428
rect 284017 319426 284083 319429
rect 291978 319426 292038 319502
rect 292573 319499 292639 319502
rect 284017 319424 292038 319426
rect 284017 319368 284022 319424
rect 284078 319368 292038 319424
rect 284017 319366 292038 319368
rect 292113 319426 292179 319429
rect 293033 319426 293099 319429
rect 292113 319424 293099 319426
rect 292113 319368 292118 319424
rect 292174 319368 293038 319424
rect 293094 319368 293099 319424
rect 292113 319366 293099 319368
rect 284017 319363 284083 319366
rect 292113 319363 292179 319366
rect 293033 319363 293099 319366
rect 294505 319426 294571 319429
rect 294822 319426 294828 319428
rect 294505 319424 294828 319426
rect 294505 319368 294510 319424
rect 294566 319368 294828 319424
rect 294505 319366 294828 319368
rect 294505 319363 294571 319366
rect 294822 319364 294828 319366
rect 294892 319364 294898 319428
rect 295558 319364 295564 319428
rect 295628 319426 295634 319428
rect 295793 319426 295859 319429
rect 295628 319424 295859 319426
rect 295628 319368 295798 319424
rect 295854 319368 295859 319424
rect 295628 319366 295859 319368
rect 295628 319364 295634 319366
rect 295793 319363 295859 319366
rect 297725 319426 297791 319429
rect 297950 319426 297956 319428
rect 297725 319424 297956 319426
rect 297725 319368 297730 319424
rect 297786 319368 297956 319424
rect 297725 319366 297956 319368
rect 297725 319363 297791 319366
rect 297950 319364 297956 319366
rect 298020 319364 298026 319428
rect 299933 319426 299999 319429
rect 300485 319428 300551 319429
rect 300158 319426 300164 319428
rect 299933 319424 300164 319426
rect 299933 319368 299938 319424
rect 299994 319368 300164 319424
rect 299933 319366 300164 319368
rect 299933 319363 299999 319366
rect 300158 319364 300164 319366
rect 300228 319364 300234 319428
rect 300485 319426 300532 319428
rect 300440 319424 300532 319426
rect 300440 319368 300490 319424
rect 300440 319366 300532 319368
rect 300485 319364 300532 319366
rect 300596 319364 300602 319428
rect 301497 319426 301563 319429
rect 301630 319426 301636 319428
rect 301497 319424 301636 319426
rect 301497 319368 301502 319424
rect 301558 319368 301636 319424
rect 301497 319366 301636 319368
rect 300485 319363 300551 319364
rect 301497 319363 301563 319366
rect 301630 319364 301636 319366
rect 301700 319364 301706 319428
rect 302190 319426 302250 319502
rect 305177 319560 305500 319562
rect 305177 319504 305182 319560
rect 305238 319504 305500 319560
rect 305177 319502 305500 319504
rect 305177 319499 305243 319502
rect 305494 319500 305500 319502
rect 305564 319500 305570 319564
rect 305729 319562 305795 319565
rect 306097 319564 306163 319565
rect 305862 319562 305868 319564
rect 305729 319560 305868 319562
rect 305729 319504 305734 319560
rect 305790 319504 305868 319560
rect 305729 319502 305868 319504
rect 305729 319499 305795 319502
rect 305862 319500 305868 319502
rect 305932 319500 305938 319564
rect 306046 319500 306052 319564
rect 306116 319562 306163 319564
rect 306741 319564 306807 319565
rect 307937 319564 308003 319565
rect 306741 319562 306788 319564
rect 306116 319560 306208 319562
rect 306158 319504 306208 319560
rect 306116 319502 306208 319504
rect 306696 319560 306788 319562
rect 306696 319504 306746 319560
rect 306696 319502 306788 319504
rect 306116 319500 306163 319502
rect 306097 319499 306163 319500
rect 306741 319500 306788 319502
rect 306852 319500 306858 319564
rect 307886 319500 307892 319564
rect 307956 319562 308003 319564
rect 308121 319562 308187 319565
rect 308438 319562 308444 319564
rect 307956 319560 308048 319562
rect 307998 319504 308048 319560
rect 307956 319502 308048 319504
rect 308121 319560 308444 319562
rect 308121 319504 308126 319560
rect 308182 319504 308444 319560
rect 308121 319502 308444 319504
rect 307956 319500 308003 319502
rect 306741 319499 306807 319500
rect 307937 319499 308003 319500
rect 308121 319499 308187 319502
rect 308438 319500 308444 319502
rect 308508 319500 308514 319564
rect 309225 319562 309291 319565
rect 309358 319562 309364 319564
rect 309225 319560 309364 319562
rect 309225 319504 309230 319560
rect 309286 319504 309364 319560
rect 309225 319502 309364 319504
rect 309225 319499 309291 319502
rect 309358 319500 309364 319502
rect 309428 319500 309434 319564
rect 309542 319500 309548 319564
rect 309612 319562 309618 319564
rect 309777 319562 309843 319565
rect 314009 319564 314075 319565
rect 309612 319560 309843 319562
rect 309612 319504 309782 319560
rect 309838 319504 309843 319560
rect 309612 319502 309843 319504
rect 309612 319500 309618 319502
rect 309777 319499 309843 319502
rect 313958 319500 313964 319564
rect 314028 319562 314075 319564
rect 317137 319562 317203 319565
rect 320633 319564 320699 319565
rect 317270 319562 317276 319564
rect 314028 319560 314120 319562
rect 314070 319504 314120 319560
rect 314028 319502 314120 319504
rect 317137 319560 317276 319562
rect 317137 319504 317142 319560
rect 317198 319504 317276 319560
rect 317137 319502 317276 319504
rect 314028 319500 314075 319502
rect 314009 319499 314075 319500
rect 317137 319499 317203 319502
rect 317270 319500 317276 319502
rect 317340 319500 317346 319564
rect 320582 319500 320588 319564
rect 320652 319562 320699 319564
rect 323485 319564 323551 319565
rect 323761 319564 323827 319565
rect 320652 319560 320744 319562
rect 320694 319504 320744 319560
rect 320652 319502 320744 319504
rect 323485 319560 323532 319564
rect 323596 319562 323602 319564
rect 323485 319504 323490 319560
rect 320652 319500 320699 319502
rect 320633 319499 320699 319500
rect 323485 319500 323532 319504
rect 323596 319502 323642 319562
rect 323596 319500 323602 319502
rect 323710 319500 323716 319564
rect 323780 319562 323827 319564
rect 325325 319564 325391 319565
rect 326613 319564 326679 319565
rect 325325 319562 325372 319564
rect 323780 319560 323872 319562
rect 323822 319504 323872 319560
rect 323780 319502 323872 319504
rect 325280 319560 325372 319562
rect 325280 319504 325330 319560
rect 325280 319502 325372 319504
rect 323780 319500 323827 319502
rect 323485 319499 323551 319500
rect 323761 319499 323827 319500
rect 325325 319500 325372 319502
rect 325436 319500 325442 319564
rect 326613 319562 326660 319564
rect 326568 319560 326660 319562
rect 326568 319504 326618 319560
rect 326568 319502 326660 319504
rect 326613 319500 326660 319502
rect 326724 319500 326730 319564
rect 326981 319562 327047 319565
rect 327441 319564 327507 319565
rect 327206 319562 327212 319564
rect 326981 319560 327212 319562
rect 326981 319504 326986 319560
rect 327042 319504 327212 319560
rect 326981 319502 327212 319504
rect 325325 319499 325391 319500
rect 326613 319499 326679 319500
rect 326981 319499 327047 319502
rect 327206 319500 327212 319502
rect 327276 319500 327282 319564
rect 327390 319500 327396 319564
rect 327460 319562 327507 319564
rect 327460 319560 327552 319562
rect 327502 319504 327552 319560
rect 327460 319502 327552 319504
rect 327460 319500 327507 319502
rect 327441 319499 327507 319500
rect 306649 319426 306715 319429
rect 307293 319428 307359 319429
rect 307293 319426 307340 319428
rect 302190 319424 306715 319426
rect 302190 319368 306654 319424
rect 306710 319368 306715 319424
rect 302190 319366 306715 319368
rect 307248 319424 307340 319426
rect 307248 319368 307298 319424
rect 307248 319366 307340 319368
rect 306649 319363 306715 319366
rect 307293 319364 307340 319366
rect 307404 319364 307410 319428
rect 307937 319426 308003 319429
rect 309685 319428 309751 319429
rect 308622 319426 308628 319428
rect 307937 319424 308628 319426
rect 307937 319368 307942 319424
rect 307998 319368 308628 319424
rect 307937 319366 308628 319368
rect 307293 319363 307359 319364
rect 307937 319363 308003 319366
rect 308622 319364 308628 319366
rect 308692 319364 308698 319428
rect 309685 319424 309732 319428
rect 309796 319426 309802 319428
rect 310973 319426 311039 319429
rect 312261 319428 312327 319429
rect 311198 319426 311204 319428
rect 309685 319368 309690 319424
rect 309685 319364 309732 319368
rect 309796 319366 309842 319426
rect 310973 319424 311204 319426
rect 310973 319368 310978 319424
rect 311034 319368 311204 319424
rect 310973 319366 311204 319368
rect 309796 319364 309802 319366
rect 309685 319363 309751 319364
rect 310973 319363 311039 319366
rect 311198 319364 311204 319366
rect 311268 319364 311274 319428
rect 312261 319426 312308 319428
rect 312216 319424 312308 319426
rect 312216 319368 312266 319424
rect 312216 319366 312308 319368
rect 312261 319364 312308 319366
rect 312372 319364 312378 319428
rect 313590 319364 313596 319428
rect 313660 319426 313666 319428
rect 314193 319426 314259 319429
rect 313660 319424 314259 319426
rect 313660 319368 314198 319424
rect 314254 319368 314259 319424
rect 313660 319366 314259 319368
rect 313660 319364 313666 319366
rect 312261 319363 312327 319364
rect 314193 319363 314259 319366
rect 318977 319426 319043 319429
rect 327717 319426 327783 319429
rect 318977 319424 327783 319426
rect 318977 319368 318982 319424
rect 319038 319368 327722 319424
rect 327778 319368 327783 319424
rect 318977 319366 327783 319368
rect 318977 319363 319043 319366
rect 327717 319363 327783 319366
rect 272885 319290 272951 319293
rect 282913 319290 282979 319293
rect 258030 319288 282979 319290
rect 258030 319232 272890 319288
rect 272946 319232 282918 319288
rect 282974 319232 282979 319288
rect 258030 319230 282979 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 272885 319227 272951 319230
rect 282913 319227 282979 319230
rect 283414 319228 283420 319292
rect 283484 319290 283490 319292
rect 283966 319290 283972 319292
rect 283484 319230 283972 319290
rect 283484 319228 283490 319230
rect 283966 319228 283972 319230
rect 284036 319228 284042 319292
rect 284477 319290 284543 319293
rect 285622 319290 285628 319292
rect 284477 319288 285628 319290
rect 284477 319232 284482 319288
rect 284538 319232 285628 319288
rect 284477 319230 285628 319232
rect 284477 319227 284543 319230
rect 285622 319228 285628 319230
rect 285692 319228 285698 319292
rect 286910 319228 286916 319292
rect 286980 319290 286986 319292
rect 287053 319290 287119 319293
rect 286980 319288 287119 319290
rect 286980 319232 287058 319288
rect 287114 319232 287119 319288
rect 286980 319230 287119 319232
rect 286980 319228 286986 319230
rect 287053 319227 287119 319230
rect 288065 319290 288131 319293
rect 288382 319290 288388 319292
rect 288065 319288 288388 319290
rect 288065 319232 288070 319288
rect 288126 319232 288388 319288
rect 288065 319230 288388 319232
rect 288065 319227 288131 319230
rect 288382 319228 288388 319230
rect 288452 319228 288458 319292
rect 288566 319228 288572 319292
rect 288636 319290 288642 319292
rect 288893 319290 288959 319293
rect 288636 319288 288959 319290
rect 288636 319232 288898 319288
rect 288954 319232 288959 319288
rect 288636 319230 288959 319232
rect 288636 319228 288642 319230
rect 288893 319227 288959 319230
rect 289077 319290 289143 319293
rect 292665 319292 292731 319293
rect 292614 319290 292620 319292
rect 289077 319288 292452 319290
rect 289077 319232 289082 319288
rect 289138 319232 292452 319288
rect 289077 319230 292452 319232
rect 292574 319230 292620 319290
rect 292684 319288 292731 319292
rect 292726 319232 292731 319288
rect 289077 319227 289143 319230
rect 287237 319154 287303 319157
rect 273210 319152 290842 319154
rect 273210 319096 287242 319152
rect 287298 319096 290842 319152
rect 273210 319094 290842 319096
rect 206921 318882 206987 318885
rect 273210 318882 273270 319094
rect 287237 319091 287303 319094
rect 278405 319018 278471 319021
rect 283230 319018 283236 319020
rect 278405 319016 283236 319018
rect 278405 318960 278410 319016
rect 278466 318960 283236 319016
rect 278405 318958 283236 318960
rect 278405 318955 278471 318958
rect 283230 318956 283236 318958
rect 283300 318956 283306 319020
rect 283598 318956 283604 319020
rect 283668 319018 283674 319020
rect 283833 319018 283899 319021
rect 284753 319020 284819 319021
rect 284702 319018 284708 319020
rect 283668 319016 283899 319018
rect 283668 318960 283838 319016
rect 283894 318960 283899 319016
rect 283668 318958 283899 318960
rect 284662 318958 284708 319018
rect 284772 319016 284819 319020
rect 284814 318960 284819 319016
rect 283668 318956 283674 318958
rect 283833 318955 283899 318958
rect 284702 318956 284708 318958
rect 284772 318956 284819 318960
rect 284886 318956 284892 319020
rect 284956 319018 284962 319020
rect 285029 319018 285095 319021
rect 287237 319020 287303 319021
rect 287237 319018 287284 319020
rect 284956 319016 285095 319018
rect 284956 318960 285034 319016
rect 285090 318960 285095 319016
rect 284956 318958 285095 318960
rect 287192 319016 287284 319018
rect 287192 318960 287242 319016
rect 287192 318958 287284 318960
rect 284956 318956 284962 318958
rect 284753 318955 284819 318956
rect 285029 318955 285095 318958
rect 287237 318956 287284 318958
rect 287348 318956 287354 319020
rect 288934 318956 288940 319020
rect 289004 319018 289010 319020
rect 289721 319018 289787 319021
rect 289004 319016 289787 319018
rect 289004 318960 289726 319016
rect 289782 318960 289787 319016
rect 289004 318958 289787 318960
rect 289004 318956 289010 318958
rect 287237 318955 287303 318956
rect 289721 318955 289787 318958
rect 206921 318880 273270 318882
rect 206921 318824 206926 318880
rect 206982 318824 273270 318880
rect 206921 318822 273270 318824
rect 277301 318882 277367 318885
rect 278313 318882 278379 318885
rect 277301 318880 278379 318882
rect 277301 318824 277306 318880
rect 277362 318824 278318 318880
rect 278374 318824 278379 318880
rect 277301 318822 278379 318824
rect 206921 318819 206987 318822
rect 277301 318819 277367 318822
rect 278313 318819 278379 318822
rect 279693 318882 279759 318885
rect 290590 318882 290596 318884
rect 279693 318880 290596 318882
rect 279693 318824 279698 318880
rect 279754 318824 290596 318880
rect 279693 318822 290596 318824
rect 279693 318819 279759 318822
rect 290590 318820 290596 318822
rect 290660 318820 290666 318884
rect 290782 318882 290842 319094
rect 291142 319092 291148 319156
rect 291212 319154 291218 319156
rect 292246 319154 292252 319156
rect 291212 319094 292252 319154
rect 291212 319092 291218 319094
rect 292246 319092 292252 319094
rect 292316 319092 292322 319156
rect 292392 319154 292452 319230
rect 292614 319228 292620 319230
rect 292684 319228 292731 319232
rect 292665 319227 292731 319228
rect 292941 319292 293007 319293
rect 292941 319288 292988 319292
rect 293052 319290 293058 319292
rect 294229 319290 294295 319293
rect 295006 319290 295012 319292
rect 292941 319232 292946 319288
rect 292941 319228 292988 319232
rect 293052 319230 293098 319290
rect 294229 319288 295012 319290
rect 294229 319232 294234 319288
rect 294290 319232 295012 319288
rect 294229 319230 295012 319232
rect 293052 319228 293058 319230
rect 292941 319227 293007 319228
rect 294229 319227 294295 319230
rect 295006 319228 295012 319230
rect 295076 319228 295082 319292
rect 295374 319228 295380 319292
rect 295444 319290 295450 319292
rect 296069 319290 296135 319293
rect 295444 319288 296135 319290
rect 295444 319232 296074 319288
rect 296130 319232 296135 319288
rect 295444 319230 296135 319232
rect 295444 319228 295450 319230
rect 296069 319227 296135 319230
rect 296713 319290 296779 319293
rect 296897 319290 296963 319293
rect 296713 319288 296963 319290
rect 296713 319232 296718 319288
rect 296774 319232 296902 319288
rect 296958 319232 296963 319288
rect 296713 319230 296963 319232
rect 296713 319227 296779 319230
rect 296897 319227 296963 319230
rect 297449 319290 297515 319293
rect 342529 319290 342595 319293
rect 297449 319288 342595 319290
rect 297449 319232 297454 319288
rect 297510 319232 342534 319288
rect 342590 319232 342595 319288
rect 297449 319230 342595 319232
rect 297449 319227 297515 319230
rect 342529 319227 342595 319230
rect 346945 319154 347011 319157
rect 292392 319152 347011 319154
rect 292392 319096 346950 319152
rect 347006 319096 347011 319152
rect 292392 319094 347011 319096
rect 346945 319091 347011 319094
rect 291745 319018 291811 319021
rect 292481 319018 292547 319021
rect 291745 319016 292547 319018
rect 291745 318960 291750 319016
rect 291806 318960 292486 319016
rect 292542 318960 292547 319016
rect 291745 318958 292547 318960
rect 291745 318955 291811 318958
rect 292481 318955 292547 318958
rect 292665 319018 292731 319021
rect 293677 319018 293743 319021
rect 295701 319020 295767 319021
rect 297357 319020 297423 319021
rect 295701 319018 295748 319020
rect 292665 319016 293743 319018
rect 292665 318960 292670 319016
rect 292726 318960 293682 319016
rect 293738 318960 293743 319016
rect 292665 318958 293743 318960
rect 295656 319016 295748 319018
rect 295656 318960 295706 319016
rect 295656 318958 295748 318960
rect 292665 318955 292731 318958
rect 293677 318955 293743 318958
rect 295701 318956 295748 318958
rect 295812 318956 295818 319020
rect 297357 319018 297404 319020
rect 297312 319016 297404 319018
rect 297312 318960 297362 319016
rect 297312 318958 297404 318960
rect 297357 318956 297404 318958
rect 297468 318956 297474 319020
rect 297541 319016 297607 319021
rect 297541 318960 297546 319016
rect 297602 318960 297607 319016
rect 295701 318955 295767 318956
rect 297357 318955 297423 318956
rect 297541 318955 297607 318960
rect 297725 319020 297791 319021
rect 298737 319020 298803 319021
rect 297725 319016 297772 319020
rect 297836 319018 297842 319020
rect 298686 319018 298692 319020
rect 297725 318960 297730 319016
rect 297725 318956 297772 318960
rect 297836 318958 297882 319018
rect 298610 318958 298692 319018
rect 298756 319018 298803 319020
rect 299381 319018 299447 319021
rect 298756 319016 299447 319018
rect 298798 318960 299386 319016
rect 299442 318960 299447 319016
rect 297836 318956 297842 318958
rect 298686 318956 298692 318958
rect 298756 318958 299447 318960
rect 298756 318956 298803 318958
rect 297725 318955 297791 318956
rect 298737 318955 298803 318956
rect 299381 318955 299447 318958
rect 300209 319018 300275 319021
rect 300342 319018 300348 319020
rect 300209 319016 300348 319018
rect 300209 318960 300214 319016
rect 300270 318960 300348 319016
rect 300209 318958 300348 318960
rect 300209 318955 300275 318958
rect 300342 318956 300348 318958
rect 300412 318956 300418 319020
rect 301681 319018 301747 319021
rect 304758 319018 304764 319020
rect 301681 319016 304764 319018
rect 301681 318960 301686 319016
rect 301742 318960 304764 319016
rect 301681 318958 304764 318960
rect 301681 318955 301747 318958
rect 304758 318956 304764 318958
rect 304828 318956 304834 319020
rect 305545 319018 305611 319021
rect 308213 319020 308279 319021
rect 312077 319020 312143 319021
rect 305678 319018 305684 319020
rect 305545 319016 305684 319018
rect 305545 318960 305550 319016
rect 305606 318960 305684 319016
rect 305545 318958 305684 318960
rect 305545 318955 305611 318958
rect 305678 318956 305684 318958
rect 305748 318956 305754 319020
rect 308213 319018 308260 319020
rect 308168 319016 308260 319018
rect 308168 318960 308218 319016
rect 308168 318958 308260 318960
rect 308213 318956 308260 318958
rect 308324 318956 308330 319020
rect 312077 319018 312124 319020
rect 312032 319016 312124 319018
rect 312032 318960 312082 319016
rect 312032 318958 312124 318960
rect 312077 318956 312124 318958
rect 312188 318956 312194 319020
rect 319478 318956 319484 319020
rect 319548 319018 319554 319020
rect 319621 319018 319687 319021
rect 319548 319016 319687 319018
rect 319548 318960 319626 319016
rect 319682 318960 319687 319016
rect 319548 318958 319687 318960
rect 319548 318956 319554 318958
rect 308213 318955 308279 318956
rect 312077 318955 312143 318956
rect 319621 318955 319687 318958
rect 319846 318956 319852 319020
rect 319916 319018 319922 319020
rect 319989 319018 320055 319021
rect 319916 319016 320055 319018
rect 319916 318960 319994 319016
rect 320050 318960 320055 319016
rect 319916 318958 320055 318960
rect 319916 318956 319922 318958
rect 319989 318955 320055 318958
rect 324446 318956 324452 319020
rect 324516 319018 324522 319020
rect 324589 319018 324655 319021
rect 324516 319016 324655 319018
rect 324516 318960 324594 319016
rect 324650 318960 324655 319016
rect 324516 318958 324655 318960
rect 324516 318956 324522 318958
rect 324589 318955 324655 318958
rect 324998 318956 325004 319020
rect 325068 319018 325074 319020
rect 328361 319018 328427 319021
rect 325068 319016 328427 319018
rect 325068 318960 328366 319016
rect 328422 318960 328427 319016
rect 325068 318958 328427 318960
rect 325068 318956 325074 318958
rect 328361 318955 328427 318958
rect 295190 318882 295196 318884
rect 290782 318822 295196 318882
rect 295190 318820 295196 318822
rect 295260 318820 295266 318884
rect 296897 318882 296963 318885
rect 297544 318882 297604 318955
rect 296897 318880 297604 318882
rect 296897 318824 296902 318880
rect 296958 318824 297604 318880
rect 296897 318822 297604 318824
rect 296897 318819 296963 318822
rect 298502 318820 298508 318884
rect 298572 318882 298578 318884
rect 299657 318882 299723 318885
rect 298572 318880 299723 318882
rect 298572 318824 299662 318880
rect 299718 318824 299723 318880
rect 298572 318822 299723 318824
rect 298572 318820 298578 318822
rect 299657 318819 299723 318822
rect 299790 318820 299796 318884
rect 299860 318882 299866 318884
rect 300117 318882 300183 318885
rect 299860 318880 300183 318882
rect 299860 318824 300122 318880
rect 300178 318824 300183 318880
rect 299860 318822 300183 318824
rect 299860 318820 299866 318822
rect 300117 318819 300183 318822
rect 307886 318820 307892 318884
rect 307956 318882 307962 318884
rect 309685 318882 309751 318885
rect 307956 318880 309751 318882
rect 307956 318824 309690 318880
rect 309746 318824 309751 318880
rect 307956 318822 309751 318824
rect 307956 318820 307962 318822
rect 309685 318819 309751 318822
rect 319713 318882 319779 318885
rect 320030 318882 320036 318884
rect 319713 318880 320036 318882
rect 319713 318824 319718 318880
rect 319774 318824 320036 318880
rect 319713 318822 320036 318824
rect 319713 318819 319779 318822
rect 320030 318820 320036 318822
rect 320100 318820 320106 318884
rect 324497 318882 324563 318885
rect 324630 318882 324636 318884
rect 324497 318880 324636 318882
rect 324497 318824 324502 318880
rect 324558 318824 324636 318880
rect 324497 318822 324636 318824
rect 324497 318819 324563 318822
rect 324630 318820 324636 318822
rect 324700 318820 324706 318884
rect 324814 318820 324820 318884
rect 324884 318882 324890 318884
rect 325049 318882 325115 318885
rect 324884 318880 325115 318882
rect 324884 318824 325054 318880
rect 325110 318824 325115 318880
rect 324884 318822 325115 318824
rect 324884 318820 324890 318822
rect 325049 318819 325115 318822
rect 325182 318820 325188 318884
rect 325252 318882 325258 318884
rect 328494 318882 328500 318884
rect 325252 318822 328500 318882
rect 325252 318820 325258 318822
rect 328494 318820 328500 318822
rect 328564 318820 328570 318884
rect 225873 318746 225939 318749
rect 283414 318746 283420 318748
rect 225873 318744 283420 318746
rect 225873 318688 225878 318744
rect 225934 318688 283420 318744
rect 225873 318686 283420 318688
rect 225873 318683 225939 318686
rect 283414 318684 283420 318686
rect 283484 318684 283490 318748
rect 286501 318746 286567 318749
rect 287830 318746 287836 318748
rect 286501 318744 287836 318746
rect 286501 318688 286506 318744
rect 286562 318688 287836 318744
rect 286501 318686 287836 318688
rect 286501 318683 286567 318686
rect 287830 318684 287836 318686
rect 287900 318684 287906 318748
rect 288341 318746 288407 318749
rect 294597 318748 294663 318749
rect 294597 318746 294644 318748
rect 288341 318744 293004 318746
rect 288341 318688 288346 318744
rect 288402 318688 293004 318744
rect 288341 318686 293004 318688
rect 294552 318744 294644 318746
rect 294552 318688 294602 318744
rect 294552 318686 294644 318688
rect 288341 318683 288407 318686
rect 230197 318610 230263 318613
rect 279601 318610 279667 318613
rect 289077 318610 289143 318613
rect 292798 318610 292804 318612
rect 230197 318608 273270 318610
rect 230197 318552 230202 318608
rect 230258 318552 273270 318608
rect 230197 318550 273270 318552
rect 230197 318547 230263 318550
rect 236494 318412 236500 318476
rect 236564 318474 236570 318476
rect 257061 318474 257127 318477
rect 236564 318472 257127 318474
rect 236564 318416 257066 318472
rect 257122 318416 257127 318472
rect 236564 318414 257127 318416
rect 273210 318474 273270 318550
rect 279601 318608 287714 318610
rect 279601 318552 279606 318608
rect 279662 318552 287714 318608
rect 279601 318550 287714 318552
rect 279601 318547 279667 318550
rect 284293 318474 284359 318477
rect 273210 318472 284359 318474
rect 273210 318416 284298 318472
rect 284354 318416 284359 318472
rect 273210 318414 284359 318416
rect 287654 318474 287714 318550
rect 289077 318608 292804 318610
rect 289077 318552 289082 318608
rect 289138 318552 292804 318608
rect 289077 318550 292804 318552
rect 289077 318547 289143 318550
rect 292798 318548 292804 318550
rect 292868 318548 292874 318612
rect 292944 318610 293004 318686
rect 294597 318684 294644 318686
rect 294708 318684 294714 318748
rect 296662 318684 296668 318748
rect 296732 318746 296738 318748
rect 297950 318746 297956 318748
rect 296732 318686 297956 318746
rect 296732 318684 296738 318686
rect 297950 318684 297956 318686
rect 298020 318684 298026 318748
rect 300577 318746 300643 318749
rect 300710 318746 300716 318748
rect 300577 318744 300716 318746
rect 300577 318688 300582 318744
rect 300638 318688 300716 318744
rect 300577 318686 300716 318688
rect 294597 318683 294663 318684
rect 300577 318683 300643 318686
rect 300710 318684 300716 318686
rect 300780 318684 300786 318748
rect 306373 318746 306439 318749
rect 307518 318746 307524 318748
rect 306373 318744 307524 318746
rect 306373 318688 306378 318744
rect 306434 318688 307524 318744
rect 306373 318686 307524 318688
rect 306373 318683 306439 318686
rect 307518 318684 307524 318686
rect 307588 318684 307594 318748
rect 308070 318684 308076 318748
rect 308140 318746 308146 318748
rect 308489 318746 308555 318749
rect 308140 318744 308555 318746
rect 308140 318688 308494 318744
rect 308550 318688 308555 318744
rect 308140 318686 308555 318688
rect 308140 318684 308146 318686
rect 308489 318683 308555 318686
rect 313641 318746 313707 318749
rect 314326 318746 314332 318748
rect 313641 318744 314332 318746
rect 313641 318688 313646 318744
rect 313702 318688 314332 318744
rect 313641 318686 314332 318688
rect 313641 318683 313707 318686
rect 314326 318684 314332 318686
rect 314396 318684 314402 318748
rect 320357 318746 320423 318749
rect 321093 318746 321159 318749
rect 325509 318748 325575 318749
rect 325509 318746 325556 318748
rect 320357 318744 321159 318746
rect 320357 318688 320362 318744
rect 320418 318688 321098 318744
rect 321154 318688 321159 318744
rect 320357 318686 321159 318688
rect 325464 318744 325556 318746
rect 325464 318688 325514 318744
rect 325464 318686 325556 318688
rect 320357 318683 320423 318686
rect 321093 318683 321159 318686
rect 325509 318684 325556 318686
rect 325620 318684 325626 318748
rect 330109 318746 330175 318749
rect 327030 318744 330175 318746
rect 327030 318688 330114 318744
rect 330170 318688 330175 318744
rect 327030 318686 330175 318688
rect 325509 318683 325575 318684
rect 295793 318610 295859 318613
rect 292944 318608 295859 318610
rect 292944 318552 295798 318608
rect 295854 318552 295859 318608
rect 292944 318550 295859 318552
rect 295793 318547 295859 318550
rect 297357 318610 297423 318613
rect 319345 318610 319411 318613
rect 323342 318610 323348 318612
rect 297357 318608 311910 318610
rect 297357 318552 297362 318608
rect 297418 318552 311910 318608
rect 297357 318550 311910 318552
rect 297357 318547 297423 318550
rect 287654 318414 292590 318474
rect 236564 318412 236570 318414
rect 257061 318411 257127 318414
rect 284293 318411 284359 318414
rect 237966 318276 237972 318340
rect 238036 318338 238042 318340
rect 272609 318338 272675 318341
rect 238036 318336 272675 318338
rect 238036 318280 272614 318336
rect 272670 318280 272675 318336
rect 238036 318278 272675 318280
rect 238036 318276 238042 318278
rect 272609 318275 272675 318278
rect 285806 318276 285812 318340
rect 285876 318338 285882 318340
rect 286225 318338 286291 318341
rect 285876 318336 286291 318338
rect 285876 318280 286230 318336
rect 286286 318280 286291 318336
rect 285876 318278 286291 318280
rect 285876 318276 285882 318278
rect 286225 318275 286291 318278
rect 289813 318338 289879 318341
rect 292062 318338 292068 318340
rect 289813 318336 292068 318338
rect 289813 318280 289818 318336
rect 289874 318280 292068 318336
rect 289813 318278 292068 318280
rect 289813 318275 289879 318278
rect 292062 318276 292068 318278
rect 292132 318276 292138 318340
rect 292530 318338 292590 318414
rect 296846 318412 296852 318476
rect 296916 318474 296922 318476
rect 297541 318474 297607 318477
rect 296916 318472 297607 318474
rect 296916 318416 297546 318472
rect 297602 318416 297607 318472
rect 296916 318414 297607 318416
rect 296916 318412 296922 318414
rect 297541 318411 297607 318414
rect 300710 318412 300716 318476
rect 300780 318474 300786 318476
rect 302233 318474 302299 318477
rect 300780 318472 302299 318474
rect 300780 318416 302238 318472
rect 302294 318416 302299 318472
rect 300780 318414 302299 318416
rect 300780 318412 300786 318414
rect 302233 318411 302299 318414
rect 306465 318474 306531 318477
rect 306966 318474 306972 318476
rect 306465 318472 306972 318474
rect 306465 318416 306470 318472
rect 306526 318416 306972 318472
rect 306465 318414 306972 318416
rect 306465 318411 306531 318414
rect 306966 318412 306972 318414
rect 307036 318412 307042 318476
rect 308305 318338 308371 318341
rect 292530 318336 308371 318338
rect 292530 318280 308310 318336
rect 308366 318280 308371 318336
rect 292530 318278 308371 318280
rect 308305 318275 308371 318278
rect 206737 318202 206803 318205
rect 263685 318202 263751 318205
rect 289537 318202 289603 318205
rect 297357 318202 297423 318205
rect 302785 318202 302851 318205
rect 206737 318200 263751 318202
rect 206737 318144 206742 318200
rect 206798 318144 263690 318200
rect 263746 318144 263751 318200
rect 206737 318142 263751 318144
rect 206737 318139 206803 318142
rect 263685 318139 263751 318142
rect 273210 318200 297423 318202
rect 273210 318144 289542 318200
rect 289598 318144 297362 318200
rect 297418 318144 297423 318200
rect 273210 318142 297423 318144
rect 210785 318066 210851 318069
rect 273210 318066 273270 318142
rect 289537 318139 289603 318142
rect 297357 318139 297423 318142
rect 300074 318200 302851 318202
rect 300074 318144 302790 318200
rect 302846 318144 302851 318200
rect 300074 318142 302851 318144
rect 311850 318202 311910 318550
rect 319345 318608 323348 318610
rect 319345 318552 319350 318608
rect 319406 318552 323348 318608
rect 319345 318550 323348 318552
rect 319345 318547 319411 318550
rect 323342 318548 323348 318550
rect 323412 318548 323418 318612
rect 324405 318610 324471 318613
rect 327030 318610 327090 318686
rect 330109 318683 330175 318686
rect 324405 318608 327090 318610
rect 324405 318552 324410 318608
rect 324466 318552 327090 318608
rect 324405 318550 327090 318552
rect 327257 318610 327323 318613
rect 331397 318610 331463 318613
rect 327257 318608 331463 318610
rect 327257 318552 327262 318608
rect 327318 318552 331402 318608
rect 331458 318552 331463 318608
rect 327257 318550 331463 318552
rect 324405 318547 324471 318550
rect 327257 318547 327323 318550
rect 331397 318547 331463 318550
rect 320081 318474 320147 318477
rect 322013 318474 322079 318477
rect 335169 318474 335235 318477
rect 320081 318472 321938 318474
rect 320081 318416 320086 318472
rect 320142 318416 321938 318472
rect 320081 318414 321938 318416
rect 320081 318411 320147 318414
rect 314653 318338 314719 318341
rect 318885 318338 318951 318341
rect 314653 318336 318951 318338
rect 314653 318280 314658 318336
rect 314714 318280 318890 318336
rect 318946 318280 318951 318336
rect 314653 318278 318951 318280
rect 314653 318275 314719 318278
rect 318885 318275 318951 318278
rect 320725 318338 320791 318341
rect 321318 318338 321324 318340
rect 320725 318336 321324 318338
rect 320725 318280 320730 318336
rect 320786 318280 321324 318336
rect 320725 318278 321324 318280
rect 320725 318275 320791 318278
rect 321318 318276 321324 318278
rect 321388 318276 321394 318340
rect 321878 318338 321938 318414
rect 322013 318472 335235 318474
rect 322013 318416 322018 318472
rect 322074 318416 335174 318472
rect 335230 318416 335235 318472
rect 322013 318414 335235 318416
rect 322013 318411 322079 318414
rect 335169 318411 335235 318414
rect 324037 318338 324103 318341
rect 328085 318338 328151 318341
rect 321878 318336 324103 318338
rect 321878 318280 324042 318336
rect 324098 318280 324103 318336
rect 321878 318278 324103 318280
rect 324037 318275 324103 318278
rect 324270 318336 328151 318338
rect 324270 318280 328090 318336
rect 328146 318280 328151 318336
rect 324270 318278 328151 318280
rect 324270 318202 324330 318278
rect 328085 318275 328151 318278
rect 311850 318142 324330 318202
rect 325877 318202 325943 318205
rect 329925 318202 329991 318205
rect 367686 318202 367692 318204
rect 325877 318200 328746 318202
rect 325877 318144 325882 318200
rect 325938 318144 328746 318200
rect 325877 318142 328746 318144
rect 210785 318064 273270 318066
rect 210785 318008 210790 318064
rect 210846 318008 273270 318064
rect 210785 318006 273270 318008
rect 210785 318003 210851 318006
rect 285622 318004 285628 318068
rect 285692 318066 285698 318068
rect 286542 318066 286548 318068
rect 285692 318006 286548 318066
rect 285692 318004 285698 318006
rect 286542 318004 286548 318006
rect 286612 318004 286618 318068
rect 287329 318066 287395 318069
rect 287605 318066 287671 318069
rect 290549 318068 290615 318069
rect 289118 318066 289124 318068
rect 287329 318064 289124 318066
rect 287329 318008 287334 318064
rect 287390 318008 287610 318064
rect 287666 318008 289124 318064
rect 287329 318006 289124 318008
rect 287329 318003 287395 318006
rect 287605 318003 287671 318006
rect 289118 318004 289124 318006
rect 289188 318004 289194 318068
rect 290549 318066 290596 318068
rect 290504 318064 290596 318066
rect 290504 318008 290554 318064
rect 290504 318006 290596 318008
rect 290549 318004 290596 318006
rect 290660 318004 290666 318068
rect 290917 318066 290983 318069
rect 292430 318066 292436 318068
rect 290917 318064 292436 318066
rect 290917 318008 290922 318064
rect 290978 318008 292436 318064
rect 290917 318006 292436 318008
rect 290549 318003 290615 318004
rect 290917 318003 290983 318006
rect 292430 318004 292436 318006
rect 292500 318004 292506 318068
rect 293401 318066 293467 318069
rect 300074 318066 300134 318142
rect 302785 318139 302851 318142
rect 325877 318139 325943 318142
rect 293401 318064 300134 318066
rect 293401 318008 293406 318064
rect 293462 318008 300134 318064
rect 293401 318006 300134 318008
rect 300209 318066 300275 318069
rect 302734 318066 302740 318068
rect 300209 318064 302740 318066
rect 300209 318008 300214 318064
rect 300270 318008 302740 318064
rect 300209 318006 302740 318008
rect 293401 318003 293467 318006
rect 300209 318003 300275 318006
rect 302734 318004 302740 318006
rect 302804 318004 302810 318068
rect 304758 318004 304764 318068
rect 304828 318066 304834 318068
rect 314929 318066 314995 318069
rect 315062 318066 315068 318068
rect 304828 318006 311910 318066
rect 304828 318004 304834 318006
rect 283925 317930 283991 317933
rect 284518 317930 284524 317932
rect 283925 317928 284524 317930
rect 283925 317872 283930 317928
rect 283986 317872 284524 317928
rect 283925 317870 284524 317872
rect 283925 317867 283991 317870
rect 284518 317868 284524 317870
rect 284588 317868 284594 317932
rect 287094 317868 287100 317932
rect 287164 317930 287170 317932
rect 287973 317930 288039 317933
rect 287164 317928 288039 317930
rect 287164 317872 287978 317928
rect 288034 317872 288039 317928
rect 287164 317870 288039 317872
rect 287164 317868 287170 317870
rect 287973 317867 288039 317870
rect 288382 317868 288388 317932
rect 288452 317930 288458 317932
rect 289169 317930 289235 317933
rect 303797 317930 303863 317933
rect 288452 317928 289235 317930
rect 288452 317872 289174 317928
rect 289230 317872 289235 317928
rect 288452 317870 289235 317872
rect 288452 317868 288458 317870
rect 289169 317867 289235 317870
rect 292530 317928 303863 317930
rect 292530 317872 303802 317928
rect 303858 317872 303863 317928
rect 292530 317870 303863 317872
rect 282637 317794 282703 317797
rect 292530 317794 292590 317870
rect 303797 317867 303863 317870
rect 306373 317930 306439 317933
rect 306598 317930 306604 317932
rect 306373 317928 306604 317930
rect 306373 317872 306378 317928
rect 306434 317872 306604 317928
rect 306373 317870 306604 317872
rect 306373 317867 306439 317870
rect 306598 317868 306604 317870
rect 306668 317868 306674 317932
rect 311850 317930 311910 318006
rect 314929 318064 315068 318066
rect 314929 318008 314934 318064
rect 314990 318008 315068 318064
rect 314929 318006 315068 318008
rect 314929 318003 314995 318006
rect 315062 318004 315068 318006
rect 315132 318004 315138 318068
rect 316534 318004 316540 318068
rect 316604 318066 316610 318068
rect 317137 318066 317203 318069
rect 316604 318064 317203 318066
rect 316604 318008 317142 318064
rect 317198 318008 317203 318064
rect 316604 318006 317203 318008
rect 316604 318004 316610 318006
rect 317137 318003 317203 318006
rect 317454 318004 317460 318068
rect 317524 318066 317530 318068
rect 318701 318066 318767 318069
rect 317524 318064 318767 318066
rect 317524 318008 318706 318064
rect 318762 318008 318767 318064
rect 317524 318006 318767 318008
rect 317524 318004 317530 318006
rect 318701 318003 318767 318006
rect 320265 318066 320331 318069
rect 326654 318066 326660 318068
rect 320265 318064 326660 318066
rect 320265 318008 320270 318064
rect 320326 318008 326660 318064
rect 320265 318006 326660 318008
rect 320265 318003 320331 318006
rect 326654 318004 326660 318006
rect 326724 318004 326730 318068
rect 328269 318066 328335 318069
rect 327214 318064 328335 318066
rect 327214 318008 328274 318064
rect 328330 318008 328335 318064
rect 327214 318006 328335 318008
rect 318149 317930 318215 317933
rect 318793 317932 318859 317933
rect 311850 317928 318215 317930
rect 311850 317872 318154 317928
rect 318210 317872 318215 317928
rect 311850 317870 318215 317872
rect 318149 317867 318215 317870
rect 318742 317868 318748 317932
rect 318812 317930 318859 317932
rect 318812 317928 318904 317930
rect 318854 317872 318904 317928
rect 318812 317870 318904 317872
rect 318812 317868 318859 317870
rect 320766 317868 320772 317932
rect 320836 317930 320842 317932
rect 321001 317930 321067 317933
rect 322841 317932 322907 317933
rect 322790 317930 322796 317932
rect 320836 317928 321067 317930
rect 320836 317872 321006 317928
rect 321062 317872 321067 317928
rect 320836 317870 321067 317872
rect 322750 317870 322796 317930
rect 322860 317928 322907 317932
rect 322902 317872 322907 317928
rect 320836 317868 320842 317870
rect 318793 317867 318859 317868
rect 321001 317867 321067 317870
rect 322790 317868 322796 317870
rect 322860 317868 322907 317872
rect 324446 317868 324452 317932
rect 324516 317930 324522 317932
rect 324957 317930 325023 317933
rect 324516 317928 325023 317930
rect 324516 317872 324962 317928
rect 325018 317872 325023 317928
rect 324516 317870 325023 317872
rect 324516 317868 324522 317870
rect 322841 317867 322907 317868
rect 324957 317867 325023 317870
rect 325877 317930 325943 317933
rect 327214 317930 327274 318006
rect 328269 318003 328335 318006
rect 325877 317928 327274 317930
rect 325877 317872 325882 317928
rect 325938 317872 327274 317928
rect 325877 317870 327274 317872
rect 327349 317930 327415 317933
rect 328686 317932 328746 318142
rect 329925 318200 367692 318202
rect 329925 318144 329930 318200
rect 329986 318144 367692 318200
rect 329925 318142 367692 318144
rect 329925 318139 329991 318142
rect 367686 318140 367692 318142
rect 367756 318140 367762 318204
rect 329833 318066 329899 318069
rect 369894 318066 369900 318068
rect 329833 318064 369900 318066
rect 329833 318008 329838 318064
rect 329894 318008 369900 318064
rect 329833 318006 369900 318008
rect 329833 318003 329899 318006
rect 369894 318004 369900 318006
rect 369964 318004 369970 318068
rect 327574 317930 327580 317932
rect 327349 317928 327580 317930
rect 327349 317872 327354 317928
rect 327410 317872 327580 317928
rect 327349 317870 327580 317872
rect 325877 317867 325943 317870
rect 327349 317867 327415 317870
rect 327574 317868 327580 317870
rect 327644 317868 327650 317932
rect 328678 317868 328684 317932
rect 328748 317930 328754 317932
rect 329557 317930 329623 317933
rect 328748 317928 329623 317930
rect 328748 317872 329562 317928
rect 329618 317872 329623 317928
rect 328748 317870 329623 317872
rect 328748 317868 328754 317870
rect 329557 317867 329623 317870
rect 300577 317796 300643 317797
rect 282637 317792 292590 317794
rect 282637 317736 282642 317792
rect 282698 317736 292590 317792
rect 282637 317734 292590 317736
rect 282637 317731 282703 317734
rect 300526 317732 300532 317796
rect 300596 317794 300643 317796
rect 300596 317792 300688 317794
rect 300638 317736 300688 317792
rect 300596 317734 300688 317736
rect 300596 317732 300643 317734
rect 301262 317732 301268 317796
rect 301332 317794 301338 317796
rect 302049 317794 302115 317797
rect 303337 317796 303403 317797
rect 303286 317794 303292 317796
rect 301332 317792 302115 317794
rect 301332 317736 302054 317792
rect 302110 317736 302115 317792
rect 301332 317734 302115 317736
rect 303246 317734 303292 317794
rect 303356 317792 303403 317796
rect 303398 317736 303403 317792
rect 301332 317732 301338 317734
rect 300577 317731 300643 317732
rect 302049 317731 302115 317734
rect 303286 317732 303292 317734
rect 303356 317732 303403 317736
rect 303337 317731 303403 317732
rect 304257 317794 304323 317797
rect 305310 317794 305316 317796
rect 304257 317792 305316 317794
rect 304257 317736 304262 317792
rect 304318 317736 305316 317792
rect 304257 317734 305316 317736
rect 304257 317731 304323 317734
rect 305310 317732 305316 317734
rect 305380 317794 305386 317796
rect 306189 317794 306255 317797
rect 305380 317792 306255 317794
rect 305380 317736 306194 317792
rect 306250 317736 306255 317792
rect 305380 317734 306255 317736
rect 305380 317732 305386 317734
rect 306189 317731 306255 317734
rect 307702 317732 307708 317796
rect 307772 317794 307778 317796
rect 308857 317794 308923 317797
rect 312905 317796 312971 317797
rect 307772 317792 308923 317794
rect 307772 317736 308862 317792
rect 308918 317736 308923 317792
rect 307772 317734 308923 317736
rect 307772 317732 307778 317734
rect 308857 317731 308923 317734
rect 309726 317732 309732 317796
rect 309796 317794 309802 317796
rect 310278 317794 310284 317796
rect 309796 317734 310284 317794
rect 309796 317732 309802 317734
rect 310278 317732 310284 317734
rect 310348 317732 310354 317796
rect 312854 317732 312860 317796
rect 312924 317794 312971 317796
rect 312924 317792 313016 317794
rect 312966 317736 313016 317792
rect 312924 317734 313016 317736
rect 312924 317732 312971 317734
rect 316166 317732 316172 317796
rect 316236 317794 316242 317796
rect 317321 317794 317387 317797
rect 316236 317792 317387 317794
rect 316236 317736 317326 317792
rect 317382 317736 317387 317792
rect 316236 317734 317387 317736
rect 316236 317732 316242 317734
rect 312905 317731 312971 317732
rect 317321 317731 317387 317734
rect 317781 317794 317847 317797
rect 318190 317794 318196 317796
rect 317781 317792 318196 317794
rect 317781 317736 317786 317792
rect 317842 317736 318196 317792
rect 317781 317734 318196 317736
rect 317781 317731 317847 317734
rect 318190 317732 318196 317734
rect 318260 317732 318266 317796
rect 318885 317794 318951 317797
rect 325550 317794 325556 317796
rect 318885 317792 325556 317794
rect 318885 317736 318890 317792
rect 318946 317736 325556 317792
rect 318885 317734 325556 317736
rect 318885 317731 318951 317734
rect 325550 317732 325556 317734
rect 325620 317732 325626 317796
rect 327022 317732 327028 317796
rect 327092 317794 327098 317796
rect 327441 317794 327507 317797
rect 327092 317792 327507 317794
rect 327092 317736 327446 317792
rect 327502 317736 327507 317792
rect 327092 317734 327507 317736
rect 327092 317732 327098 317734
rect 327441 317731 327507 317734
rect 263685 317658 263751 317661
rect 264881 317658 264947 317661
rect 284661 317658 284727 317661
rect 263685 317656 284727 317658
rect 263685 317600 263690 317656
rect 263746 317600 264886 317656
rect 264942 317600 284666 317656
rect 284722 317600 284727 317656
rect 263685 317598 284727 317600
rect 263685 317595 263751 317598
rect 264881 317595 264947 317598
rect 284661 317595 284727 317598
rect 286225 317658 286291 317661
rect 286501 317658 286567 317661
rect 286225 317656 286567 317658
rect 286225 317600 286230 317656
rect 286286 317600 286506 317656
rect 286562 317600 286567 317656
rect 286225 317598 286567 317600
rect 286225 317595 286291 317598
rect 286501 317595 286567 317598
rect 287329 317658 287395 317661
rect 322013 317658 322079 317661
rect 287329 317656 322079 317658
rect 287329 317600 287334 317656
rect 287390 317600 322018 317656
rect 322074 317600 322079 317656
rect 287329 317598 322079 317600
rect 287329 317595 287395 317598
rect 322013 317595 322079 317598
rect 322197 317658 322263 317661
rect 322790 317658 322796 317660
rect 322197 317656 322796 317658
rect 322197 317600 322202 317656
rect 322258 317600 322796 317656
rect 322197 317598 322796 317600
rect 322197 317595 322263 317598
rect 322790 317596 322796 317598
rect 322860 317596 322866 317660
rect 323485 317658 323551 317661
rect 327441 317658 327507 317661
rect 323485 317656 327507 317658
rect 323485 317600 323490 317656
rect 323546 317600 327446 317656
rect 327502 317600 327507 317656
rect 323485 317598 327507 317600
rect 323485 317595 323551 317598
rect 327441 317595 327507 317598
rect 278313 317522 278379 317525
rect 279601 317522 279667 317525
rect 278313 317520 279667 317522
rect 278313 317464 278318 317520
rect 278374 317464 279606 317520
rect 279662 317464 279667 317520
rect 278313 317462 279667 317464
rect 278313 317459 278379 317462
rect 279601 317459 279667 317462
rect 283046 317460 283052 317524
rect 283116 317522 283122 317524
rect 283557 317522 283623 317525
rect 283116 317520 283623 317522
rect 283116 317464 283562 317520
rect 283618 317464 283623 317520
rect 283116 317462 283623 317464
rect 283116 317460 283122 317462
rect 283557 317459 283623 317462
rect 284334 317460 284340 317524
rect 284404 317522 284410 317524
rect 284937 317522 285003 317525
rect 284404 317520 285003 317522
rect 284404 317464 284942 317520
rect 284998 317464 285003 317520
rect 284404 317462 285003 317464
rect 284404 317460 284410 317462
rect 284937 317459 285003 317462
rect 285121 317522 285187 317525
rect 290774 317522 290780 317524
rect 285121 317520 290780 317522
rect 285121 317464 285126 317520
rect 285182 317464 290780 317520
rect 285121 317462 290780 317464
rect 285121 317459 285187 317462
rect 290774 317460 290780 317462
rect 290844 317522 290850 317524
rect 291694 317522 291700 317524
rect 290844 317462 291700 317522
rect 290844 317460 290850 317462
rect 291694 317460 291700 317462
rect 291764 317460 291770 317524
rect 299606 317460 299612 317524
rect 299676 317522 299682 317524
rect 300117 317522 300183 317525
rect 299676 317520 300183 317522
rect 299676 317464 300122 317520
rect 300178 317464 300183 317520
rect 299676 317462 300183 317464
rect 299676 317460 299682 317462
rect 300117 317459 300183 317462
rect 301078 317460 301084 317524
rect 301148 317522 301154 317524
rect 301405 317522 301471 317525
rect 301148 317520 301471 317522
rect 301148 317464 301410 317520
rect 301466 317464 301471 317520
rect 301148 317462 301471 317464
rect 301148 317460 301154 317462
rect 301405 317459 301471 317462
rect 301773 317522 301839 317525
rect 301998 317522 302004 317524
rect 301773 317520 302004 317522
rect 301773 317464 301778 317520
rect 301834 317464 302004 317520
rect 301773 317462 302004 317464
rect 301773 317459 301839 317462
rect 301998 317460 302004 317462
rect 302068 317460 302074 317524
rect 302601 317522 302667 317525
rect 302734 317522 302740 317524
rect 302601 317520 302740 317522
rect 302601 317464 302606 317520
rect 302662 317464 302740 317520
rect 302601 317462 302740 317464
rect 302601 317459 302667 317462
rect 302734 317460 302740 317462
rect 302804 317460 302810 317524
rect 303153 317522 303219 317525
rect 303470 317522 303476 317524
rect 303153 317520 303476 317522
rect 303153 317464 303158 317520
rect 303214 317464 303476 317520
rect 303153 317462 303476 317464
rect 303153 317459 303219 317462
rect 303470 317460 303476 317462
rect 303540 317460 303546 317524
rect 305494 317460 305500 317524
rect 305564 317522 305570 317524
rect 306281 317522 306347 317525
rect 306833 317524 306899 317525
rect 306782 317522 306788 317524
rect 305564 317520 306347 317522
rect 305564 317464 306286 317520
rect 306342 317464 306347 317520
rect 305564 317462 306347 317464
rect 306742 317462 306788 317522
rect 306852 317520 306899 317524
rect 306894 317464 306899 317520
rect 305564 317460 305570 317462
rect 306281 317459 306347 317462
rect 306782 317460 306788 317462
rect 306852 317460 306899 317464
rect 306833 317459 306899 317460
rect 307753 317522 307819 317525
rect 309777 317524 309843 317525
rect 309961 317524 310027 317525
rect 308254 317522 308260 317524
rect 307753 317520 308260 317522
rect 307753 317464 307758 317520
rect 307814 317464 308260 317520
rect 307753 317462 308260 317464
rect 307753 317459 307819 317462
rect 308254 317460 308260 317462
rect 308324 317460 308330 317524
rect 309726 317522 309732 317524
rect 309686 317462 309732 317522
rect 309796 317520 309843 317524
rect 309838 317464 309843 317520
rect 309726 317460 309732 317462
rect 309796 317460 309843 317464
rect 309910 317460 309916 317524
rect 309980 317522 310027 317524
rect 311893 317522 311959 317525
rect 313038 317522 313044 317524
rect 309980 317520 310072 317522
rect 310022 317464 310072 317520
rect 309980 317462 310072 317464
rect 311893 317520 313044 317522
rect 311893 317464 311898 317520
rect 311954 317464 313044 317520
rect 311893 317462 313044 317464
rect 309980 317460 310027 317462
rect 309777 317459 309843 317460
rect 309961 317459 310027 317460
rect 311893 317459 311959 317462
rect 313038 317460 313044 317462
rect 313108 317460 313114 317524
rect 313406 317460 313412 317524
rect 313476 317522 313482 317524
rect 313825 317522 313891 317525
rect 313476 317520 313891 317522
rect 313476 317464 313830 317520
rect 313886 317464 313891 317520
rect 313476 317462 313891 317464
rect 313476 317460 313482 317462
rect 313825 317459 313891 317462
rect 314469 317524 314535 317525
rect 314469 317520 314516 317524
rect 314580 317522 314586 317524
rect 318057 317522 318123 317525
rect 318374 317522 318380 317524
rect 314469 317464 314474 317520
rect 314469 317460 314516 317464
rect 314580 317462 314626 317522
rect 318057 317520 318380 317522
rect 318057 317464 318062 317520
rect 318118 317464 318380 317520
rect 318057 317462 318380 317464
rect 314580 317460 314586 317462
rect 314469 317459 314535 317460
rect 318057 317459 318123 317462
rect 318374 317460 318380 317462
rect 318444 317460 318450 317524
rect 320582 317460 320588 317524
rect 320652 317522 320658 317524
rect 320909 317522 320975 317525
rect 320652 317520 320975 317522
rect 320652 317464 320914 317520
rect 320970 317464 320975 317520
rect 320652 317462 320975 317464
rect 320652 317460 320658 317462
rect 320909 317459 320975 317462
rect 321093 317522 321159 317525
rect 322657 317524 322723 317525
rect 322606 317522 322612 317524
rect 321093 317520 322490 317522
rect 321093 317464 321098 317520
rect 321154 317464 322490 317520
rect 321093 317462 322490 317464
rect 322566 317462 322612 317522
rect 322676 317520 322723 317524
rect 325877 317522 325943 317525
rect 322718 317464 322723 317520
rect 321093 317459 321159 317462
rect 269849 317386 269915 317389
rect 284385 317386 284451 317389
rect 258030 317384 284451 317386
rect 258030 317328 269854 317384
rect 269910 317328 284390 317384
rect 284446 317328 284451 317384
rect 258030 317326 284451 317328
rect 223246 317052 223252 317116
rect 223316 317114 223322 317116
rect 244273 317114 244339 317117
rect 223316 317112 244339 317114
rect 223316 317056 244278 317112
rect 244334 317056 244339 317112
rect 223316 317054 244339 317056
rect 223316 317052 223322 317054
rect 244273 317051 244339 317054
rect 223430 316916 223436 316980
rect 223500 316978 223506 316980
rect 253749 316978 253815 316981
rect 223500 316976 253815 316978
rect 223500 316920 253754 316976
rect 253810 316920 253815 316976
rect 223500 316918 253815 316920
rect 223500 316916 223506 316918
rect 253749 316915 253815 316918
rect 215109 316842 215175 316845
rect 258030 316842 258090 317326
rect 269849 317323 269915 317326
rect 284385 317323 284451 317326
rect 287646 317324 287652 317388
rect 287716 317386 287722 317388
rect 292430 317386 292436 317388
rect 287716 317326 292436 317386
rect 287716 317324 287722 317326
rect 292430 317324 292436 317326
rect 292500 317324 292506 317388
rect 322430 317386 322490 317462
rect 322606 317460 322612 317462
rect 322676 317460 322723 317464
rect 322657 317459 322723 317460
rect 322798 317520 325943 317522
rect 322798 317464 325882 317520
rect 325938 317464 325943 317520
rect 322798 317462 325943 317464
rect 322798 317386 322858 317462
rect 325877 317459 325943 317462
rect 326245 317522 326311 317525
rect 326797 317524 326863 317525
rect 326245 317520 326722 317522
rect 326245 317464 326250 317520
rect 326306 317464 326722 317520
rect 326245 317462 326722 317464
rect 326245 317459 326311 317462
rect 322430 317326 322858 317386
rect 325049 317386 325115 317389
rect 326521 317386 326587 317389
rect 325049 317384 326587 317386
rect 325049 317328 325054 317384
rect 325110 317328 326526 317384
rect 326582 317328 326587 317384
rect 325049 317326 326587 317328
rect 326662 317386 326722 317462
rect 326797 317520 326844 317524
rect 326908 317522 326914 317524
rect 326797 317464 326802 317520
rect 326797 317460 326844 317464
rect 326908 317462 326954 317522
rect 326908 317460 326914 317462
rect 326797 317459 326863 317460
rect 327901 317386 327967 317389
rect 385493 317386 385559 317389
rect 326662 317384 385559 317386
rect 326662 317328 327906 317384
rect 327962 317328 385498 317384
rect 385554 317328 385559 317384
rect 326662 317326 385559 317328
rect 325049 317323 325115 317326
rect 326521 317323 326587 317326
rect 327901 317323 327967 317326
rect 385493 317323 385559 317326
rect 271413 317250 271479 317253
rect 303654 317250 303660 317252
rect 271413 317248 303660 317250
rect 271413 317192 271418 317248
rect 271474 317192 303660 317248
rect 271413 317190 303660 317192
rect 271413 317187 271479 317190
rect 303654 317188 303660 317190
rect 303724 317188 303730 317252
rect 322473 317250 322539 317253
rect 352741 317250 352807 317253
rect 322473 317248 352807 317250
rect 322473 317192 322478 317248
rect 322534 317192 352746 317248
rect 352802 317192 352807 317248
rect 322473 317190 352807 317192
rect 322473 317187 322539 317190
rect 352741 317187 352807 317190
rect 274449 317114 274515 317117
rect 288433 317114 288499 317117
rect 274449 317112 288499 317114
rect 274449 317056 274454 317112
rect 274510 317056 288438 317112
rect 288494 317056 288499 317112
rect 274449 317054 288499 317056
rect 274449 317051 274515 317054
rect 288433 317051 288499 317054
rect 314837 317114 314903 317117
rect 336733 317114 336799 317117
rect 337929 317114 337995 317117
rect 339493 317114 339559 317117
rect 340689 317114 340755 317117
rect 314837 317112 337995 317114
rect 314837 317056 314842 317112
rect 314898 317056 336738 317112
rect 336794 317056 337934 317112
rect 337990 317056 337995 317112
rect 314837 317054 337995 317056
rect 314837 317051 314903 317054
rect 336733 317051 336799 317054
rect 337929 317051 337995 317054
rect 338438 317112 340755 317114
rect 338438 317056 339498 317112
rect 339554 317056 340694 317112
rect 340750 317056 340755 317112
rect 338438 317054 340755 317056
rect 281390 316916 281396 316980
rect 281460 316978 281466 316980
rect 315297 316978 315363 316981
rect 281460 316976 315363 316978
rect 281460 316920 315302 316976
rect 315358 316920 315363 316976
rect 281460 316918 315363 316920
rect 281460 316916 281466 316918
rect 315297 316915 315363 316918
rect 326654 316916 326660 316980
rect 326724 316978 326730 316980
rect 338438 316978 338498 317054
rect 339493 317051 339559 317054
rect 340689 317051 340755 317054
rect 326724 316918 338498 316978
rect 326724 316916 326730 316918
rect 215109 316840 258090 316842
rect 215109 316784 215114 316840
rect 215170 316784 258090 316840
rect 215109 316782 258090 316784
rect 282361 316842 282427 316845
rect 316677 316842 316743 316845
rect 282361 316840 316743 316842
rect 282361 316784 282366 316840
rect 282422 316784 316682 316840
rect 316738 316784 316743 316840
rect 282361 316782 316743 316784
rect 215109 316779 215175 316782
rect 282361 316779 282427 316782
rect 316677 316779 316743 316782
rect 325550 316780 325556 316844
rect 325620 316842 325626 316844
rect 338113 316842 338179 316845
rect 325620 316840 338179 316842
rect 325620 316784 338118 316840
rect 338174 316784 338179 316840
rect 325620 316782 338179 316784
rect 325620 316780 325626 316782
rect 338113 316779 338179 316782
rect 205449 316706 205515 316709
rect 284109 316706 284175 316709
rect 205449 316704 284175 316706
rect 205449 316648 205454 316704
rect 205510 316648 284114 316704
rect 284170 316648 284175 316704
rect 205449 316646 284175 316648
rect 205449 316643 205515 316646
rect 284109 316643 284175 316646
rect 296621 316706 296687 316709
rect 321737 316706 321803 316709
rect 322473 316706 322539 316709
rect 296621 316704 322539 316706
rect 296621 316648 296626 316704
rect 296682 316648 321742 316704
rect 321798 316648 322478 316704
rect 322534 316648 322539 316704
rect 296621 316646 322539 316648
rect 296621 316643 296687 316646
rect 321737 316643 321803 316646
rect 322473 316643 322539 316646
rect 326981 316706 327047 316709
rect 330109 316706 330175 316709
rect 340822 316706 340828 316708
rect 326981 316704 340828 316706
rect 326981 316648 326986 316704
rect 327042 316648 330114 316704
rect 330170 316648 340828 316704
rect 326981 316646 340828 316648
rect 326981 316643 327047 316646
rect 330109 316643 330175 316646
rect 340822 316644 340828 316646
rect 340892 316644 340898 316708
rect 298645 316570 298711 316573
rect 299422 316570 299428 316572
rect 298645 316568 299428 316570
rect 298645 316512 298650 316568
rect 298706 316512 299428 316568
rect 298645 316510 299428 316512
rect 298645 316507 298711 316510
rect 299422 316508 299428 316510
rect 299492 316508 299498 316572
rect 335353 316570 335419 316573
rect 335905 316570 335971 316573
rect 335310 316568 335971 316570
rect 335310 316512 335358 316568
rect 335414 316512 335910 316568
rect 335966 316512 335971 316568
rect 335310 316510 335971 316512
rect 335310 316507 335419 316510
rect 335905 316507 335971 316510
rect 298369 316434 298435 316437
rect 299238 316434 299244 316436
rect 298369 316432 299244 316434
rect 298369 316376 298374 316432
rect 298430 316376 299244 316432
rect 298369 316374 299244 316376
rect 298369 316371 298435 316374
rect 299238 316372 299244 316374
rect 299308 316372 299314 316436
rect 324037 316434 324103 316437
rect 335310 316434 335370 316507
rect 324037 316432 335370 316434
rect 324037 316376 324042 316432
rect 324098 316376 335370 316432
rect 324037 316374 335370 316376
rect 324037 316371 324103 316374
rect 298553 316298 298619 316301
rect 298870 316298 298876 316300
rect 298553 316296 298876 316298
rect 298553 316240 298558 316296
rect 298614 316240 298876 316296
rect 298553 316238 298876 316240
rect 298553 316235 298619 316238
rect 298870 316236 298876 316238
rect 298940 316236 298946 316300
rect 323669 316298 323735 316301
rect 327257 316298 327323 316301
rect 323669 316296 327323 316298
rect 323669 316240 323674 316296
rect 323730 316240 327262 316296
rect 327318 316240 327323 316296
rect 323669 316238 327323 316240
rect 323669 316235 323735 316238
rect 327257 316235 327323 316238
rect 281073 316162 281139 316165
rect 299473 316162 299539 316165
rect 281073 316160 299539 316162
rect 281073 316104 281078 316160
rect 281134 316104 299478 316160
rect 299534 316104 299539 316160
rect 281073 316102 299539 316104
rect 281073 316099 281139 316102
rect 299473 316099 299539 316102
rect 322381 316162 322447 316165
rect 323761 316162 323827 316165
rect 322381 316160 323827 316162
rect 322381 316104 322386 316160
rect 322442 316104 323766 316160
rect 323822 316104 323827 316160
rect 322381 316102 323827 316104
rect 322381 316099 322447 316102
rect 323761 316099 323827 316102
rect 222694 315964 222700 316028
rect 222764 316026 222770 316028
rect 264789 316026 264855 316029
rect 222764 316024 264855 316026
rect 222764 315968 264794 316024
rect 264850 315968 264855 316024
rect 222764 315966 264855 315968
rect 222764 315964 222770 315966
rect 264789 315963 264855 315966
rect 269573 316026 269639 316029
rect 284845 316026 284911 316029
rect 269573 316024 284911 316026
rect 269573 315968 269578 316024
rect 269634 315968 284850 316024
rect 284906 315968 284911 316024
rect 269573 315966 284911 315968
rect 269573 315963 269639 315966
rect 284845 315963 284911 315966
rect 298502 315964 298508 316028
rect 298572 316026 298578 316028
rect 299289 316026 299355 316029
rect 298572 316024 299355 316026
rect 298572 315968 299294 316024
rect 299350 315968 299355 316024
rect 298572 315966 299355 315968
rect 298572 315964 298578 315966
rect 299289 315963 299355 315966
rect 317045 316026 317111 316029
rect 377029 316026 377095 316029
rect 317045 316024 377095 316026
rect 317045 315968 317050 316024
rect 317106 315968 377034 316024
rect 377090 315968 377095 316024
rect 317045 315966 377095 315968
rect 317045 315963 317111 315966
rect 377029 315963 377095 315966
rect 214925 315890 214991 315893
rect 271045 315890 271111 315893
rect 214925 315888 271111 315890
rect 214925 315832 214930 315888
rect 214986 315832 271050 315888
rect 271106 315832 271111 315888
rect 214925 315830 271111 315832
rect 214925 315827 214991 315830
rect 271045 315827 271111 315830
rect 273621 315890 273687 315893
rect 296478 315890 296484 315892
rect 273621 315888 296484 315890
rect 273621 315832 273626 315888
rect 273682 315832 296484 315888
rect 273621 315830 296484 315832
rect 273621 315827 273687 315830
rect 296478 315828 296484 315830
rect 296548 315828 296554 315892
rect 326061 315890 326127 315893
rect 385125 315890 385191 315893
rect 326061 315888 385191 315890
rect 326061 315832 326066 315888
rect 326122 315832 385130 315888
rect 385186 315832 385191 315888
rect 326061 315830 385191 315832
rect 326061 315827 326127 315830
rect 385125 315827 385191 315830
rect 210877 315754 210943 315757
rect 268561 315754 268627 315757
rect 210877 315752 268627 315754
rect 210877 315696 210882 315752
rect 210938 315696 268566 315752
rect 268622 315696 268627 315752
rect 210877 315694 268627 315696
rect 210877 315691 210943 315694
rect 268561 315691 268627 315694
rect 269849 315754 269915 315757
rect 310053 315756 310119 315757
rect 296294 315754 296300 315756
rect 269849 315752 296300 315754
rect 269849 315696 269854 315752
rect 269910 315696 296300 315752
rect 269849 315694 296300 315696
rect 269849 315691 269915 315694
rect 296294 315692 296300 315694
rect 296364 315692 296370 315756
rect 310053 315752 310100 315756
rect 310164 315754 310170 315756
rect 326521 315754 326587 315757
rect 328453 315754 328519 315757
rect 310053 315696 310058 315752
rect 310053 315692 310100 315696
rect 310164 315694 310210 315754
rect 326521 315752 328519 315754
rect 326521 315696 326526 315752
rect 326582 315696 328458 315752
rect 328514 315696 328519 315752
rect 326521 315694 328519 315696
rect 310164 315692 310170 315694
rect 310053 315691 310119 315692
rect 326521 315691 326587 315694
rect 328453 315691 328519 315694
rect 328913 315754 328979 315757
rect 381905 315754 381971 315757
rect 328913 315752 381971 315754
rect 328913 315696 328918 315752
rect 328974 315696 381910 315752
rect 381966 315696 381971 315752
rect 328913 315694 381971 315696
rect 328913 315691 328979 315694
rect 381905 315691 381971 315694
rect 236678 315556 236684 315620
rect 236748 315618 236754 315620
rect 297030 315618 297036 315620
rect 236748 315558 297036 315618
rect 236748 315556 236754 315558
rect 297030 315556 297036 315558
rect 297100 315556 297106 315620
rect 310513 315618 310579 315621
rect 311157 315618 311223 315621
rect 365110 315618 365116 315620
rect 310513 315616 365116 315618
rect 310513 315560 310518 315616
rect 310574 315560 311162 315616
rect 311218 315560 365116 315616
rect 310513 315558 365116 315560
rect 310513 315555 310579 315558
rect 311157 315555 311223 315558
rect 365110 315556 365116 315558
rect 365180 315618 365186 315620
rect 367093 315618 367159 315621
rect 365180 315616 367159 315618
rect 365180 315560 367098 315616
rect 367154 315560 367159 315616
rect 365180 315558 367159 315560
rect 365180 315556 365186 315558
rect 367093 315555 367159 315558
rect 237046 315420 237052 315484
rect 237116 315482 237122 315484
rect 297398 315482 297404 315484
rect 237116 315422 297404 315482
rect 237116 315420 237122 315422
rect 297398 315420 297404 315422
rect 297468 315420 297474 315484
rect 324221 315482 324287 315485
rect 352414 315482 352420 315484
rect 324221 315480 352420 315482
rect 324221 315424 324226 315480
rect 324282 315424 352420 315480
rect 324221 315422 352420 315424
rect 324221 315419 324287 315422
rect 352414 315420 352420 315422
rect 352484 315420 352490 315484
rect 209589 315346 209655 315349
rect 276749 315346 276815 315349
rect 209589 315344 276815 315346
rect 209589 315288 209594 315344
rect 209650 315288 276754 315344
rect 276810 315288 276815 315344
rect 209589 315286 276815 315288
rect 209589 315283 209655 315286
rect 276749 315283 276815 315286
rect 319253 315346 319319 315349
rect 336917 315346 336983 315349
rect 319253 315344 336983 315346
rect 319253 315288 319258 315344
rect 319314 315288 336922 315344
rect 336978 315288 336983 315344
rect 319253 315286 336983 315288
rect 319253 315283 319319 315286
rect 336917 315283 336983 315286
rect 224718 315148 224724 315212
rect 224788 315210 224794 315212
rect 247033 315210 247099 315213
rect 224788 315208 247099 315210
rect 224788 315152 247038 315208
rect 247094 315152 247099 315208
rect 224788 315150 247099 315152
rect 224788 315148 224794 315150
rect 247033 315147 247099 315150
rect 268561 315210 268627 315213
rect 301078 315210 301084 315212
rect 268561 315208 301084 315210
rect 268561 315152 268566 315208
rect 268622 315152 301084 315208
rect 268561 315150 301084 315152
rect 268561 315147 268627 315150
rect 301078 315148 301084 315150
rect 301148 315148 301154 315212
rect 321553 315210 321619 315213
rect 328913 315210 328979 315213
rect 321553 315208 328979 315210
rect 321553 315152 321558 315208
rect 321614 315152 328918 315208
rect 328974 315152 328979 315208
rect 321553 315150 328979 315152
rect 321553 315147 321619 315150
rect 328913 315147 328979 315150
rect 244774 314604 244780 314668
rect 244844 314666 244850 314668
rect 275921 314666 275987 314669
rect 244844 314664 275987 314666
rect 244844 314608 275926 314664
rect 275982 314608 275987 314664
rect 244844 314606 275987 314608
rect 244844 314604 244850 314606
rect 275921 314603 275987 314606
rect 283649 314666 283715 314669
rect 288198 314666 288204 314668
rect 283649 314664 288204 314666
rect 283649 314608 283654 314664
rect 283710 314608 288204 314664
rect 283649 314606 288204 314608
rect 283649 314603 283715 314606
rect 288198 314604 288204 314606
rect 288268 314604 288274 314668
rect 306373 314666 306439 314669
rect 312445 314668 312511 314669
rect 306782 314666 306788 314668
rect 306373 314664 306788 314666
rect 306373 314608 306378 314664
rect 306434 314608 306788 314664
rect 306373 314606 306788 314608
rect 306373 314603 306439 314606
rect 306782 314604 306788 314606
rect 306852 314604 306858 314668
rect 312445 314664 312492 314668
rect 312556 314666 312562 314668
rect 312445 314608 312450 314664
rect 312445 314604 312492 314608
rect 312556 314606 312602 314666
rect 312556 314604 312562 314606
rect 312854 314604 312860 314668
rect 312924 314666 312930 314668
rect 313089 314666 313155 314669
rect 312924 314664 313155 314666
rect 312924 314608 313094 314664
rect 313150 314608 313155 314664
rect 312924 314606 313155 314608
rect 312924 314604 312930 314606
rect 312445 314603 312511 314604
rect 313089 314603 313155 314606
rect 319161 314666 319227 314669
rect 319897 314666 319963 314669
rect 319161 314664 319963 314666
rect 319161 314608 319166 314664
rect 319222 314608 319902 314664
rect 319958 314608 319963 314664
rect 319161 314606 319963 314608
rect 319161 314603 319227 314606
rect 319897 314603 319963 314606
rect 322289 314666 322355 314669
rect 322657 314666 322723 314669
rect 330845 314666 330911 314669
rect 389357 314666 389423 314669
rect 322289 314664 330402 314666
rect 322289 314608 322294 314664
rect 322350 314608 322662 314664
rect 322718 314608 330402 314664
rect 322289 314606 330402 314608
rect 322289 314603 322355 314606
rect 322657 314603 322723 314606
rect 232262 314468 232268 314532
rect 232332 314530 232338 314532
rect 269021 314530 269087 314533
rect 232332 314528 269087 314530
rect 232332 314472 269026 314528
rect 269082 314472 269087 314528
rect 232332 314470 269087 314472
rect 232332 314468 232338 314470
rect 269021 314467 269087 314470
rect 271597 314530 271663 314533
rect 301262 314530 301268 314532
rect 271597 314528 301268 314530
rect 271597 314472 271602 314528
rect 271658 314472 301268 314528
rect 271597 314470 301268 314472
rect 271597 314467 271663 314470
rect 301262 314468 301268 314470
rect 301332 314468 301338 314532
rect 312670 314468 312676 314532
rect 312740 314530 312746 314532
rect 312813 314530 312879 314533
rect 312740 314528 312879 314530
rect 312740 314472 312818 314528
rect 312874 314472 312879 314528
rect 312740 314470 312879 314472
rect 312740 314468 312746 314470
rect 312813 314467 312879 314470
rect 325325 314530 325391 314533
rect 330201 314530 330267 314533
rect 325325 314528 330267 314530
rect 325325 314472 325330 314528
rect 325386 314472 330206 314528
rect 330262 314472 330267 314528
rect 325325 314470 330267 314472
rect 330342 314530 330402 314606
rect 330845 314664 389423 314666
rect 330845 314608 330850 314664
rect 330906 314608 389362 314664
rect 389418 314608 389423 314664
rect 330845 314606 389423 314608
rect 330845 314603 330911 314606
rect 389357 314603 389423 314606
rect 388069 314530 388135 314533
rect 330342 314528 388135 314530
rect 330342 314472 388074 314528
rect 388130 314472 388135 314528
rect 330342 314470 388135 314472
rect 325325 314467 325391 314470
rect 330201 314467 330267 314470
rect 388069 314467 388135 314470
rect 232814 314332 232820 314396
rect 232884 314394 232890 314396
rect 274081 314394 274147 314397
rect 293217 314394 293283 314397
rect 232884 314392 293283 314394
rect 232884 314336 274086 314392
rect 274142 314336 293222 314392
rect 293278 314336 293283 314392
rect 232884 314334 293283 314336
rect 232884 314332 232890 314334
rect 274081 314331 274147 314334
rect 293217 314331 293283 314334
rect 325417 314394 325483 314397
rect 389449 314394 389515 314397
rect 325417 314392 389515 314394
rect 325417 314336 325422 314392
rect 325478 314336 389454 314392
rect 389510 314336 389515 314392
rect 325417 314334 389515 314336
rect 325417 314331 325483 314334
rect 389449 314331 389515 314334
rect 245510 314196 245516 314260
rect 245580 314258 245586 314260
rect 304574 314258 304580 314260
rect 245580 314198 304580 314258
rect 245580 314196 245586 314198
rect 304574 314196 304580 314198
rect 304644 314196 304650 314260
rect 326429 314258 326495 314261
rect 330017 314258 330083 314261
rect 326429 314256 330083 314258
rect 326429 314200 326434 314256
rect 326490 314200 330022 314256
rect 330078 314200 330083 314256
rect 326429 314198 330083 314200
rect 326429 314195 326495 314198
rect 330017 314195 330083 314198
rect 330201 314258 330267 314261
rect 387977 314258 388043 314261
rect 330201 314256 388043 314258
rect 330201 314200 330206 314256
rect 330262 314200 387982 314256
rect 388038 314200 388043 314256
rect 330201 314198 388043 314200
rect 330201 314195 330267 314198
rect 387977 314195 388043 314198
rect 242566 314060 242572 314124
rect 242636 314122 242642 314124
rect 302550 314122 302556 314124
rect 242636 314062 302556 314122
rect 242636 314060 242642 314062
rect 302550 314060 302556 314062
rect 302620 314060 302626 314124
rect 319529 314122 319595 314125
rect 379789 314122 379855 314125
rect 319529 314120 383670 314122
rect 319529 314064 319534 314120
rect 319590 314064 379794 314120
rect 379850 314064 383670 314120
rect 319529 314062 383670 314064
rect 319529 314059 319595 314062
rect 379789 314059 379855 314062
rect 241278 313924 241284 313988
rect 241348 313986 241354 313988
rect 299473 313986 299539 313989
rect 241348 313984 299539 313986
rect 241348 313928 299478 313984
rect 299534 313928 299539 313984
rect 241348 313926 299539 313928
rect 241348 313924 241354 313926
rect 299473 313923 299539 313926
rect 319897 313986 319963 313989
rect 356830 313986 356836 313988
rect 319897 313984 356836 313986
rect 319897 313928 319902 313984
rect 319958 313928 356836 313984
rect 319897 313926 356836 313928
rect 319897 313923 319963 313926
rect 356830 313924 356836 313926
rect 356900 313924 356906 313988
rect 383610 313986 383670 314062
rect 477493 313986 477559 313989
rect 383610 313984 477559 313986
rect 383610 313928 477498 313984
rect 477554 313928 477559 313984
rect 383610 313926 477559 313928
rect 477493 313923 477559 313926
rect 242750 313788 242756 313852
rect 242820 313850 242826 313852
rect 271597 313850 271663 313853
rect 242820 313848 271663 313850
rect 242820 313792 271602 313848
rect 271658 313792 271663 313848
rect 242820 313790 271663 313792
rect 242820 313788 242826 313790
rect 271597 313787 271663 313790
rect 287697 313850 287763 313853
rect 323853 313850 323919 313853
rect 330845 313850 330911 313853
rect 287697 313848 330911 313850
rect 287697 313792 287702 313848
rect 287758 313792 323858 313848
rect 323914 313792 330850 313848
rect 330906 313792 330911 313848
rect 287697 313790 330911 313792
rect 287697 313787 287763 313790
rect 323853 313787 323919 313790
rect 330845 313787 330911 313790
rect 269021 313714 269087 313717
rect 292757 313714 292823 313717
rect 269021 313712 292823 313714
rect 269021 313656 269026 313712
rect 269082 313656 292762 313712
rect 292818 313656 292823 313712
rect 269021 313654 292823 313656
rect 269021 313651 269087 313654
rect 292757 313651 292823 313654
rect 320817 313306 320883 313309
rect 321553 313306 321619 313309
rect 320817 313304 321619 313306
rect 320817 313248 320822 313304
rect 320878 313248 321558 313304
rect 321614 313248 321619 313304
rect 320817 313246 321619 313248
rect 320817 313243 320883 313246
rect 321553 313243 321619 313246
rect 309777 313172 309843 313173
rect 234102 313108 234108 313172
rect 234172 313170 234178 313172
rect 293350 313170 293356 313172
rect 234172 313110 293356 313170
rect 234172 313108 234178 313110
rect 293350 313108 293356 313110
rect 293420 313108 293426 313172
rect 309726 313108 309732 313172
rect 309796 313170 309843 313172
rect 312537 313170 312603 313173
rect 320766 313170 320772 313172
rect 309796 313168 309888 313170
rect 309838 313112 309888 313168
rect 309796 313110 309888 313112
rect 312537 313168 320772 313170
rect 312537 313112 312542 313168
rect 312598 313112 320772 313168
rect 312537 313110 320772 313112
rect 309796 313108 309843 313110
rect 309777 313107 309843 313108
rect 312537 313107 312603 313110
rect 320766 313108 320772 313110
rect 320836 313108 320842 313172
rect 323158 313108 323164 313172
rect 323228 313170 323234 313172
rect 323577 313170 323643 313173
rect 323228 313168 323643 313170
rect 323228 313112 323582 313168
rect 323638 313112 323643 313168
rect 323228 313110 323643 313112
rect 323228 313108 323234 313110
rect 323577 313107 323643 313110
rect 324221 313170 324287 313173
rect 392209 313170 392275 313173
rect 324221 313168 392275 313170
rect 324221 313112 324226 313168
rect 324282 313112 392214 313168
rect 392270 313112 392275 313168
rect 324221 313110 392275 313112
rect 324221 313107 324287 313110
rect 392209 313107 392275 313110
rect 249558 312972 249564 313036
rect 249628 313034 249634 313036
rect 309174 313034 309180 313036
rect 249628 312974 309180 313034
rect 249628 312972 249634 312974
rect 309174 312972 309180 312974
rect 309244 312972 309250 313036
rect 323117 313034 323183 313037
rect 324129 313034 324195 313037
rect 323117 313032 324195 313034
rect 323117 312976 323122 313032
rect 323178 312976 324134 313032
rect 324190 312976 324195 313032
rect 323117 312974 324195 312976
rect 323117 312971 323183 312974
rect 324129 312971 324195 312974
rect 326521 313034 326587 313037
rect 326889 313034 326955 313037
rect 326521 313032 393330 313034
rect 326521 312976 326526 313032
rect 326582 312976 326894 313032
rect 326950 312976 393330 313032
rect 326521 312974 393330 312976
rect 326521 312971 326587 312974
rect 326889 312971 326955 312974
rect 251030 312836 251036 312900
rect 251100 312898 251106 312900
rect 310513 312898 310579 312901
rect 251100 312896 310579 312898
rect 251100 312840 310518 312896
rect 310574 312840 310579 312896
rect 251100 312838 310579 312840
rect 251100 312836 251106 312838
rect 310513 312835 310579 312838
rect 326613 312898 326679 312901
rect 387333 312898 387399 312901
rect 326613 312896 387399 312898
rect 326613 312840 326618 312896
rect 326674 312840 387338 312896
rect 387394 312840 387399 312896
rect 326613 312838 387399 312840
rect 326613 312835 326679 312838
rect 387333 312835 387399 312838
rect 234470 312700 234476 312764
rect 234540 312762 234546 312764
rect 294638 312762 294644 312764
rect 234540 312702 294644 312762
rect 234540 312700 234546 312702
rect 294638 312700 294644 312702
rect 294708 312700 294714 312764
rect 316166 312700 316172 312764
rect 316236 312762 316242 312764
rect 317137 312762 317203 312765
rect 316236 312760 317203 312762
rect 316236 312704 317142 312760
rect 317198 312704 317203 312760
rect 316236 312702 317203 312704
rect 316236 312700 316242 312702
rect 317137 312699 317203 312702
rect 323577 312762 323643 312765
rect 382549 312762 382615 312765
rect 323577 312760 382615 312762
rect 323577 312704 323582 312760
rect 323638 312704 382554 312760
rect 382610 312704 382615 312760
rect 323577 312702 382615 312704
rect 323577 312699 323643 312702
rect 382549 312699 382615 312702
rect 233550 312564 233556 312628
rect 233620 312626 233626 312628
rect 294270 312626 294276 312628
rect 233620 312566 294276 312626
rect 233620 312564 233626 312566
rect 294270 312564 294276 312566
rect 294340 312564 294346 312628
rect 294689 312626 294755 312629
rect 315062 312626 315068 312628
rect 294689 312624 315068 312626
rect 294689 312568 294694 312624
rect 294750 312568 315068 312624
rect 294689 312566 315068 312568
rect 294689 312563 294755 312566
rect 315062 312564 315068 312566
rect 315132 312564 315138 312628
rect 324129 312626 324195 312629
rect 363689 312626 363755 312629
rect 324129 312624 363755 312626
rect 324129 312568 324134 312624
rect 324190 312568 363694 312624
rect 363750 312568 363755 312624
rect 324129 312566 363755 312568
rect 324129 312563 324195 312566
rect 363689 312563 363755 312566
rect 233734 312428 233740 312492
rect 233804 312490 233810 312492
rect 294454 312490 294460 312492
rect 233804 312430 294460 312490
rect 233804 312428 233810 312430
rect 294454 312428 294460 312430
rect 294524 312428 294530 312492
rect 296529 312490 296595 312493
rect 324313 312490 324379 312493
rect 343541 312490 343607 312493
rect 296529 312488 343607 312490
rect 296529 312432 296534 312488
rect 296590 312432 324318 312488
rect 324374 312432 343546 312488
rect 343602 312432 343607 312488
rect 296529 312430 343607 312432
rect 393270 312490 393330 312974
rect 394785 312490 394851 312493
rect 572805 312490 572871 312493
rect 393270 312488 572871 312490
rect 393270 312432 394790 312488
rect 394846 312432 572810 312488
rect 572866 312432 572871 312488
rect 393270 312430 572871 312432
rect 296529 312427 296595 312430
rect 324313 312427 324379 312430
rect 343541 312427 343607 312430
rect 394785 312427 394851 312430
rect 572805 312427 572871 312430
rect 250846 312292 250852 312356
rect 250916 312354 250922 312356
rect 309685 312354 309751 312357
rect 250916 312352 309751 312354
rect 250916 312296 309690 312352
rect 309746 312296 309751 312352
rect 250916 312294 309751 312296
rect 250916 312292 250922 312294
rect 309685 312291 309751 312294
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 583520 311932 584960 312022
rect 232630 311748 232636 311812
rect 232700 311810 232706 311812
rect 271689 311810 271755 311813
rect 292021 311810 292087 311813
rect 392117 311810 392183 311813
rect 232700 311808 292087 311810
rect 232700 311752 271694 311808
rect 271750 311752 292026 311808
rect 292082 311752 292087 311808
rect 232700 311750 292087 311752
rect 232700 311748 232706 311750
rect 271689 311747 271755 311750
rect 292021 311747 292087 311750
rect 321510 311808 392183 311810
rect 321510 311752 392122 311808
rect 392178 311752 392183 311808
rect 321510 311750 392183 311752
rect 270125 311674 270191 311677
rect 317689 311674 317755 311677
rect 321510 311674 321570 311750
rect 392117 311747 392183 311750
rect 270125 311672 321570 311674
rect 270125 311616 270130 311672
rect 270186 311616 317694 311672
rect 317750 311616 321570 311672
rect 270125 311614 321570 311616
rect 324589 311674 324655 311677
rect 325141 311674 325207 311677
rect 324589 311672 393330 311674
rect 324589 311616 324594 311672
rect 324650 311616 325146 311672
rect 325202 311616 393330 311672
rect 324589 311614 393330 311616
rect 270125 311611 270191 311614
rect 317689 311611 317755 311614
rect 324589 311611 324655 311614
rect 325141 311611 325207 311614
rect 259310 311476 259316 311540
rect 259380 311538 259386 311540
rect 318057 311538 318123 311541
rect 259380 311536 318123 311538
rect 259380 311480 318062 311536
rect 318118 311480 318123 311536
rect 259380 311478 318123 311480
rect 259380 311476 259386 311478
rect 318057 311475 318123 311478
rect 326981 311538 327047 311541
rect 392025 311538 392091 311541
rect 326981 311536 392091 311538
rect 326981 311480 326986 311536
rect 327042 311480 392030 311536
rect 392086 311480 392091 311536
rect 326981 311478 392091 311480
rect 326981 311475 327047 311478
rect 392025 311475 392091 311478
rect 231526 311340 231532 311404
rect 231596 311402 231602 311404
rect 291101 311402 291167 311405
rect 231596 311400 291167 311402
rect 231596 311344 291106 311400
rect 291162 311344 291167 311400
rect 231596 311342 291167 311344
rect 231596 311340 231602 311342
rect 291101 311339 291167 311342
rect 316401 311402 316467 311405
rect 375557 311402 375623 311405
rect 316401 311400 375623 311402
rect 316401 311344 316406 311400
rect 316462 311344 375562 311400
rect 375618 311344 375623 311400
rect 316401 311342 375623 311344
rect 316401 311339 316467 311342
rect 375557 311339 375623 311342
rect 231710 311204 231716 311268
rect 231780 311266 231786 311268
rect 290181 311266 290247 311269
rect 231780 311264 290247 311266
rect 231780 311208 290186 311264
rect 290242 311208 290247 311264
rect 231780 311206 290247 311208
rect 231780 311204 231786 311206
rect 290181 311203 290247 311206
rect 291101 311266 291167 311269
rect 325785 311266 325851 311269
rect 326981 311266 327047 311269
rect 291101 311264 327047 311266
rect 291101 311208 291106 311264
rect 291162 311208 325790 311264
rect 325846 311208 326986 311264
rect 327042 311208 327047 311264
rect 291101 311206 327047 311208
rect 291101 311203 291167 311206
rect 325785 311203 325851 311206
rect 326981 311203 327047 311206
rect 231158 311068 231164 311132
rect 231228 311130 231234 311132
rect 231228 311070 277410 311130
rect 231228 311068 231234 311070
rect 277350 310994 277410 311070
rect 291694 311068 291700 311132
rect 291764 311130 291770 311132
rect 313774 311130 313780 311132
rect 291764 311070 313780 311130
rect 291764 311068 291770 311070
rect 313774 311068 313780 311070
rect 313844 311068 313850 311132
rect 322606 311068 322612 311132
rect 322676 311130 322682 311132
rect 328453 311130 328519 311133
rect 382457 311130 382523 311133
rect 322676 311128 382523 311130
rect 322676 311072 328458 311128
rect 328514 311072 382462 311128
rect 382518 311072 382523 311128
rect 322676 311070 382523 311072
rect 393270 311130 393330 311614
rect 394693 311130 394759 311133
rect 556245 311130 556311 311133
rect 393270 311128 556311 311130
rect 393270 311072 394698 311128
rect 394754 311072 556250 311128
rect 556306 311072 556311 311128
rect 393270 311070 556311 311072
rect 322676 311068 322682 311070
rect 328453 311067 328519 311070
rect 382457 311067 382523 311070
rect 394693 311067 394759 311070
rect 556245 311067 556311 311070
rect 291878 310994 291884 310996
rect 277350 310934 291884 310994
rect 291878 310932 291884 310934
rect 291948 310932 291954 310996
rect 318057 310994 318123 310997
rect 330753 310994 330819 310997
rect 318057 310992 330819 310994
rect 318057 310936 318062 310992
rect 318118 310936 330758 310992
rect 330814 310936 330819 310992
rect 318057 310934 330819 310936
rect 318057 310931 318123 310934
rect 330753 310931 330819 310934
rect 283741 310586 283807 310589
rect 295333 310586 295399 310589
rect 283741 310584 295399 310586
rect 283741 310528 283746 310584
rect 283802 310528 295338 310584
rect 295394 310528 295399 310584
rect 283741 310526 295399 310528
rect 283741 310523 283807 310526
rect 295333 310523 295399 310526
rect 316401 310586 316467 310589
rect 317137 310586 317203 310589
rect 316401 310584 317203 310586
rect 316401 310528 316406 310584
rect 316462 310528 317142 310584
rect 317198 310528 317203 310584
rect 316401 310526 317203 310528
rect 316401 310523 316467 310526
rect 317137 310523 317203 310526
rect 227478 310388 227484 310452
rect 227548 310450 227554 310452
rect 257153 310450 257219 310453
rect 257889 310450 257955 310453
rect 227548 310448 257955 310450
rect 227548 310392 257158 310448
rect 257214 310392 257894 310448
rect 257950 310392 257955 310448
rect 227548 310390 257955 310392
rect 227548 310388 227554 310390
rect 257153 310387 257219 310390
rect 257889 310387 257955 310390
rect 259269 310450 259335 310453
rect 289353 310450 289419 310453
rect 259269 310448 289419 310450
rect 259269 310392 259274 310448
rect 259330 310392 289358 310448
rect 289414 310392 289419 310448
rect 259269 310390 289419 310392
rect 259269 310387 259335 310390
rect 289353 310387 289419 310390
rect 290457 310450 290523 310453
rect 297582 310450 297588 310452
rect 290457 310448 297588 310450
rect 290457 310392 290462 310448
rect 290518 310392 297588 310448
rect 290457 310390 297588 310392
rect 290457 310387 290523 310390
rect 297582 310388 297588 310390
rect 297652 310388 297658 310452
rect 326429 310450 326495 310453
rect 326838 310450 326844 310452
rect 326429 310448 326844 310450
rect 326429 310392 326434 310448
rect 326490 310392 326844 310448
rect 326429 310390 326844 310392
rect 326429 310387 326495 310390
rect 326838 310388 326844 310390
rect 326908 310450 326914 310452
rect 387149 310450 387215 310453
rect 326908 310448 387215 310450
rect 326908 310392 387154 310448
rect 387210 310392 387215 310448
rect 326908 310390 387215 310392
rect 326908 310388 326914 310390
rect 387149 310387 387215 310390
rect 239990 310252 239996 310316
rect 240060 310314 240066 310316
rect 270401 310314 270467 310317
rect 299606 310314 299612 310316
rect 240060 310312 299612 310314
rect 240060 310256 270406 310312
rect 270462 310256 299612 310312
rect 240060 310254 299612 310256
rect 240060 310252 240066 310254
rect 270401 310251 270467 310254
rect 299606 310252 299612 310254
rect 299676 310252 299682 310316
rect 321737 310314 321803 310317
rect 322657 310314 322723 310317
rect 380893 310314 380959 310317
rect 321737 310312 380959 310314
rect 321737 310256 321742 310312
rect 321798 310256 322662 310312
rect 322718 310256 380898 310312
rect 380954 310256 380959 310312
rect 321737 310254 380959 310256
rect 321737 310251 321803 310254
rect 322657 310251 322723 310254
rect 380893 310251 380959 310254
rect 226190 310116 226196 310180
rect 226260 310178 226266 310180
rect 260649 310178 260715 310181
rect 286133 310178 286199 310181
rect 226260 310176 286199 310178
rect 226260 310120 260654 310176
rect 260710 310120 286138 310176
rect 286194 310120 286199 310176
rect 226260 310118 286199 310120
rect 226260 310116 226266 310118
rect 260649 310115 260715 310118
rect 286133 310115 286199 310118
rect 324497 310178 324563 310181
rect 325049 310178 325115 310181
rect 383837 310178 383903 310181
rect 324497 310176 383903 310178
rect 324497 310120 324502 310176
rect 324558 310120 325054 310176
rect 325110 310120 383842 310176
rect 383898 310120 383903 310176
rect 324497 310118 383903 310120
rect 324497 310115 324563 310118
rect 325049 310115 325115 310118
rect 383837 310115 383903 310118
rect 241094 309980 241100 310044
rect 241164 310042 241170 310044
rect 300526 310042 300532 310044
rect 241164 309982 300532 310042
rect 241164 309980 241170 309982
rect 300526 309980 300532 309982
rect 300596 309980 300602 310044
rect 320541 310042 320607 310045
rect 321093 310042 321159 310045
rect 375966 310042 375972 310044
rect 320541 310040 375972 310042
rect 320541 309984 320546 310040
rect 320602 309984 321098 310040
rect 321154 309984 375972 310040
rect 320541 309982 375972 309984
rect 320541 309979 320607 309982
rect 321093 309979 321159 309982
rect 375966 309980 375972 309982
rect 376036 309980 376042 310044
rect 231342 309844 231348 309908
rect 231412 309906 231418 309908
rect 291326 309906 291332 309908
rect 231412 309846 291332 309906
rect 231412 309844 231418 309846
rect 291326 309844 291332 309846
rect 291396 309844 291402 309908
rect 230238 309708 230244 309772
rect 230308 309770 230314 309772
rect 290774 309770 290780 309772
rect 230308 309710 290780 309770
rect 230308 309708 230314 309710
rect 290774 309708 290780 309710
rect 290844 309708 290850 309772
rect 291837 309770 291903 309773
rect 299105 309770 299171 309773
rect 291837 309768 299171 309770
rect 291837 309712 291842 309768
rect 291898 309712 299110 309768
rect 299166 309712 299171 309768
rect 291837 309710 299171 309712
rect 291837 309707 291903 309710
rect 299105 309707 299171 309710
rect 228950 309572 228956 309636
rect 229020 309634 229026 309636
rect 259269 309634 259335 309637
rect 287881 309634 287947 309637
rect 229020 309632 259335 309634
rect 229020 309576 259274 309632
rect 259330 309576 259335 309632
rect 229020 309574 259335 309576
rect 229020 309572 229026 309574
rect 259269 309571 259335 309574
rect 277350 309632 287947 309634
rect 277350 309576 287886 309632
rect 287942 309576 287947 309632
rect 277350 309574 287947 309576
rect 257153 309498 257219 309501
rect 277350 309498 277410 309574
rect 287881 309571 287947 309574
rect 257153 309496 277410 309498
rect 257153 309440 257158 309496
rect 257214 309440 277410 309496
rect 257153 309438 277410 309440
rect 288249 309498 288315 309501
rect 328678 309498 328684 309500
rect 288249 309496 328684 309498
rect 288249 309440 288254 309496
rect 288310 309440 328684 309496
rect 288249 309438 328684 309440
rect 257153 309435 257219 309438
rect 288249 309435 288315 309438
rect 328678 309436 328684 309438
rect 328748 309436 328754 309500
rect 285673 309362 285739 309365
rect 324957 309362 325023 309365
rect 285673 309360 325023 309362
rect 285673 309304 285678 309360
rect 285734 309304 324962 309360
rect 325018 309304 325023 309360
rect 285673 309302 325023 309304
rect 285673 309299 285739 309302
rect 324957 309299 325023 309302
rect 284334 309090 284340 309092
rect 267690 309030 284340 309090
rect 206369 308546 206435 308549
rect 263501 308546 263567 308549
rect 267690 308546 267750 309030
rect 284334 309028 284340 309030
rect 284404 309028 284410 309092
rect 323117 309090 323183 309093
rect 323669 309090 323735 309093
rect 323117 309088 323735 309090
rect 323117 309032 323122 309088
rect 323178 309032 323674 309088
rect 323730 309032 323735 309088
rect 323117 309030 323735 309032
rect 323117 309027 323183 309030
rect 323669 309027 323735 309030
rect 324405 308954 324471 308957
rect 325601 308954 325667 308957
rect 384849 308954 384915 308957
rect 324405 308952 384915 308954
rect 324405 308896 324410 308952
rect 324466 308896 325606 308952
rect 325662 308896 384854 308952
rect 384910 308896 384915 308952
rect 324405 308894 384915 308896
rect 324405 308891 324471 308894
rect 325601 308891 325667 308894
rect 384849 308891 384915 308894
rect 301405 308818 301471 308821
rect 358302 308818 358308 308820
rect 301405 308816 358308 308818
rect 301405 308760 301410 308816
rect 301466 308760 358308 308816
rect 301405 308758 358308 308760
rect 301405 308755 301471 308758
rect 358302 308756 358308 308758
rect 358372 308756 358378 308820
rect 269665 308682 269731 308685
rect 319662 308682 319668 308684
rect 269665 308680 319668 308682
rect 269665 308624 269670 308680
rect 269726 308624 319668 308680
rect 269665 308622 319668 308624
rect 269665 308619 269731 308622
rect 319662 308620 319668 308622
rect 319732 308620 319738 308684
rect 323669 308682 323735 308685
rect 383193 308682 383259 308685
rect 323669 308680 383259 308682
rect 323669 308624 323674 308680
rect 323730 308624 383198 308680
rect 383254 308624 383259 308680
rect 323669 308622 383259 308624
rect 323669 308619 323735 308622
rect 383193 308619 383259 308622
rect 206369 308544 267750 308546
rect 206369 308488 206374 308544
rect 206430 308488 263506 308544
rect 263562 308488 267750 308544
rect 206369 308486 267750 308488
rect 206369 308483 206435 308486
rect 263501 308483 263567 308486
rect 270350 308484 270356 308548
rect 270420 308546 270426 308548
rect 327441 308546 327507 308549
rect 270420 308544 327507 308546
rect 270420 308488 327446 308544
rect 327502 308488 327507 308544
rect 270420 308486 327507 308488
rect 270420 308484 270426 308486
rect 327441 308483 327507 308486
rect 218973 308410 219039 308413
rect 301405 308410 301471 308413
rect 218973 308408 301471 308410
rect 218973 308352 218978 308408
rect 219034 308352 301410 308408
rect 301466 308352 301471 308408
rect 218973 308350 301471 308352
rect 218973 308347 219039 308350
rect 301405 308347 301471 308350
rect 314009 308410 314075 308413
rect 356462 308410 356468 308412
rect 314009 308408 356468 308410
rect 314009 308352 314014 308408
rect 314070 308352 356468 308408
rect 314009 308350 356468 308352
rect 314009 308347 314075 308350
rect 356462 308348 356468 308350
rect 356532 308348 356538 308412
rect 210233 307866 210299 307869
rect 313457 307866 313523 307869
rect 314009 307866 314075 307869
rect 210233 307864 302066 307866
rect 210233 307808 210238 307864
rect 210294 307808 302066 307864
rect 210233 307806 302066 307808
rect 210233 307803 210299 307806
rect 267690 307670 277410 307730
rect 204897 307186 204963 307189
rect 266261 307186 266327 307189
rect 267690 307186 267750 307670
rect 277350 307594 277410 307670
rect 281390 307668 281396 307732
rect 281460 307730 281466 307732
rect 283005 307730 283071 307733
rect 281460 307728 283071 307730
rect 281460 307672 283010 307728
rect 283066 307672 283071 307728
rect 281460 307670 283071 307672
rect 302006 307730 302066 307806
rect 313457 307864 314075 307866
rect 313457 307808 313462 307864
rect 313518 307808 314014 307864
rect 314070 307808 314075 307864
rect 313457 307806 314075 307808
rect 313457 307803 313523 307806
rect 314009 307803 314075 307806
rect 302734 307730 302740 307732
rect 302006 307670 302740 307730
rect 281460 307668 281466 307670
rect 283005 307667 283071 307670
rect 302734 307668 302740 307670
rect 302804 307730 302810 307732
rect 362718 307730 362724 307732
rect 302804 307670 362724 307730
rect 302804 307668 302810 307670
rect 362718 307668 362724 307670
rect 362788 307668 362794 307732
rect 282862 307594 282868 307596
rect 277350 307534 282868 307594
rect 282862 307532 282868 307534
rect 282932 307532 282938 307596
rect 322197 307594 322263 307597
rect 322790 307594 322796 307596
rect 322197 307592 322796 307594
rect 322197 307536 322202 307592
rect 322258 307536 322796 307592
rect 322197 307534 322796 307536
rect 322197 307531 322263 307534
rect 322790 307532 322796 307534
rect 322860 307594 322866 307596
rect 380934 307594 380940 307596
rect 322860 307534 380940 307594
rect 322860 307532 322866 307534
rect 380934 307532 380940 307534
rect 381004 307532 381010 307596
rect 304533 307458 304599 307461
rect 312353 307458 312419 307461
rect 369158 307458 369164 307460
rect 304533 307456 369164 307458
rect 304533 307400 304538 307456
rect 304594 307400 312358 307456
rect 312414 307400 369164 307456
rect 304533 307398 369164 307400
rect 304533 307395 304599 307398
rect 312353 307395 312419 307398
rect 369158 307396 369164 307398
rect 369228 307396 369234 307460
rect 312261 307322 312327 307325
rect 312721 307322 312787 307325
rect 359406 307322 359412 307324
rect 312261 307320 359412 307322
rect 312261 307264 312266 307320
rect 312322 307264 312726 307320
rect 312782 307264 359412 307320
rect 312261 307262 359412 307264
rect 312261 307259 312327 307262
rect 312721 307259 312787 307262
rect 359406 307260 359412 307262
rect 359476 307260 359482 307324
rect 204897 307184 267750 307186
rect 204897 307128 204902 307184
rect 204958 307128 266266 307184
rect 266322 307128 267750 307184
rect 204897 307126 267750 307128
rect 204897 307123 204963 307126
rect 266261 307123 266327 307126
rect 271086 307124 271092 307188
rect 271156 307186 271162 307188
rect 330109 307186 330175 307189
rect 271156 307184 330175 307186
rect 271156 307128 330114 307184
rect 330170 307128 330175 307184
rect 271156 307126 330175 307128
rect 271156 307124 271162 307126
rect 330109 307123 330175 307126
rect 220169 307050 220235 307053
rect 313406 307050 313412 307052
rect 220169 307048 313412 307050
rect 220169 306992 220174 307048
rect 220230 306992 313412 307048
rect 220169 306990 313412 306992
rect 220169 306987 220235 306990
rect 313406 306988 313412 306990
rect 313476 307050 313482 307052
rect 314469 307050 314535 307053
rect 313476 307048 314535 307050
rect 313476 306992 314474 307048
rect 314530 306992 314535 307048
rect 313476 306990 314535 306992
rect 313476 306988 313482 306990
rect 314469 306987 314535 306990
rect 314837 307050 314903 307053
rect 315481 307050 315547 307053
rect 345054 307050 345060 307052
rect 314837 307048 345060 307050
rect 314837 306992 314842 307048
rect 314898 306992 315486 307048
rect 315542 306992 345060 307048
rect 314837 306990 345060 306992
rect 314837 306987 314903 306990
rect 315481 306987 315547 306990
rect 345054 306988 345060 306990
rect 345124 306988 345130 307052
rect 327574 306444 327580 306508
rect 327644 306506 327650 306508
rect 571977 306506 572043 306509
rect 327644 306504 572043 306506
rect 327644 306448 571982 306504
rect 572038 306448 572043 306504
rect 327644 306446 572043 306448
rect 327644 306444 327650 306446
rect 571977 306443 572043 306446
rect 306833 306370 306899 306373
rect 307293 306370 307359 306373
rect 364926 306370 364932 306372
rect 306833 306368 364932 306370
rect -960 306234 480 306324
rect 306833 306312 306838 306368
rect 306894 306312 307298 306368
rect 307354 306312 364932 306368
rect 306833 306310 364932 306312
rect 306833 306307 306899 306310
rect 307293 306307 307359 306310
rect 364926 306308 364932 306310
rect 364996 306308 365002 306372
rect 4061 306234 4127 306237
rect -960 306232 4127 306234
rect -960 306176 4066 306232
rect 4122 306176 4127 306232
rect -960 306174 4127 306176
rect -960 306084 480 306174
rect 4061 306171 4127 306174
rect 297725 306234 297791 306237
rect 312169 306234 312235 306237
rect 363454 306234 363460 306236
rect 297725 306232 363460 306234
rect 297725 306176 297730 306232
rect 297786 306176 312174 306232
rect 312230 306176 363460 306232
rect 297725 306174 363460 306176
rect 297725 306171 297791 306174
rect 312169 306171 312235 306174
rect 363454 306172 363460 306174
rect 363524 306172 363530 306236
rect 308673 306098 308739 306101
rect 358118 306098 358124 306100
rect 296670 306096 358124 306098
rect 296670 306040 308678 306096
rect 308734 306040 358124 306096
rect 296670 306038 358124 306040
rect 296253 305962 296319 305965
rect 296670 305962 296730 306038
rect 308673 306035 308739 306038
rect 358118 306036 358124 306038
rect 358188 306036 358194 306100
rect 309501 305962 309567 305965
rect 357934 305962 357940 305964
rect 296253 305960 296730 305962
rect 296253 305904 296258 305960
rect 296314 305904 296730 305960
rect 296253 305902 296730 305904
rect 306330 305960 357940 305962
rect 306330 305904 309506 305960
rect 309562 305904 357940 305960
rect 306330 305902 357940 305904
rect 296253 305899 296319 305902
rect 223982 305764 223988 305828
rect 224052 305826 224058 305828
rect 283925 305826 283991 305829
rect 224052 305824 283991 305826
rect 224052 305768 283930 305824
rect 283986 305768 283991 305824
rect 224052 305766 283991 305768
rect 224052 305764 224058 305766
rect 283925 305763 283991 305766
rect 294873 305826 294939 305829
rect 306330 305826 306390 305902
rect 309501 305899 309567 305902
rect 357934 305900 357940 305902
rect 358004 305900 358010 305964
rect 314745 305826 314811 305829
rect 356646 305826 356652 305828
rect 294873 305824 306390 305826
rect 294873 305768 294878 305824
rect 294934 305768 306390 305824
rect 294873 305766 306390 305768
rect 311850 305824 356652 305826
rect 311850 305768 314750 305824
rect 314806 305768 356652 305824
rect 311850 305766 356652 305768
rect 294873 305763 294939 305766
rect 221641 305690 221707 305693
rect 311850 305690 311910 305766
rect 314745 305763 314811 305766
rect 356646 305764 356652 305766
rect 356716 305764 356722 305828
rect 221641 305688 311910 305690
rect 221641 305632 221646 305688
rect 221702 305632 311910 305688
rect 221641 305630 311910 305632
rect 221641 305627 221707 305630
rect 246982 304948 246988 305012
rect 247052 305010 247058 305012
rect 307109 305010 307175 305013
rect 307661 305010 307727 305013
rect 247052 305008 307727 305010
rect 247052 304952 307114 305008
rect 307170 304952 307666 305008
rect 307722 304952 307727 305008
rect 247052 304950 307727 304952
rect 247052 304948 247058 304950
rect 307109 304947 307175 304950
rect 307661 304947 307727 304950
rect 320582 304948 320588 305012
rect 320652 305010 320658 305012
rect 320909 305010 320975 305013
rect 320652 305008 320975 305010
rect 320652 304952 320914 305008
rect 320970 304952 320975 305008
rect 320652 304950 320975 304952
rect 320652 304948 320658 304950
rect 320909 304947 320975 304950
rect 301446 304812 301452 304876
rect 301516 304874 301522 304876
rect 360694 304874 360700 304876
rect 301516 304814 360700 304874
rect 301516 304812 301522 304814
rect 360694 304812 360700 304814
rect 360764 304812 360770 304876
rect 320449 304738 320515 304741
rect 321277 304738 321343 304741
rect 377305 304738 377371 304741
rect 320449 304736 377371 304738
rect 320449 304680 320454 304736
rect 320510 304680 321282 304736
rect 321338 304680 377310 304736
rect 377366 304680 377371 304736
rect 320449 304678 377371 304680
rect 320449 304675 320515 304678
rect 321277 304675 321343 304678
rect 377305 304675 377371 304678
rect 322381 304602 322447 304605
rect 377254 304602 377260 304604
rect 322381 304600 377260 304602
rect 322381 304544 322386 304600
rect 322442 304544 377260 304600
rect 322381 304542 377260 304544
rect 322381 304539 322447 304542
rect 377254 304540 377260 304542
rect 377324 304540 377330 304604
rect 315665 304330 315731 304333
rect 335537 304330 335603 304333
rect 336457 304330 336523 304333
rect 315665 304328 336523 304330
rect 315665 304272 315670 304328
rect 315726 304272 335542 304328
rect 335598 304272 336462 304328
rect 336518 304272 336523 304328
rect 315665 304270 336523 304272
rect 315665 304267 315731 304270
rect 335537 304267 335603 304270
rect 336457 304267 336523 304270
rect 246798 304132 246804 304196
rect 246868 304194 246874 304196
rect 305494 304194 305500 304196
rect 246868 304134 305500 304194
rect 246868 304132 246874 304134
rect 305494 304132 305500 304134
rect 305564 304194 305570 304196
rect 305564 304134 306390 304194
rect 305564 304132 305570 304134
rect 306330 303650 306390 304134
rect 307753 303650 307819 303653
rect 306330 303648 307819 303650
rect 306330 303592 307758 303648
rect 307814 303592 307819 303648
rect 306330 303590 307819 303592
rect 307753 303587 307819 303590
rect 317505 303516 317571 303517
rect 317454 303514 317460 303516
rect 317414 303454 317460 303514
rect 317524 303512 317571 303516
rect 317566 303456 317571 303512
rect 317454 303452 317460 303454
rect 317524 303452 317571 303456
rect 317505 303451 317571 303452
rect 323945 303514 324011 303517
rect 327257 303514 327323 303517
rect 391933 303514 391999 303517
rect 323945 303512 391999 303514
rect 323945 303456 323950 303512
rect 324006 303456 327262 303512
rect 327318 303456 391938 303512
rect 391994 303456 391999 303512
rect 323945 303454 391999 303456
rect 323945 303451 324011 303454
rect 327257 303451 327323 303454
rect 391933 303451 391999 303454
rect 306649 303378 306715 303381
rect 367318 303378 367324 303380
rect 306649 303376 367324 303378
rect 306649 303320 306654 303376
rect 306710 303320 367324 303376
rect 306649 303318 367324 303320
rect 306649 303315 306715 303318
rect 367318 303316 367324 303318
rect 367388 303316 367394 303380
rect 323025 303242 323091 303245
rect 324037 303242 324103 303245
rect 383009 303242 383075 303245
rect 323025 303240 383075 303242
rect 323025 303184 323030 303240
rect 323086 303184 324042 303240
rect 324098 303184 383014 303240
rect 383070 303184 383075 303240
rect 323025 303182 383075 303184
rect 323025 303179 323091 303182
rect 324037 303179 324103 303182
rect 383009 303179 383075 303182
rect 304758 302908 304764 302972
rect 304828 302970 304834 302972
rect 305361 302970 305427 302973
rect 304828 302968 305427 302970
rect 304828 302912 305366 302968
rect 305422 302912 305427 302968
rect 304828 302910 305427 302912
rect 304828 302908 304834 302910
rect 305361 302907 305427 302910
rect 239438 302772 239444 302836
rect 239508 302834 239514 302836
rect 300025 302834 300091 302837
rect 239508 302832 300091 302834
rect 239508 302776 300030 302832
rect 300086 302776 300091 302832
rect 239508 302774 300091 302776
rect 239508 302772 239514 302774
rect 300025 302771 300091 302774
rect 301865 302834 301931 302837
rect 317505 302834 317571 302837
rect 301865 302832 317571 302834
rect 301865 302776 301870 302832
rect 301926 302776 317510 302832
rect 317566 302776 317571 302832
rect 301865 302774 317571 302776
rect 301865 302771 301931 302774
rect 317505 302771 317571 302774
rect 306649 302290 306715 302293
rect 307109 302290 307175 302293
rect 306649 302288 307175 302290
rect 306649 302232 306654 302288
rect 306710 302232 307114 302288
rect 307170 302232 307175 302288
rect 306649 302230 307175 302232
rect 306649 302227 306715 302230
rect 307109 302227 307175 302230
rect 262121 302154 262187 302157
rect 287329 302154 287395 302157
rect 262121 302152 287395 302154
rect 262121 302096 262126 302152
rect 262182 302096 287334 302152
rect 287390 302096 287395 302152
rect 262121 302094 287395 302096
rect 262121 302091 262187 302094
rect 287329 302091 287395 302094
rect 296161 302154 296227 302157
rect 299197 302154 299263 302157
rect 358854 302154 358860 302156
rect 296161 302152 358860 302154
rect 296161 302096 296166 302152
rect 296222 302096 299202 302152
rect 299258 302096 358860 302152
rect 296161 302094 358860 302096
rect 296161 302091 296227 302094
rect 299197 302091 299263 302094
rect 358854 302092 358860 302094
rect 358924 302092 358930 302156
rect 313038 301956 313044 302020
rect 313108 302018 313114 302020
rect 313108 301958 335370 302018
rect 313108 301956 313114 301958
rect 335310 301746 335370 301958
rect 343633 301746 343699 301749
rect 344921 301746 344987 301749
rect 335310 301744 344987 301746
rect 335310 301688 343638 301744
rect 343694 301688 344926 301744
rect 344982 301688 344987 301744
rect 335310 301686 344987 301688
rect 343633 301683 343699 301686
rect 344921 301683 344987 301686
rect 235206 301548 235212 301612
rect 235276 301610 235282 301612
rect 262121 301610 262187 301613
rect 300761 301612 300827 301613
rect 235276 301608 262187 301610
rect 235276 301552 262126 301608
rect 262182 301552 262187 301608
rect 235276 301550 262187 301552
rect 235276 301548 235282 301550
rect 262121 301547 262187 301550
rect 299606 301548 299612 301612
rect 299676 301610 299682 301612
rect 300710 301610 300716 301612
rect 299676 301550 300716 301610
rect 300780 301610 300827 301612
rect 300780 301608 300908 301610
rect 300822 301552 300908 301608
rect 299676 301548 299682 301550
rect 300710 301548 300716 301550
rect 300780 301550 300908 301552
rect 300780 301548 300827 301550
rect 300761 301547 300827 301548
rect 240910 301412 240916 301476
rect 240980 301474 240986 301476
rect 300894 301474 300900 301476
rect 240980 301414 300900 301474
rect 240980 301412 240986 301414
rect 300894 301412 300900 301414
rect 300964 301412 300970 301476
rect 317454 300732 317460 300796
rect 317524 300794 317530 300796
rect 318374 300794 318380 300796
rect 317524 300734 318380 300794
rect 317524 300732 317530 300734
rect 318374 300732 318380 300734
rect 318444 300794 318450 300796
rect 318701 300794 318767 300797
rect 318444 300792 318767 300794
rect 318444 300736 318706 300792
rect 318762 300736 318767 300792
rect 318444 300734 318767 300736
rect 318444 300732 318450 300734
rect 318701 300731 318767 300734
rect 271270 300188 271276 300252
rect 271340 300250 271346 300252
rect 330702 300250 330708 300252
rect 271340 300190 330708 300250
rect 271340 300188 271346 300190
rect 330702 300188 330708 300190
rect 330772 300188 330778 300252
rect 269614 300052 269620 300116
rect 269684 300114 269690 300116
rect 331765 300114 331831 300117
rect 269684 300112 331831 300114
rect 269684 300056 331770 300112
rect 331826 300056 331831 300112
rect 269684 300054 331831 300056
rect 269684 300052 269690 300054
rect 331765 300051 331831 300054
rect 237782 299372 237788 299436
rect 237852 299434 237858 299436
rect 299381 299434 299447 299437
rect 237852 299432 299447 299434
rect 237852 299376 299386 299432
rect 299442 299376 299447 299432
rect 237852 299374 299447 299376
rect 237852 299372 237858 299374
rect 299381 299371 299447 299374
rect 309726 299372 309732 299436
rect 309796 299434 309802 299436
rect 310329 299434 310395 299437
rect 309796 299432 310395 299434
rect 309796 299376 310334 299432
rect 310390 299376 310395 299432
rect 309796 299374 310395 299376
rect 309796 299372 309802 299374
rect 310329 299371 310395 299374
rect 313774 299372 313780 299436
rect 313844 299434 313850 299436
rect 314510 299434 314516 299436
rect 313844 299374 314516 299434
rect 313844 299372 313850 299374
rect 314510 299372 314516 299374
rect 314580 299434 314586 299436
rect 375414 299434 375420 299436
rect 314580 299374 375420 299434
rect 314580 299372 314586 299374
rect 375414 299372 375420 299374
rect 375484 299372 375490 299436
rect 292430 299236 292436 299300
rect 292500 299298 292506 299300
rect 292849 299298 292915 299301
rect 350574 299298 350580 299300
rect 292500 299296 292915 299298
rect 292500 299240 292854 299296
rect 292910 299240 292915 299296
rect 292500 299238 292915 299240
rect 292500 299236 292506 299238
rect 292849 299235 292915 299238
rect 292990 299238 350580 299298
rect 283925 299026 283991 299029
rect 289997 299026 290063 299029
rect 292990 299026 293050 299238
rect 350574 299236 350580 299238
rect 350644 299236 350650 299300
rect 349286 299162 349292 299164
rect 283925 299024 293050 299026
rect 283925 298968 283930 299024
rect 283986 298968 290002 299024
rect 290058 298968 293050 299024
rect 283925 298966 293050 298968
rect 296670 299102 349292 299162
rect 283925 298963 283991 298966
rect 289997 298963 290063 298966
rect 288801 298890 288867 298893
rect 296670 298890 296730 299102
rect 349286 299100 349292 299102
rect 349356 299100 349362 299164
rect 370446 299026 370452 299028
rect 315990 298966 370452 299026
rect 277350 298888 296730 298890
rect 277350 298832 288806 298888
rect 288862 298832 296730 298888
rect 277350 298830 296730 298832
rect 298921 298890 298987 298893
rect 311617 298890 311683 298893
rect 315990 298890 316050 298966
rect 370446 298964 370452 298966
rect 370516 298964 370522 299028
rect 298921 298888 316050 298890
rect 298921 298832 298926 298888
rect 298982 298832 311622 298888
rect 311678 298832 316050 298888
rect 298921 298830 316050 298832
rect 211981 298754 212047 298757
rect 277350 298754 277410 298830
rect 288801 298827 288867 298830
rect 298921 298827 298987 298830
rect 311617 298827 311683 298830
rect 318190 298828 318196 298892
rect 318260 298890 318266 298892
rect 318701 298890 318767 298893
rect 318260 298888 318767 298890
rect 318260 298832 318706 298888
rect 318762 298832 318767 298888
rect 318260 298830 318767 298832
rect 318260 298828 318266 298830
rect 318701 298827 318767 298830
rect 211981 298752 277410 298754
rect 211981 298696 211986 298752
rect 212042 298696 277410 298752
rect 211981 298694 277410 298696
rect 292849 298754 292915 298757
rect 349102 298754 349108 298756
rect 292849 298752 349108 298754
rect 292849 298696 292854 298752
rect 292910 298696 349108 298752
rect 292849 298694 349108 298696
rect 211981 298691 212047 298694
rect 292849 298691 292915 298694
rect 349102 298692 349108 298694
rect 349172 298692 349178 298756
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 288065 298210 288131 298213
rect 310053 298210 310119 298213
rect 288065 298208 310119 298210
rect 288065 298152 288070 298208
rect 288126 298152 310058 298208
rect 310114 298152 310119 298208
rect 288065 298150 310119 298152
rect 288065 298147 288131 298150
rect 310053 298147 310119 298150
rect 223798 298012 223804 298076
rect 223868 298074 223874 298076
rect 225873 298074 225939 298077
rect 223868 298072 225939 298074
rect 223868 298016 225878 298072
rect 225934 298016 225939 298072
rect 223868 298014 225939 298016
rect 223868 298012 223874 298014
rect 225873 298011 225939 298014
rect 286409 298074 286475 298077
rect 286777 298074 286843 298077
rect 286409 298072 286843 298074
rect 286409 298016 286414 298072
rect 286470 298016 286782 298072
rect 286838 298016 286843 298072
rect 286409 298014 286843 298016
rect 286409 298011 286475 298014
rect 286777 298011 286843 298014
rect 308254 298012 308260 298076
rect 308324 298074 308330 298076
rect 309041 298074 309107 298077
rect 308324 298072 309107 298074
rect 308324 298016 309046 298072
rect 309102 298016 309107 298072
rect 308324 298014 309107 298016
rect 308324 298012 308330 298014
rect 309041 298011 309107 298014
rect 303286 297876 303292 297940
rect 303356 297938 303362 297940
rect 363086 297938 363092 297940
rect 303356 297878 363092 297938
rect 303356 297876 303362 297878
rect 363086 297876 363092 297878
rect 363156 297876 363162 297940
rect 303470 297740 303476 297804
rect 303540 297802 303546 297804
rect 362902 297802 362908 297804
rect 303540 297742 362908 297802
rect 303540 297740 303546 297742
rect 362902 297740 362908 297742
rect 362972 297740 362978 297804
rect 286777 297666 286843 297669
rect 307702 297666 307708 297668
rect 286777 297664 307708 297666
rect 286777 297608 286782 297664
rect 286838 297608 307708 297664
rect 286777 297606 307708 297608
rect 286777 297603 286843 297606
rect 307702 297604 307708 297606
rect 307772 297666 307778 297668
rect 309041 297666 309107 297669
rect 307772 297664 309107 297666
rect 307772 297608 309046 297664
rect 309102 297608 309107 297664
rect 307772 297606 309107 297608
rect 307772 297604 307778 297606
rect 309041 297603 309107 297606
rect 310278 297604 310284 297668
rect 310348 297666 310354 297668
rect 362534 297666 362540 297668
rect 310348 297606 362540 297666
rect 310348 297604 310354 297606
rect 362534 297604 362540 297606
rect 362604 297604 362610 297668
rect 239254 297468 239260 297532
rect 239324 297530 239330 297532
rect 298369 297530 298435 297533
rect 239324 297528 298435 297530
rect 239324 297472 298374 297528
rect 298430 297472 298435 297528
rect 239324 297470 298435 297472
rect 239324 297468 239330 297470
rect 298369 297467 298435 297470
rect 316861 297530 316927 297533
rect 368974 297530 368980 297532
rect 316861 297528 368980 297530
rect 316861 297472 316866 297528
rect 316922 297472 368980 297528
rect 316861 297470 368980 297472
rect 316861 297467 316927 297470
rect 368974 297468 368980 297470
rect 369044 297468 369050 297532
rect 238334 297332 238340 297396
rect 238404 297394 238410 297396
rect 298318 297394 298324 297396
rect 238404 297334 298324 297394
rect 238404 297332 238410 297334
rect 298318 297332 298324 297334
rect 298388 297332 298394 297396
rect 289445 297258 289511 297261
rect 318701 297258 318767 297261
rect 289445 297256 318767 297258
rect 289445 297200 289450 297256
rect 289506 297200 318706 297256
rect 318762 297200 318767 297256
rect 289445 297198 318767 297200
rect 289445 297195 289511 297198
rect 318701 297195 318767 297198
rect 285397 297122 285463 297125
rect 307569 297122 307635 297125
rect 308949 297122 309015 297125
rect 285397 297120 309015 297122
rect 285397 297064 285402 297120
rect 285458 297064 307574 297120
rect 307630 297064 308954 297120
rect 309010 297064 309015 297120
rect 285397 297062 309015 297064
rect 285397 297059 285463 297062
rect 307569 297059 307635 297062
rect 308949 297059 309015 297062
rect 286409 296986 286475 296989
rect 346342 296986 346348 296988
rect 286409 296984 346348 296986
rect 286409 296928 286414 296984
rect 286470 296928 346348 296984
rect 286409 296926 346348 296928
rect 286409 296923 286475 296926
rect 346342 296924 346348 296926
rect 346412 296924 346418 296988
rect 315297 296850 315363 296853
rect 316861 296850 316927 296853
rect 315297 296848 316927 296850
rect 315297 296792 315302 296848
rect 315358 296792 316866 296848
rect 316922 296792 316927 296848
rect 315297 296790 316927 296792
rect 315297 296787 315363 296790
rect 316861 296787 316927 296790
rect 227294 296516 227300 296580
rect 227364 296578 227370 296580
rect 285622 296578 285628 296580
rect 227364 296518 285628 296578
rect 227364 296516 227370 296518
rect 285622 296516 285628 296518
rect 285692 296516 285698 296580
rect 225822 296380 225828 296444
rect 225892 296442 225898 296444
rect 285806 296442 285812 296444
rect 225892 296382 285812 296442
rect 225892 296380 225898 296382
rect 285806 296380 285812 296382
rect 285876 296380 285882 296444
rect 227110 296244 227116 296308
rect 227180 296306 227186 296308
rect 288341 296306 288407 296309
rect 227180 296304 288407 296306
rect 227180 296248 288346 296304
rect 288402 296248 288407 296304
rect 227180 296246 288407 296248
rect 227180 296244 227186 296246
rect 288341 296243 288407 296246
rect 228766 296108 228772 296172
rect 228836 296170 228842 296172
rect 288709 296170 288775 296173
rect 228836 296168 288775 296170
rect 228836 296112 288714 296168
rect 288770 296112 288775 296168
rect 228836 296110 288775 296112
rect 228836 296108 228842 296110
rect 288709 296107 288775 296110
rect 226926 295972 226932 296036
rect 226996 296034 227002 296036
rect 287605 296034 287671 296037
rect 226996 296032 287671 296034
rect 226996 295976 287610 296032
rect 287666 295976 287671 296032
rect 226996 295974 287671 295976
rect 226996 295972 227002 295974
rect 287605 295971 287671 295974
rect 229686 295156 229692 295220
rect 229756 295218 229762 295220
rect 288750 295218 288756 295220
rect 229756 295158 288756 295218
rect 229756 295156 229762 295158
rect 288750 295156 288756 295158
rect 288820 295156 288826 295220
rect 292205 295218 292271 295221
rect 354438 295218 354444 295220
rect 292205 295216 354444 295218
rect 292205 295160 292210 295216
rect 292266 295160 354444 295216
rect 292205 295158 354444 295160
rect 292205 295155 292271 295158
rect 354438 295156 354444 295158
rect 354508 295156 354514 295220
rect 223062 295020 223068 295084
rect 223132 295082 223138 295084
rect 284017 295082 284083 295085
rect 223132 295080 284083 295082
rect 223132 295024 284022 295080
rect 284078 295024 284083 295080
rect 223132 295022 284083 295024
rect 223132 295020 223138 295022
rect 284017 295019 284083 295022
rect 290733 295082 290799 295085
rect 352046 295082 352052 295084
rect 290733 295080 352052 295082
rect 290733 295024 290738 295080
rect 290794 295024 352052 295080
rect 290733 295022 352052 295024
rect 290733 295019 290799 295022
rect 352046 295020 352052 295022
rect 352116 295020 352122 295084
rect 227846 294884 227852 294948
rect 227916 294946 227922 294948
rect 288617 294946 288683 294949
rect 227916 294944 288683 294946
rect 227916 294888 288622 294944
rect 288678 294888 288683 294944
rect 227916 294886 288683 294888
rect 227916 294884 227922 294886
rect 288617 294883 288683 294886
rect 229870 294748 229876 294812
rect 229940 294810 229946 294812
rect 289905 294810 289971 294813
rect 229940 294808 289971 294810
rect 229940 294752 289910 294808
rect 289966 294752 289971 294808
rect 229940 294750 289971 294752
rect 229940 294748 229946 294750
rect 289905 294747 289971 294750
rect 290549 294810 290615 294813
rect 317638 294810 317644 294812
rect 290549 294808 317644 294810
rect 290549 294752 290554 294808
rect 290610 294752 317644 294808
rect 290549 294750 317644 294752
rect 290549 294747 290615 294750
rect 317638 294748 317644 294750
rect 317708 294748 317714 294812
rect 223614 294612 223620 294676
rect 223684 294674 223690 294676
rect 230197 294674 230263 294677
rect 223684 294672 230263 294674
rect 223684 294616 230202 294672
rect 230258 294616 230263 294672
rect 223684 294614 230263 294616
rect 223684 294612 223690 294614
rect 230197 294611 230263 294614
rect 231301 294674 231367 294677
rect 289721 294674 289787 294677
rect 347814 294674 347820 294676
rect 231301 294672 347820 294674
rect 231301 294616 231306 294672
rect 231362 294616 289726 294672
rect 289782 294616 347820 294672
rect 231301 294614 347820 294616
rect 231301 294611 231367 294614
rect 289721 294611 289787 294614
rect 347814 294612 347820 294614
rect 347884 294612 347890 294676
rect 230054 294476 230060 294540
rect 230124 294538 230130 294540
rect 291009 294538 291075 294541
rect 230124 294536 291075 294538
rect 230124 294480 291014 294536
rect 291070 294480 291075 294536
rect 230124 294478 291075 294480
rect 230124 294476 230130 294478
rect 291009 294475 291075 294478
rect 228214 294340 228220 294404
rect 228284 294402 228290 294404
rect 231301 294402 231367 294405
rect 291142 294402 291148 294404
rect 228284 294400 231367 294402
rect 228284 294344 231306 294400
rect 231362 294344 231367 294400
rect 228284 294342 231367 294344
rect 228284 294340 228290 294342
rect 231301 294339 231367 294342
rect 238710 294342 291148 294402
rect 232446 294204 232452 294268
rect 232516 294266 232522 294268
rect 238710 294266 238770 294342
rect 291142 294340 291148 294342
rect 291212 294340 291218 294404
rect 232516 294206 238770 294266
rect 232516 294204 232522 294206
rect 245142 293524 245148 293588
rect 245212 293586 245218 293588
rect 304022 293586 304028 293588
rect 245212 293526 304028 293586
rect 245212 293524 245218 293526
rect 304022 293524 304028 293526
rect 304092 293524 304098 293588
rect 238150 293388 238156 293452
rect 238220 293450 238226 293452
rect 298134 293450 298140 293452
rect 238220 293390 298140 293450
rect 238220 293388 238226 293390
rect 298134 293388 298140 293390
rect 298204 293388 298210 293452
rect -960 293178 480 293268
rect 236862 293252 236868 293316
rect 236932 293314 236938 293316
rect 297909 293314 297975 293317
rect 236932 293312 297975 293314
rect 236932 293256 297914 293312
rect 297970 293256 297975 293312
rect 236932 293254 297975 293256
rect 236932 293252 236938 293254
rect 297909 293251 297975 293254
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 239070 293116 239076 293180
rect 239140 293178 239146 293180
rect 300577 293178 300643 293181
rect 239140 293176 300643 293178
rect 239140 293120 300582 293176
rect 300638 293120 300643 293176
rect 239140 293118 300643 293120
rect 239140 293116 239146 293118
rect 300577 293115 300643 293118
rect 224217 292906 224283 292909
rect 224677 292906 224743 292909
rect 219390 292904 224743 292906
rect 219390 292848 224222 292904
rect 224278 292848 224682 292904
rect 224738 292848 224743 292904
rect 219390 292846 224743 292848
rect 164325 292770 164391 292773
rect 219390 292770 219450 292846
rect 224217 292843 224283 292846
rect 224677 292843 224743 292846
rect 164325 292768 219450 292770
rect 164325 292712 164330 292768
rect 164386 292712 219450 292768
rect 164325 292710 219450 292712
rect 164325 292707 164391 292710
rect 162761 292634 162827 292637
rect 225781 292634 225847 292637
rect 162761 292632 225847 292634
rect 162761 292576 162766 292632
rect 162822 292576 225786 292632
rect 225842 292576 225847 292632
rect 162761 292574 225847 292576
rect 162761 292571 162827 292574
rect 225781 292571 225847 292574
rect 218697 292226 218763 292229
rect 252553 292226 252619 292229
rect 218697 292224 252619 292226
rect 218697 292168 218702 292224
rect 218758 292168 252558 292224
rect 252614 292168 252619 292224
rect 218697 292166 252619 292168
rect 218697 292163 218763 292166
rect 252553 292163 252619 292166
rect 251173 292090 251239 292093
rect 261477 292090 261543 292093
rect 251173 292088 261543 292090
rect 251173 292032 251178 292088
rect 251234 292032 261482 292088
rect 261538 292032 261543 292088
rect 251173 292030 261543 292032
rect 251173 292027 251239 292030
rect 261477 292027 261543 292030
rect 220261 291954 220327 291957
rect 224585 291954 224651 291957
rect 220261 291952 224651 291954
rect 220261 291896 220266 291952
rect 220322 291896 224590 291952
rect 224646 291896 224651 291952
rect 220261 291894 224651 291896
rect 220261 291891 220327 291894
rect 224585 291891 224651 291894
rect 250805 291954 250871 291957
rect 267181 291954 267247 291957
rect 250805 291952 267247 291954
rect 250805 291896 250810 291952
rect 250866 291896 267186 291952
rect 267242 291896 267247 291952
rect 250805 291894 267247 291896
rect 250805 291891 250871 291894
rect 267181 291891 267247 291894
rect 217133 291818 217199 291821
rect 229461 291818 229527 291821
rect 229921 291818 229987 291821
rect 217133 291816 229987 291818
rect 217133 291760 217138 291816
rect 217194 291760 229466 291816
rect 229522 291760 229926 291816
rect 229982 291760 229987 291816
rect 217133 291758 229987 291760
rect 217133 291755 217199 291758
rect 229461 291755 229527 291758
rect 229921 291755 229987 291758
rect 246614 291756 246620 291820
rect 246684 291818 246690 291820
rect 306598 291818 306604 291820
rect 246684 291758 306604 291818
rect 246684 291756 246690 291758
rect 306598 291756 306604 291758
rect 306668 291756 306674 291820
rect 220721 291682 220787 291685
rect 224401 291682 224467 291685
rect 220721 291680 224467 291682
rect 220721 291624 220726 291680
rect 220782 291624 224406 291680
rect 224462 291624 224467 291680
rect 220721 291622 224467 291624
rect 220721 291619 220787 291622
rect 224401 291619 224467 291622
rect 224585 291682 224651 291685
rect 249149 291682 249215 291685
rect 224585 291680 249215 291682
rect 224585 291624 224590 291680
rect 224646 291624 249154 291680
rect 249210 291624 249215 291680
rect 224585 291622 249215 291624
rect 224585 291619 224651 291622
rect 249149 291619 249215 291622
rect 220118 291484 220124 291548
rect 220188 291546 220194 291548
rect 250621 291546 250687 291549
rect 220188 291544 250687 291546
rect 220188 291488 250626 291544
rect 250682 291488 250687 291544
rect 220188 291486 250687 291488
rect 220188 291484 220194 291486
rect 250621 291483 250687 291486
rect 219934 291348 219940 291412
rect 220004 291410 220010 291412
rect 251541 291410 251607 291413
rect 251909 291410 251975 291413
rect 220004 291408 251975 291410
rect 220004 291352 251546 291408
rect 251602 291352 251914 291408
rect 251970 291352 251975 291408
rect 220004 291350 251975 291352
rect 220004 291348 220010 291350
rect 251541 291347 251607 291350
rect 251909 291347 251975 291350
rect 221222 291212 221228 291276
rect 221292 291274 221298 291276
rect 225505 291274 225571 291277
rect 226149 291274 226215 291277
rect 221292 291272 226215 291274
rect 221292 291216 225510 291272
rect 225566 291216 226154 291272
rect 226210 291216 226215 291272
rect 221292 291214 226215 291216
rect 221292 291212 221298 291214
rect 225505 291211 225571 291214
rect 226149 291211 226215 291214
rect 190637 290730 190703 290733
rect 248321 290730 248387 290733
rect 190637 290728 248387 290730
rect 190637 290672 190642 290728
rect 190698 290672 248326 290728
rect 248382 290672 248387 290728
rect 190637 290670 248387 290672
rect 190637 290667 190703 290670
rect 248321 290667 248387 290670
rect 249701 290730 249767 290733
rect 279366 290730 279372 290732
rect 249701 290728 279372 290730
rect 249701 290672 249706 290728
rect 249762 290672 279372 290728
rect 249701 290670 279372 290672
rect 249701 290667 249767 290670
rect 279366 290668 279372 290670
rect 279436 290668 279442 290732
rect 192201 290594 192267 290597
rect 252829 290594 252895 290597
rect 192201 290592 252895 290594
rect 192201 290536 192206 290592
rect 192262 290536 252834 290592
rect 252890 290536 252895 290592
rect 192201 290534 252895 290536
rect 192201 290531 192267 290534
rect 252829 290531 252895 290534
rect 192017 290458 192083 290461
rect 251909 290458 251975 290461
rect 267089 290458 267155 290461
rect 192017 290456 251834 290458
rect 192017 290400 192022 290456
rect 192078 290400 251834 290456
rect 192017 290398 251834 290400
rect 192017 290395 192083 290398
rect 251774 290325 251834 290398
rect 251909 290456 267155 290458
rect 251909 290400 251914 290456
rect 251970 290400 267094 290456
rect 267150 290400 267155 290456
rect 251909 290398 267155 290400
rect 251909 290395 251975 290398
rect 267089 290395 267155 290398
rect 220721 290324 220787 290325
rect 220670 290322 220676 290324
rect 220594 290262 220676 290322
rect 220740 290322 220787 290324
rect 227621 290322 227687 290325
rect 220740 290320 227687 290322
rect 220782 290264 227626 290320
rect 227682 290264 227687 290320
rect 220670 290260 220676 290262
rect 220740 290262 227687 290264
rect 220740 290260 220787 290262
rect 220721 290259 220787 290260
rect 227621 290259 227687 290262
rect 245694 290260 245700 290324
rect 245764 290322 245770 290324
rect 251173 290322 251239 290325
rect 251774 290322 251883 290325
rect 252093 290322 252159 290325
rect 245764 290320 251239 290322
rect 245764 290264 251178 290320
rect 251234 290264 251239 290320
rect 245764 290262 251239 290264
rect 251690 290320 252159 290322
rect 251690 290264 251822 290320
rect 251878 290264 252098 290320
rect 252154 290264 252159 290320
rect 251690 290262 252159 290264
rect 245764 290260 245770 290262
rect 251173 290259 251239 290262
rect 251817 290259 251883 290262
rect 252093 290259 252159 290262
rect 221825 290186 221891 290189
rect 249701 290186 249767 290189
rect 221825 290184 249767 290186
rect 221825 290128 221830 290184
rect 221886 290128 249706 290184
rect 249762 290128 249767 290184
rect 221825 290126 249767 290128
rect 221825 290123 221891 290126
rect 249701 290123 249767 290126
rect 191833 290050 191899 290053
rect 251725 290050 251791 290053
rect 191833 290048 251791 290050
rect 191833 289992 191838 290048
rect 191894 289992 251730 290048
rect 251786 289992 251791 290048
rect 191833 289990 251791 289992
rect 191833 289987 191899 289990
rect 251725 289987 251791 289990
rect 190453 289914 190519 289917
rect 245694 289914 245700 289916
rect 190453 289912 245700 289914
rect 190453 289856 190458 289912
rect 190514 289856 245700 289912
rect 190453 289854 245700 289856
rect 190453 289851 190519 289854
rect 245694 289852 245700 289854
rect 245764 289852 245770 289916
rect 247677 289914 247743 289917
rect 245886 289912 247743 289914
rect 245886 289856 247682 289912
rect 247738 289856 247743 289912
rect 245886 289854 247743 289856
rect 245886 289778 245946 289854
rect 247677 289851 247743 289854
rect 248965 289778 249031 289781
rect 219390 289718 245946 289778
rect 246070 289776 249031 289778
rect 246070 289720 248970 289776
rect 249026 289720 249031 289776
rect 246070 289718 249031 289720
rect 189809 289506 189875 289509
rect 219390 289506 219450 289718
rect 225454 289580 225460 289644
rect 225524 289642 225530 289644
rect 226057 289642 226123 289645
rect 246070 289642 246130 289718
rect 248965 289715 249031 289718
rect 246389 289644 246455 289645
rect 246389 289642 246436 289644
rect 225524 289640 226123 289642
rect 225524 289584 226062 289640
rect 226118 289584 226123 289640
rect 225524 289582 226123 289584
rect 225524 289580 225530 289582
rect 226057 289579 226123 289582
rect 233926 289582 246130 289642
rect 246344 289640 246436 289642
rect 246344 289584 246394 289640
rect 246344 289582 246436 289584
rect 189809 289504 219450 289506
rect 189809 289448 189814 289504
rect 189870 289448 219450 289504
rect 189809 289446 219450 289448
rect 189809 289443 189875 289446
rect 187785 289234 187851 289237
rect 233926 289234 233986 289582
rect 246389 289580 246436 289582
rect 246500 289580 246506 289644
rect 247166 289580 247172 289644
rect 247236 289642 247242 289644
rect 248137 289642 248203 289645
rect 247236 289640 248203 289642
rect 247236 289584 248142 289640
rect 248198 289584 248203 289640
rect 247236 289582 248203 289584
rect 247236 289580 247242 289582
rect 246389 289579 246455 289580
rect 248137 289579 248203 289582
rect 253890 289582 258090 289642
rect 246246 289444 246252 289508
rect 246316 289506 246322 289508
rect 247033 289506 247099 289509
rect 246316 289504 247099 289506
rect 246316 289448 247038 289504
rect 247094 289448 247099 289504
rect 246316 289446 247099 289448
rect 246316 289444 246322 289446
rect 247033 289443 247099 289446
rect 247534 289444 247540 289508
rect 247604 289506 247610 289508
rect 248045 289506 248111 289509
rect 247604 289504 248111 289506
rect 247604 289448 248050 289504
rect 248106 289448 248111 289504
rect 247604 289446 248111 289448
rect 247604 289444 247610 289446
rect 248045 289443 248111 289446
rect 251766 289444 251772 289508
rect 251836 289506 251842 289508
rect 252461 289506 252527 289509
rect 251836 289504 252527 289506
rect 251836 289448 252466 289504
rect 252522 289448 252527 289504
rect 251836 289446 252527 289448
rect 251836 289444 251842 289446
rect 252461 289443 252527 289446
rect 252686 289444 252692 289508
rect 252756 289506 252762 289508
rect 253657 289506 253723 289509
rect 252756 289504 253723 289506
rect 252756 289448 253662 289504
rect 253718 289448 253723 289504
rect 252756 289446 253723 289448
rect 252756 289444 252762 289446
rect 253657 289443 253723 289446
rect 237925 289370 237991 289373
rect 187785 289232 233986 289234
rect 187785 289176 187790 289232
rect 187846 289176 233986 289232
rect 187785 289174 233986 289176
rect 234570 289368 237991 289370
rect 234570 289312 237930 289368
rect 237986 289312 237991 289368
rect 234570 289310 237991 289312
rect 187785 289171 187851 289174
rect 176745 289098 176811 289101
rect 234570 289098 234630 289310
rect 237925 289307 237991 289310
rect 240726 289308 240732 289372
rect 240796 289370 240802 289372
rect 241237 289370 241303 289373
rect 240796 289368 241303 289370
rect 240796 289312 241242 289368
rect 241298 289312 241303 289368
rect 240796 289310 241303 289312
rect 240796 289308 240802 289310
rect 241237 289307 241303 289310
rect 244038 289308 244044 289372
rect 244108 289370 244114 289372
rect 253890 289370 253950 289582
rect 244108 289310 253950 289370
rect 258030 289370 258090 289582
rect 303245 289370 303311 289373
rect 258030 289368 303311 289370
rect 258030 289312 303250 289368
rect 303306 289312 303311 289368
rect 258030 289310 303311 289312
rect 244108 289308 244114 289310
rect 303245 289307 303311 289310
rect 176745 289096 234630 289098
rect 176745 289040 176750 289096
rect 176806 289040 234630 289096
rect 176745 289038 234630 289040
rect 176745 289035 176811 289038
rect 244958 289036 244964 289100
rect 245028 289098 245034 289100
rect 306097 289098 306163 289101
rect 245028 289096 306163 289098
rect 245028 289040 306102 289096
rect 306158 289040 306163 289096
rect 245028 289038 306163 289040
rect 245028 289036 245034 289038
rect 306097 289035 306163 289038
rect 186405 288690 186471 288693
rect 246430 288690 246436 288692
rect 186405 288688 246436 288690
rect 186405 288632 186410 288688
rect 186466 288632 246436 288688
rect 186405 288630 246436 288632
rect 186405 288627 186471 288630
rect 246430 288628 246436 288630
rect 246500 288690 246506 288692
rect 272701 288690 272767 288693
rect 246500 288688 272767 288690
rect 246500 288632 272706 288688
rect 272762 288632 272767 288688
rect 246500 288630 272767 288632
rect 246500 288628 246506 288630
rect 272701 288627 272767 288630
rect 180885 288554 180951 288557
rect 240726 288554 240732 288556
rect 180885 288552 240732 288554
rect 180885 288496 180890 288552
rect 180946 288496 240732 288552
rect 180885 288494 240732 288496
rect 180885 288491 180951 288494
rect 240726 288492 240732 288494
rect 240796 288554 240802 288556
rect 267457 288554 267523 288557
rect 240796 288552 267523 288554
rect 240796 288496 267462 288552
rect 267518 288496 267523 288552
rect 240796 288494 267523 288496
rect 240796 288492 240802 288494
rect 267457 288491 267523 288494
rect 250662 287676 250668 287740
rect 250732 287738 250738 287740
rect 311709 287738 311775 287741
rect 250732 287736 311775 287738
rect 250732 287680 311714 287736
rect 311770 287680 311775 287736
rect 250732 287678 311775 287680
rect 250732 287676 250738 287678
rect 311709 287675 311775 287678
rect 257102 286316 257108 286380
rect 257172 286378 257178 286380
rect 316534 286378 316540 286380
rect 257172 286318 316540 286378
rect 257172 286316 257178 286318
rect 316534 286316 316540 286318
rect 316604 286316 316610 286380
rect 583520 285276 584960 285516
rect 220905 285154 220971 285157
rect 221549 285154 221615 285157
rect 220905 285152 221615 285154
rect 220905 285096 220910 285152
rect 220966 285096 221554 285152
rect 221610 285096 221615 285152
rect 220905 285094 221615 285096
rect 220905 285091 220971 285094
rect 221549 285091 221615 285094
rect 165705 282162 165771 282165
rect 221222 282162 221228 282164
rect 165705 282160 221228 282162
rect 165705 282104 165710 282160
rect 165766 282104 221228 282160
rect 165705 282102 221228 282104
rect 165705 282099 165771 282102
rect 221222 282100 221228 282102
rect 221292 282100 221298 282164
rect -960 279972 480 280212
rect 220905 276722 220971 276725
rect 222009 276722 222075 276725
rect 220905 276720 222075 276722
rect 220905 276664 220910 276720
rect 220966 276664 222014 276720
rect 222070 276664 222075 276720
rect 220905 276662 222075 276664
rect 220905 276659 220971 276662
rect 222009 276659 222075 276662
rect 190545 272506 190611 272509
rect 220118 272506 220124 272508
rect 190545 272504 220124 272506
rect 190545 272448 190550 272504
rect 190606 272448 220124 272504
rect 190545 272446 220124 272448
rect 190545 272443 190611 272446
rect 220118 272444 220124 272446
rect 220188 272444 220194 272508
rect 580625 272234 580691 272237
rect 583520 272234 584960 272324
rect 580625 272232 584960 272234
rect 580625 272176 580630 272232
rect 580686 272176 584960 272232
rect 580625 272174 584960 272176
rect 580625 272171 580691 272174
rect 583520 272084 584960 272174
rect 265014 271084 265020 271148
rect 265084 271146 265090 271148
rect 325141 271146 325207 271149
rect 265084 271144 325207 271146
rect 265084 271088 325146 271144
rect 325202 271088 325207 271144
rect 265084 271086 325207 271088
rect 265084 271084 265090 271086
rect 325141 271083 325207 271086
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 256918 267140 256924 267204
rect 256988 267202 256994 267204
rect 316350 267202 316356 267204
rect 256988 267142 316356 267202
rect 256988 267140 256994 267142
rect 316350 267140 316356 267142
rect 316420 267140 316426 267204
rect 255814 267004 255820 267068
rect 255884 267066 255890 267068
rect 316769 267066 316835 267069
rect 255884 267064 316835 267066
rect 255884 267008 316774 267064
rect 316830 267008 316835 267064
rect 255884 267006 316835 267008
rect 255884 267004 255890 267006
rect 316769 267003 316835 267006
rect 256366 265508 256372 265572
rect 256436 265570 256442 265572
rect 314878 265570 314884 265572
rect 256436 265510 314884 265570
rect 256436 265508 256442 265510
rect 314878 265508 314884 265510
rect 314948 265508 314954 265572
rect 260598 264284 260604 264348
rect 260668 264346 260674 264348
rect 318926 264346 318932 264348
rect 260668 264286 318932 264346
rect 260668 264284 260674 264286
rect 318926 264284 318932 264286
rect 318996 264284 319002 264348
rect 267590 264148 267596 264212
rect 267660 264210 267666 264212
rect 326705 264210 326771 264213
rect 267660 264208 326771 264210
rect 267660 264152 326710 264208
rect 326766 264152 326771 264208
rect 267660 264150 326771 264152
rect 267660 264148 267666 264150
rect 326705 264147 326771 264150
rect 259126 260068 259132 260132
rect 259196 260130 259202 260132
rect 318149 260130 318215 260133
rect 259196 260128 318215 260130
rect 259196 260072 318154 260128
rect 318210 260072 318215 260128
rect 259196 260070 318215 260072
rect 259196 260068 259202 260070
rect 318149 260067 318215 260070
rect 580533 258906 580599 258909
rect 583520 258906 584960 258996
rect 580533 258904 584960 258906
rect 580533 258848 580538 258904
rect 580594 258848 584960 258904
rect 580533 258846 584960 258848
rect 580533 258843 580599 258846
rect 262806 258708 262812 258772
rect 262876 258770 262882 258772
rect 322381 258770 322447 258773
rect 262876 258768 322447 258770
rect 262876 258712 322386 258768
rect 322442 258712 322447 258768
rect 583520 258756 584960 258846
rect 262876 258710 322447 258712
rect 262876 258708 262882 258710
rect 322381 258707 322447 258710
rect 270217 257546 270283 257549
rect 287094 257546 287100 257548
rect 270217 257544 287100 257546
rect 270217 257488 270222 257544
rect 270278 257488 287100 257544
rect 270217 257486 287100 257488
rect 270217 257483 270283 257486
rect 287094 257484 287100 257486
rect 287164 257484 287170 257548
rect 256182 257348 256188 257412
rect 256252 257410 256258 257412
rect 315573 257410 315639 257413
rect 256252 257408 315639 257410
rect 256252 257352 315578 257408
rect 315634 257352 315639 257408
rect 256252 257350 315639 257352
rect 256252 257348 256258 257350
rect 315573 257347 315639 257350
rect 267549 257274 267615 257277
rect 327073 257274 327139 257277
rect 267549 257272 327139 257274
rect 267549 257216 267554 257272
rect 267610 257216 327078 257272
rect 327134 257216 327139 257272
rect 267549 257214 327139 257216
rect 267549 257211 267615 257214
rect 327073 257211 327139 257214
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 260966 253132 260972 253196
rect 261036 253194 261042 253196
rect 321001 253194 321067 253197
rect 261036 253192 321067 253194
rect 261036 253136 321006 253192
rect 321062 253136 321067 253192
rect 261036 253134 321067 253136
rect 261036 253132 261042 253134
rect 321001 253131 321067 253134
rect 268009 250610 268075 250613
rect 326521 250610 326587 250613
rect 268009 250608 326587 250610
rect 268009 250552 268014 250608
rect 268070 250552 326526 250608
rect 326582 250552 326587 250608
rect 268009 250550 326587 250552
rect 268009 250547 268075 250550
rect 326521 250547 326587 250550
rect 264462 250412 264468 250476
rect 264532 250474 264538 250476
rect 325049 250474 325115 250477
rect 264532 250472 325115 250474
rect 264532 250416 325054 250472
rect 325110 250416 325115 250472
rect 264532 250414 325115 250416
rect 264532 250412 264538 250414
rect 325049 250411 325115 250414
rect 267549 249250 267615 249253
rect 327022 249250 327028 249252
rect 267549 249248 327028 249250
rect 267549 249192 267554 249248
rect 267610 249192 327028 249248
rect 267549 249190 327028 249192
rect 267549 249187 267615 249190
rect 327022 249188 327028 249190
rect 327092 249188 327098 249252
rect 262254 249052 262260 249116
rect 262324 249114 262330 249116
rect 322197 249114 322263 249117
rect 262324 249112 322263 249114
rect 262324 249056 322202 249112
rect 322258 249056 322263 249112
rect 262324 249054 322263 249056
rect 262324 249052 262330 249054
rect 322197 249051 322263 249054
rect 268837 247890 268903 247893
rect 290590 247890 290596 247892
rect 268837 247888 290596 247890
rect 268837 247832 268842 247888
rect 268898 247832 290596 247888
rect 268837 247830 290596 247832
rect 268837 247827 268903 247830
rect 290590 247828 290596 247830
rect 290660 247828 290666 247892
rect 269113 247754 269179 247757
rect 326429 247754 326495 247757
rect 269113 247752 326495 247754
rect 269113 247696 269118 247752
rect 269174 247696 326434 247752
rect 326490 247696 326495 247752
rect 269113 247694 326495 247696
rect 269113 247691 269179 247694
rect 326429 247691 326495 247694
rect 267733 247618 267799 247621
rect 323669 247618 323735 247621
rect 267733 247616 323735 247618
rect 267733 247560 267738 247616
rect 267794 247560 323674 247616
rect 323730 247560 323735 247616
rect 267733 247558 323735 247560
rect 267733 247555 267799 247558
rect 323669 247555 323735 247558
rect 270401 246394 270467 246397
rect 325693 246394 325759 246397
rect 270401 246392 325759 246394
rect 270401 246336 270406 246392
rect 270462 246336 325698 246392
rect 325754 246336 325759 246392
rect 270401 246334 325759 246336
rect 270401 246331 270467 246334
rect 325693 246331 325759 246334
rect 262438 246196 262444 246260
rect 262508 246258 262514 246260
rect 323577 246258 323643 246261
rect 262508 246256 323643 246258
rect 262508 246200 323582 246256
rect 323638 246200 323643 246256
rect 262508 246198 323643 246200
rect 262508 246196 262514 246198
rect 323577 246195 323643 246198
rect 579613 245578 579679 245581
rect 583520 245578 584960 245668
rect 579613 245576 584960 245578
rect 579613 245520 579618 245576
rect 579674 245520 584960 245576
rect 579613 245518 584960 245520
rect 579613 245515 579679 245518
rect 270769 245442 270835 245445
rect 289302 245442 289308 245444
rect 270769 245440 289308 245442
rect 270769 245384 270774 245440
rect 270830 245384 289308 245440
rect 270769 245382 289308 245384
rect 270769 245379 270835 245382
rect 289302 245380 289308 245382
rect 289372 245380 289378 245444
rect 583520 245428 584960 245518
rect 281165 245306 281231 245309
rect 305126 245306 305132 245308
rect 281165 245304 305132 245306
rect 281165 245248 281170 245304
rect 281226 245248 305132 245304
rect 281165 245246 305132 245248
rect 281165 245243 281231 245246
rect 305126 245244 305132 245246
rect 305196 245244 305202 245308
rect 277117 245170 277183 245173
rect 316166 245170 316172 245172
rect 277117 245168 316172 245170
rect 277117 245112 277122 245168
rect 277178 245112 316172 245168
rect 277117 245110 316172 245112
rect 277117 245107 277183 245110
rect 316166 245108 316172 245110
rect 316236 245108 316242 245172
rect 264830 244972 264836 245036
rect 264900 245034 264906 245036
rect 325509 245034 325575 245037
rect 264900 245032 325575 245034
rect 264900 244976 325514 245032
rect 325570 244976 325575 245032
rect 264900 244974 325575 244976
rect 264900 244972 264906 244974
rect 325509 244971 325575 244974
rect 266118 244836 266124 244900
rect 266188 244898 266194 244900
rect 326337 244898 326403 244901
rect 266188 244896 326403 244898
rect 266188 244840 326342 244896
rect 326398 244840 326403 244896
rect 266188 244838 326403 244840
rect 266188 244836 266194 244838
rect 326337 244835 326403 244838
rect 260782 243748 260788 243812
rect 260852 243810 260858 243812
rect 272149 243810 272215 243813
rect 278773 243810 278839 243813
rect 322974 243810 322980 243812
rect 260852 243808 276030 243810
rect 260852 243752 272154 243808
rect 272210 243752 276030 243808
rect 260852 243750 276030 243752
rect 260852 243748 260858 243750
rect 272149 243747 272215 243750
rect 275970 243674 276030 243750
rect 278773 243808 322980 243810
rect 278773 243752 278778 243808
rect 278834 243752 322980 243808
rect 278773 243750 322980 243752
rect 278773 243747 278839 243750
rect 322974 243748 322980 243750
rect 323044 243748 323050 243812
rect 320950 243674 320956 243676
rect 275970 243614 320956 243674
rect 320950 243612 320956 243614
rect 321020 243612 321026 243676
rect 265014 243476 265020 243540
rect 265084 243538 265090 243540
rect 324446 243538 324452 243540
rect 265084 243478 324452 243538
rect 265084 243476 265090 243478
rect 324446 243476 324452 243478
rect 324516 243476 324522 243540
rect 267406 243068 267412 243132
rect 267476 243130 267482 243132
rect 268653 243130 268719 243133
rect 267476 243128 268719 243130
rect 267476 243072 268658 243128
rect 268714 243072 268719 243128
rect 267476 243070 268719 243072
rect 267476 243068 267482 243070
rect 268653 243067 268719 243070
rect 268653 242994 268719 242997
rect 278773 242994 278839 242997
rect 268653 242992 278839 242994
rect 268653 242936 268658 242992
rect 268714 242936 278778 242992
rect 278834 242936 278839 242992
rect 268653 242934 278839 242936
rect 268653 242931 268719 242934
rect 278773 242931 278839 242934
rect 265934 242796 265940 242860
rect 266004 242858 266010 242860
rect 286225 242858 286291 242861
rect 266004 242856 286291 242858
rect 266004 242800 286230 242856
rect 286286 242800 286291 242856
rect 266004 242798 286291 242800
rect 266004 242796 266010 242798
rect 286225 242795 286291 242798
rect 263726 242660 263732 242724
rect 263796 242722 263802 242724
rect 285489 242722 285555 242725
rect 263796 242720 285555 242722
rect 263796 242664 285494 242720
rect 285550 242664 285555 242720
rect 263796 242662 285555 242664
rect 263796 242660 263802 242662
rect 285489 242659 285555 242662
rect 272333 242586 272399 242589
rect 320081 242586 320147 242589
rect 272333 242584 320147 242586
rect 272333 242528 272338 242584
rect 272394 242528 320086 242584
rect 320142 242528 320147 242584
rect 272333 242526 320147 242528
rect 272333 242523 272399 242526
rect 320081 242523 320147 242526
rect 259862 242388 259868 242452
rect 259932 242450 259938 242452
rect 319529 242450 319595 242453
rect 259932 242448 319595 242450
rect 259932 242392 319534 242448
rect 319590 242392 319595 242448
rect 259932 242390 319595 242392
rect 259932 242388 259938 242390
rect 319529 242387 319595 242390
rect 257286 242252 257292 242316
rect 257356 242314 257362 242316
rect 316902 242314 316908 242316
rect 257356 242254 316908 242314
rect 257356 242252 257362 242254
rect 316902 242252 316908 242254
rect 316972 242252 316978 242316
rect 190729 242178 190795 242181
rect 219934 242178 219940 242180
rect 190729 242176 219940 242178
rect 190729 242120 190734 242176
rect 190790 242120 219940 242176
rect 190729 242118 219940 242120
rect 190729 242115 190795 242118
rect 219934 242116 219940 242118
rect 220004 242116 220010 242180
rect 260230 242116 260236 242180
rect 260300 242178 260306 242180
rect 320909 242178 320975 242181
rect 260300 242176 320975 242178
rect 260300 242120 320914 242176
rect 320970 242120 320975 242176
rect 260300 242118 320975 242120
rect 260300 242116 260306 242118
rect 320909 242115 320975 242118
rect 264646 241980 264652 242044
rect 264716 242042 264722 242044
rect 264716 241982 266370 242042
rect 264716 241980 264722 241982
rect 266310 241906 266370 241982
rect 273846 241980 273852 242044
rect 273916 242042 273922 242044
rect 274541 242042 274607 242045
rect 273916 242040 274607 242042
rect 273916 241984 274546 242040
rect 274602 241984 274607 242040
rect 273916 241982 274607 241984
rect 273916 241980 273922 241982
rect 274541 241979 274607 241982
rect 274541 241906 274607 241909
rect 266310 241904 274607 241906
rect 266310 241848 274546 241904
rect 274602 241848 274607 241904
rect 266310 241846 274607 241848
rect 274541 241843 274607 241846
rect 158621 241770 158687 241773
rect 222878 241770 222884 241772
rect 158621 241768 222884 241770
rect 158621 241712 158626 241768
rect 158682 241712 222884 241768
rect 158621 241710 222884 241712
rect 158621 241707 158687 241710
rect 222878 241708 222884 241710
rect 222948 241708 222954 241772
rect 226006 241708 226012 241772
rect 226076 241770 226082 241772
rect 237966 241770 237972 241772
rect 226076 241710 237972 241770
rect 226076 241708 226082 241710
rect 237966 241708 237972 241710
rect 238036 241708 238042 241772
rect 265750 241708 265756 241772
rect 265820 241770 265826 241772
rect 273846 241770 273852 241772
rect 265820 241710 273852 241770
rect 265820 241708 265826 241710
rect 273846 241708 273852 241710
rect 273916 241708 273922 241772
rect 151721 241634 151787 241637
rect 228214 241634 228220 241636
rect 151721 241632 228220 241634
rect 151721 241576 151726 241632
rect 151782 241576 228220 241632
rect 151721 241574 228220 241576
rect 151721 241571 151787 241574
rect 228214 241572 228220 241574
rect 228284 241572 228290 241636
rect 231894 241572 231900 241636
rect 231964 241634 231970 241636
rect 231964 241574 233204 241634
rect 231964 241572 231970 241574
rect 159909 241498 159975 241501
rect 217409 241498 217475 241501
rect 232998 241498 233004 241500
rect 159909 241496 233004 241498
rect 159909 241440 159914 241496
rect 159970 241440 217414 241496
rect 217470 241440 233004 241496
rect 159909 241438 233004 241440
rect 159909 241435 159975 241438
rect 217409 241435 217475 241438
rect 232998 241436 233004 241438
rect 233068 241436 233074 241500
rect 207933 241362 207999 241365
rect 219341 241362 219407 241365
rect 200070 241360 219407 241362
rect 200070 241304 207938 241360
rect 207994 241304 219346 241360
rect 219402 241304 219407 241360
rect 200070 241302 219407 241304
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 155861 241090 155927 241093
rect 200070 241090 200130 241302
rect 207933 241299 207999 241302
rect 219341 241299 219407 241302
rect 232078 241300 232084 241364
rect 232148 241362 232154 241364
rect 232630 241362 232636 241364
rect 232148 241302 232636 241362
rect 232148 241300 232154 241302
rect 232630 241300 232636 241302
rect 232700 241300 232706 241364
rect 233144 241362 233204 241574
rect 234838 241572 234844 241636
rect 234908 241634 234914 241636
rect 234908 241574 252570 241634
rect 234908 241572 234914 241574
rect 252510 241498 252570 241574
rect 256550 241572 256556 241636
rect 256620 241634 256626 241636
rect 270217 241634 270283 241637
rect 256620 241632 270283 241634
rect 256620 241576 270222 241632
rect 270278 241576 270283 241632
rect 256620 241574 270283 241576
rect 256620 241572 256626 241574
rect 270217 241571 270283 241574
rect 271689 241634 271755 241637
rect 271822 241634 271828 241636
rect 271689 241632 271828 241634
rect 271689 241576 271694 241632
rect 271750 241576 271828 241632
rect 271689 241574 271828 241576
rect 271689 241571 271755 241574
rect 271822 241572 271828 241574
rect 271892 241572 271898 241636
rect 288382 241498 288388 241500
rect 252510 241438 288388 241498
rect 288382 241436 288388 241438
rect 288452 241436 288458 241500
rect 283373 241362 283439 241365
rect 233144 241360 283439 241362
rect 233144 241304 283378 241360
rect 283434 241304 283439 241360
rect 233144 241302 283439 241304
rect 283373 241299 283439 241302
rect 226742 241164 226748 241228
rect 226812 241226 226818 241228
rect 285581 241226 285647 241229
rect 226812 241224 285647 241226
rect 226812 241168 285586 241224
rect 285642 241168 285647 241224
rect 226812 241166 285647 241168
rect 226812 241164 226818 241166
rect 285581 241163 285647 241166
rect 155861 241088 200130 241090
rect 155861 241032 155866 241088
rect 155922 241032 200130 241088
rect 155861 241030 200130 241032
rect 155861 241027 155927 241030
rect 225270 241028 225276 241092
rect 225340 241090 225346 241092
rect 284293 241090 284359 241093
rect 225340 241088 284359 241090
rect 225340 241032 284298 241088
rect 284354 241032 284359 241088
rect 225340 241030 284359 241032
rect 225340 241028 225346 241030
rect 284293 241027 284359 241030
rect 154481 240954 154547 240957
rect 210601 240954 210667 240957
rect 220353 240954 220419 240957
rect 154481 240952 220419 240954
rect 154481 240896 154486 240952
rect 154542 240896 210606 240952
rect 210662 240896 220358 240952
rect 220414 240896 220419 240952
rect 154481 240894 220419 240896
rect 154481 240891 154547 240894
rect 210601 240891 210667 240894
rect 220353 240891 220419 240894
rect 221273 240954 221339 240957
rect 232630 240954 232636 240956
rect 221273 240952 232636 240954
rect 221273 240896 221278 240952
rect 221334 240896 232636 240952
rect 221273 240894 232636 240896
rect 221273 240891 221339 240894
rect 232630 240892 232636 240894
rect 232700 240892 232706 240956
rect 233366 240892 233372 240956
rect 233436 240954 233442 240956
rect 292614 240954 292620 240956
rect 233436 240894 292620 240954
rect 233436 240892 233442 240894
rect 292614 240892 292620 240894
rect 292684 240892 292690 240956
rect 218973 240818 219039 240821
rect 242014 240818 242020 240820
rect 218973 240816 242020 240818
rect 218973 240760 218978 240816
rect 219034 240760 242020 240816
rect 218973 240758 242020 240760
rect 218973 240755 219039 240758
rect 242014 240756 242020 240758
rect 242084 240756 242090 240820
rect 270033 240818 270099 240821
rect 252510 240816 270099 240818
rect 252510 240760 270038 240816
rect 270094 240760 270099 240816
rect 252510 240758 270099 240760
rect 220813 240682 220879 240685
rect 233918 240682 233924 240684
rect 220813 240680 233924 240682
rect 220813 240624 220818 240680
rect 220874 240624 233924 240680
rect 220813 240622 233924 240624
rect 220813 240619 220879 240622
rect 233918 240620 233924 240622
rect 233988 240620 233994 240684
rect 234286 240620 234292 240684
rect 234356 240682 234362 240684
rect 252510 240682 252570 240758
rect 270033 240755 270099 240758
rect 270861 240818 270927 240821
rect 328494 240818 328500 240820
rect 270861 240816 328500 240818
rect 270861 240760 270866 240816
rect 270922 240760 328500 240816
rect 270861 240758 328500 240760
rect 270861 240755 270927 240758
rect 328494 240756 328500 240758
rect 328564 240756 328570 240820
rect 234356 240622 252570 240682
rect 234356 240620 234362 240622
rect 265382 240620 265388 240684
rect 265452 240682 265458 240684
rect 269205 240682 269271 240685
rect 265452 240680 269271 240682
rect 265452 240624 269210 240680
rect 269266 240624 269271 240680
rect 265452 240622 269271 240624
rect 265452 240620 265458 240622
rect 269205 240619 269271 240622
rect 235022 240546 235028 240548
rect 215250 240486 235028 240546
rect 213269 240410 213335 240413
rect 215250 240410 215310 240486
rect 235022 240484 235028 240486
rect 235092 240484 235098 240548
rect 213269 240408 215310 240410
rect 213269 240352 213274 240408
rect 213330 240352 215310 240408
rect 213269 240350 215310 240352
rect 217133 240410 217199 240413
rect 218973 240410 219039 240413
rect 217133 240408 219039 240410
rect 217133 240352 217138 240408
rect 217194 240352 218978 240408
rect 219034 240352 219039 240408
rect 217133 240350 219039 240352
rect 213269 240347 213335 240350
rect 217133 240347 217199 240350
rect 218973 240347 219039 240350
rect 222694 240348 222700 240412
rect 222764 240410 222770 240412
rect 223430 240410 223436 240412
rect 222764 240350 223436 240410
rect 222764 240348 222770 240350
rect 223430 240348 223436 240350
rect 223500 240348 223506 240412
rect 232630 240348 232636 240412
rect 232700 240410 232706 240412
rect 238886 240410 238892 240412
rect 232700 240350 238892 240410
rect 232700 240348 232706 240350
rect 238886 240348 238892 240350
rect 238956 240348 238962 240412
rect 268101 240410 268167 240413
rect 258950 240408 268167 240410
rect 258950 240352 268106 240408
rect 268162 240352 268167 240408
rect 258950 240350 268167 240352
rect 154205 240274 154271 240277
rect 225270 240274 225276 240276
rect 154205 240272 225276 240274
rect 154205 240216 154210 240272
rect 154266 240216 225276 240272
rect 154205 240214 225276 240216
rect 154205 240211 154271 240214
rect 225270 240212 225276 240214
rect 225340 240212 225346 240276
rect 228030 240212 228036 240276
rect 228100 240274 228106 240276
rect 235206 240274 235212 240276
rect 228100 240214 235212 240274
rect 228100 240212 228106 240214
rect 235206 240212 235212 240214
rect 235276 240212 235282 240276
rect 236310 240212 236316 240276
rect 236380 240274 236386 240276
rect 236862 240274 236868 240276
rect 236380 240214 236868 240274
rect 236380 240212 236386 240214
rect 236862 240212 236868 240214
rect 236932 240212 236938 240276
rect 237330 240214 241530 240274
rect 213453 240138 213519 240141
rect 221089 240138 221155 240141
rect 213453 240136 221155 240138
rect 213453 240080 213458 240136
rect 213514 240080 221094 240136
rect 221150 240080 221155 240136
rect 213453 240078 221155 240080
rect 213453 240075 213519 240078
rect 221089 240075 221155 240078
rect 222009 240138 222075 240141
rect 222009 240136 225752 240138
rect 222009 240080 222014 240136
rect 222070 240080 225752 240136
rect 222009 240078 225752 240080
rect 222009 240075 222075 240078
rect 222975 239900 223041 239903
rect 222975 239898 223084 239900
rect 211061 239866 211127 239869
rect 222975 239866 222980 239898
rect 211061 239864 222980 239866
rect 211061 239808 211066 239864
rect 211122 239842 222980 239864
rect 223036 239842 223084 239898
rect 211122 239808 223084 239842
rect 211061 239806 223084 239808
rect 223665 239866 223731 239869
rect 225275 239868 225341 239869
rect 225459 239868 225525 239869
rect 224718 239866 224724 239868
rect 223665 239864 224724 239866
rect 223665 239808 223670 239864
rect 223726 239808 224724 239864
rect 223665 239806 224724 239808
rect 211061 239803 211127 239806
rect 223665 239803 223731 239806
rect 224718 239804 224724 239806
rect 224788 239804 224794 239868
rect 225270 239866 225276 239868
rect 225184 239806 225276 239866
rect 225270 239804 225276 239806
rect 225340 239804 225346 239868
rect 225454 239804 225460 239868
rect 225524 239866 225530 239868
rect 225524 239806 225616 239866
rect 225524 239804 225530 239806
rect 225275 239803 225341 239804
rect 225459 239803 225525 239804
rect 225692 239733 225752 240078
rect 226374 240076 226380 240140
rect 226444 240138 226450 240140
rect 237330 240138 237390 240214
rect 226444 240078 237390 240138
rect 241470 240138 241530 240214
rect 258950 240138 259010 240350
rect 268101 240347 268167 240350
rect 269205 240410 269271 240413
rect 269614 240410 269620 240412
rect 269205 240408 269620 240410
rect 269205 240352 269210 240408
rect 269266 240352 269620 240408
rect 269205 240350 269620 240352
rect 269205 240347 269271 240350
rect 269614 240348 269620 240350
rect 269684 240348 269690 240412
rect 281533 240274 281599 240277
rect 282453 240274 282519 240277
rect 241470 240078 247004 240138
rect 226444 240076 226450 240078
rect 225822 239940 225828 240004
rect 225892 240002 225898 240004
rect 225892 239942 226304 240002
rect 225892 239940 225898 239942
rect 226244 239869 226304 239942
rect 227846 239940 227852 240004
rect 227916 240002 227922 240004
rect 230422 240002 230428 240004
rect 227916 239942 230428 240002
rect 227916 239940 227922 239942
rect 228958 239869 229018 239942
rect 230422 239940 230428 239942
rect 230492 239940 230498 240004
rect 233734 239940 233740 240004
rect 233804 240002 233810 240004
rect 233804 239942 234354 240002
rect 233804 239940 233810 239942
rect 234294 239869 234354 239942
rect 226244 239864 226353 239869
rect 226244 239808 226292 239864
rect 226348 239808 226353 239864
rect 226244 239806 226353 239808
rect 226287 239803 226353 239806
rect 226425 239866 226491 239869
rect 227115 239868 227181 239869
rect 226558 239866 226564 239868
rect 226425 239864 226564 239866
rect 226425 239808 226430 239864
rect 226486 239808 226564 239864
rect 226425 239806 226564 239808
rect 226425 239803 226491 239806
rect 226558 239804 226564 239806
rect 226628 239804 226634 239868
rect 227110 239866 227116 239868
rect 227024 239806 227116 239866
rect 227110 239804 227116 239806
rect 227180 239804 227186 239868
rect 227575 239866 227641 239869
rect 227989 239868 228055 239869
rect 227846 239866 227852 239868
rect 227575 239864 227852 239866
rect 227575 239808 227580 239864
rect 227636 239808 227852 239864
rect 227575 239806 227852 239808
rect 227115 239803 227181 239804
rect 227575 239803 227641 239806
rect 227846 239804 227852 239806
rect 227916 239804 227922 239868
rect 227989 239864 228036 239868
rect 228100 239866 228106 239868
rect 227989 239808 227994 239864
rect 227989 239804 228036 239808
rect 228100 239806 228146 239866
rect 228955 239864 229021 239869
rect 228955 239808 228960 239864
rect 229016 239808 229021 239864
rect 228100 239804 228106 239806
rect 227989 239803 228055 239804
rect 228955 239803 229021 239808
rect 229134 239804 229140 239868
rect 229204 239866 229210 239868
rect 229691 239866 229757 239869
rect 229204 239864 229757 239866
rect 229204 239808 229696 239864
rect 229752 239808 229757 239864
rect 229204 239806 229757 239808
rect 229204 239804 229210 239806
rect 229691 239803 229757 239806
rect 229870 239804 229876 239868
rect 229940 239866 229946 239868
rect 230335 239866 230401 239869
rect 230611 239868 230677 239869
rect 230606 239866 230612 239868
rect 229940 239864 230401 239866
rect 229940 239808 230340 239864
rect 230396 239808 230401 239864
rect 229940 239806 230401 239808
rect 230520 239806 230612 239866
rect 229940 239804 229946 239806
rect 230335 239803 230401 239806
rect 230606 239804 230612 239806
rect 230676 239804 230682 239868
rect 230887 239866 230953 239869
rect 231710 239866 231716 239868
rect 230887 239864 231716 239866
rect 230887 239808 230892 239864
rect 230948 239808 231716 239864
rect 230887 239806 231716 239808
rect 230611 239803 230677 239804
rect 230887 239803 230953 239806
rect 231710 239804 231716 239806
rect 231780 239804 231786 239868
rect 231991 239866 232057 239869
rect 232446 239866 232452 239868
rect 231991 239864 232452 239866
rect 231991 239808 231996 239864
rect 232052 239808 232452 239864
rect 231991 239806 232452 239808
rect 231991 239803 232057 239806
rect 232446 239804 232452 239806
rect 232516 239804 232522 239868
rect 232814 239804 232820 239868
rect 232884 239866 232890 239868
rect 233187 239866 233253 239869
rect 232884 239864 233253 239866
rect 232884 239808 233192 239864
rect 233248 239808 233253 239864
rect 232884 239806 233253 239808
rect 232884 239804 232890 239806
rect 233187 239803 233253 239806
rect 233366 239804 233372 239868
rect 233436 239866 233442 239868
rect 233509 239866 233575 239869
rect 233436 239864 233575 239866
rect 233436 239808 233514 239864
rect 233570 239808 233575 239864
rect 233436 239806 233575 239808
rect 233436 239804 233442 239806
rect 233509 239803 233575 239806
rect 233785 239866 233851 239869
rect 234102 239866 234108 239868
rect 233785 239864 234108 239866
rect 233785 239808 233790 239864
rect 233846 239808 234108 239864
rect 233785 239806 234108 239808
rect 233785 239803 233851 239806
rect 234102 239804 234108 239806
rect 234172 239804 234178 239868
rect 234245 239864 234354 239869
rect 234245 239808 234250 239864
rect 234306 239808 234354 239864
rect 234475 239898 234541 239903
rect 236775 239900 236841 239903
rect 234475 239842 234480 239898
rect 234536 239866 234541 239898
rect 236732 239898 236841 239900
rect 234654 239866 234660 239868
rect 234536 239842 234660 239866
rect 234475 239837 234660 239842
rect 234245 239806 234354 239808
rect 234478 239806 234660 239837
rect 234245 239803 234311 239806
rect 234654 239804 234660 239806
rect 234724 239804 234730 239868
rect 236310 239804 236316 239868
rect 236380 239866 236386 239868
rect 236732 239866 236780 239898
rect 236380 239842 236780 239866
rect 236836 239842 236841 239898
rect 238707 239898 238773 239903
rect 237603 239868 237669 239869
rect 237598 239866 237604 239868
rect 236380 239837 236841 239842
rect 236380 239806 236792 239837
rect 237512 239806 237604 239866
rect 236380 239804 236386 239806
rect 237598 239804 237604 239806
rect 237668 239804 237674 239868
rect 237782 239804 237788 239868
rect 237852 239866 237858 239868
rect 238707 239866 238712 239898
rect 237852 239842 238712 239866
rect 238768 239842 238773 239898
rect 239259 239900 239325 239903
rect 239627 239900 239693 239903
rect 240271 239900 240337 239903
rect 240639 239900 240705 239903
rect 242111 239900 242177 239903
rect 239259 239898 239382 239900
rect 239259 239868 239264 239898
rect 239320 239868 239382 239898
rect 239627 239898 239750 239900
rect 239627 239868 239632 239898
rect 239688 239868 239750 239898
rect 237852 239837 238773 239842
rect 237852 239806 238770 239837
rect 237852 239804 237858 239806
rect 237603 239803 237669 239804
rect 230890 239733 230950 239803
rect 238710 239733 238770 239806
rect 239254 239804 239260 239868
rect 239324 239840 239382 239868
rect 239324 239804 239330 239840
rect 239622 239804 239628 239868
rect 239692 239840 239750 239868
rect 240136 239898 240337 239900
rect 240136 239842 240276 239898
rect 240332 239842 240337 239898
rect 240596 239898 240705 239900
rect 240596 239868 240644 239898
rect 240136 239840 240337 239842
rect 239692 239804 239698 239840
rect 239811 239764 239877 239767
rect 239811 239762 239934 239764
rect 222745 239730 222811 239733
rect 223389 239732 223455 239733
rect 223246 239730 223252 239732
rect 222745 239728 223252 239730
rect 222745 239672 222750 239728
rect 222806 239672 223252 239728
rect 222745 239670 223252 239672
rect 222745 239667 222811 239670
rect 223246 239668 223252 239670
rect 223316 239668 223322 239732
rect 223389 239728 223436 239732
rect 223500 239730 223506 239732
rect 223389 239672 223394 239728
rect 223389 239668 223436 239672
rect 223500 239670 223546 239730
rect 223500 239668 223506 239670
rect 223798 239668 223804 239732
rect 223868 239730 223874 239732
rect 223941 239730 224007 239733
rect 223868 239728 224007 239730
rect 223868 239672 223946 239728
rect 224002 239672 224007 239728
rect 223868 239670 224007 239672
rect 223868 239668 223874 239670
rect 223389 239667 223455 239668
rect 223941 239667 224007 239670
rect 224166 239668 224172 239732
rect 224236 239730 224242 239732
rect 224953 239730 225019 239733
rect 224236 239728 225019 239730
rect 224236 239672 224958 239728
rect 225014 239672 225019 239728
rect 224236 239670 225019 239672
rect 224236 239668 224242 239670
rect 224953 239667 225019 239670
rect 225689 239728 225755 239733
rect 225689 239672 225694 239728
rect 225750 239672 225755 239728
rect 225689 239667 225755 239672
rect 226885 239730 226951 239733
rect 227161 239730 227227 239733
rect 226885 239728 227227 239730
rect 226885 239672 226890 239728
rect 226946 239672 227166 239728
rect 227222 239672 227227 239728
rect 226885 239670 227227 239672
rect 226885 239667 226951 239670
rect 227161 239667 227227 239670
rect 227989 239730 228055 239733
rect 228725 239732 228791 239733
rect 228725 239730 228772 239732
rect 227989 239728 228772 239730
rect 227989 239672 227994 239728
rect 228050 239672 228730 239728
rect 227989 239670 228772 239672
rect 227989 239667 228055 239670
rect 228725 239668 228772 239670
rect 228836 239668 228842 239732
rect 230151 239730 230217 239733
rect 230606 239730 230612 239732
rect 230151 239728 230612 239730
rect 230151 239672 230156 239728
rect 230212 239672 230612 239728
rect 230151 239670 230612 239672
rect 228725 239667 228791 239668
rect 230151 239667 230217 239670
rect 230606 239668 230612 239670
rect 230676 239668 230682 239732
rect 230890 239728 230999 239733
rect 231117 239732 231183 239733
rect 231393 239732 231459 239733
rect 231117 239730 231164 239732
rect 230890 239672 230938 239728
rect 230994 239672 230999 239728
rect 230890 239670 230999 239672
rect 231072 239728 231164 239730
rect 231072 239672 231122 239728
rect 231072 239670 231164 239672
rect 230933 239667 230999 239670
rect 231117 239668 231164 239670
rect 231228 239668 231234 239732
rect 231342 239668 231348 239732
rect 231412 239730 231459 239732
rect 231853 239730 231919 239733
rect 232078 239730 232084 239732
rect 231412 239728 231504 239730
rect 231454 239672 231504 239728
rect 231412 239670 231504 239672
rect 231853 239728 232084 239730
rect 231853 239672 231858 239728
rect 231914 239672 232084 239728
rect 231853 239670 232084 239672
rect 231412 239668 231459 239670
rect 231117 239667 231183 239668
rect 231393 239667 231459 239668
rect 231853 239667 231919 239670
rect 232078 239668 232084 239670
rect 232148 239668 232154 239732
rect 232262 239668 232268 239732
rect 232332 239730 232338 239732
rect 233233 239730 233299 239733
rect 232332 239728 233299 239730
rect 232332 239672 233238 239728
rect 233294 239672 233299 239728
rect 232332 239670 233299 239672
rect 232332 239668 232338 239670
rect 233233 239667 233299 239670
rect 233601 239730 233667 239733
rect 233877 239730 233943 239733
rect 234286 239730 234292 239732
rect 233601 239728 234292 239730
rect 233601 239672 233606 239728
rect 233662 239672 233882 239728
rect 233938 239672 234292 239728
rect 233601 239670 234292 239672
rect 233601 239667 233667 239670
rect 233877 239667 233943 239670
rect 234286 239668 234292 239670
rect 234356 239668 234362 239732
rect 234470 239668 234476 239732
rect 234540 239730 234546 239732
rect 234613 239730 234679 239733
rect 234540 239728 234679 239730
rect 234540 239672 234618 239728
rect 234674 239672 234679 239728
rect 234540 239670 234679 239672
rect 234540 239668 234546 239670
rect 234613 239667 234679 239670
rect 235022 239668 235028 239732
rect 235092 239730 235098 239732
rect 236177 239730 236243 239733
rect 235092 239728 236243 239730
rect 235092 239672 236182 239728
rect 236238 239672 236243 239728
rect 235092 239670 236243 239672
rect 235092 239668 235098 239670
rect 236177 239667 236243 239670
rect 236678 239668 236684 239732
rect 236748 239730 236754 239732
rect 236821 239730 236887 239733
rect 236748 239728 236887 239730
rect 236748 239672 236826 239728
rect 236882 239672 236887 239728
rect 236748 239670 236887 239672
rect 236748 239668 236754 239670
rect 236821 239667 236887 239670
rect 237419 239730 237485 239733
rect 237649 239730 237715 239733
rect 237419 239728 237715 239730
rect 237419 239672 237424 239728
rect 237480 239672 237654 239728
rect 237710 239672 237715 239728
rect 237419 239670 237715 239672
rect 237419 239667 237485 239670
rect 237649 239667 237715 239670
rect 238201 239730 238267 239733
rect 238385 239732 238451 239733
rect 238334 239730 238340 239732
rect 238201 239728 238340 239730
rect 238404 239728 238451 239732
rect 238201 239672 238206 239728
rect 238262 239672 238340 239728
rect 238446 239672 238451 239728
rect 238201 239670 238340 239672
rect 238201 239667 238267 239670
rect 238334 239668 238340 239670
rect 238404 239668 238451 239672
rect 238385 239667 238451 239668
rect 238661 239728 238770 239733
rect 238661 239672 238666 239728
rect 238722 239672 238770 239728
rect 238661 239670 238770 239672
rect 238661 239667 238727 239670
rect 238886 239668 238892 239732
rect 238956 239730 238962 239732
rect 239213 239730 239279 239733
rect 239811 239732 239816 239762
rect 239872 239732 239934 239762
rect 238956 239728 239279 239730
rect 238956 239672 239218 239728
rect 239274 239672 239279 239728
rect 238956 239670 239279 239672
rect 238956 239668 238962 239670
rect 239213 239667 239279 239670
rect 239806 239668 239812 239732
rect 239876 239704 239934 239732
rect 240136 239730 240196 239840
rect 240271 239837 240337 239840
rect 240542 239804 240548 239868
rect 240612 239842 240644 239868
rect 240700 239866 240705 239898
rect 242068 239898 242177 239900
rect 241094 239866 241100 239868
rect 240700 239842 241100 239866
rect 240612 239806 241100 239842
rect 240612 239804 240618 239806
rect 241094 239804 241100 239806
rect 241164 239804 241170 239868
rect 241559 239866 241625 239869
rect 242068 239868 242116 239898
rect 241286 239864 241625 239866
rect 241286 239808 241564 239864
rect 241620 239808 241625 239864
rect 241286 239806 241625 239808
rect 240317 239730 240383 239733
rect 240136 239728 240383 239730
rect 239876 239668 239882 239704
rect 240136 239672 240322 239728
rect 240378 239672 240383 239728
rect 240136 239670 240383 239672
rect 240317 239667 240383 239670
rect 240542 239668 240548 239732
rect 240612 239730 240618 239732
rect 240777 239730 240843 239733
rect 240910 239730 240916 239732
rect 240612 239728 240916 239730
rect 240612 239672 240782 239728
rect 240838 239672 240916 239728
rect 240612 239670 240916 239672
rect 240612 239668 240618 239670
rect 240777 239667 240843 239670
rect 240910 239668 240916 239670
rect 240980 239668 240986 239732
rect 241094 239668 241100 239732
rect 241164 239730 241170 239732
rect 241286 239730 241346 239806
rect 241559 239803 241625 239806
rect 242014 239804 242020 239868
rect 242084 239842 242116 239868
rect 242172 239842 242177 239898
rect 245883 239898 245949 239903
rect 242084 239837 242177 239842
rect 242084 239806 242128 239837
rect 242084 239804 242090 239806
rect 242566 239804 242572 239868
rect 242636 239866 242642 239868
rect 244043 239866 244109 239869
rect 244779 239866 244845 239869
rect 245510 239866 245516 239868
rect 242636 239806 242864 239866
rect 242636 239804 242642 239806
rect 242804 239733 242864 239806
rect 244043 239864 244336 239866
rect 244043 239808 244048 239864
rect 244104 239808 244336 239864
rect 244043 239806 244336 239808
rect 244043 239803 244109 239806
rect 241164 239670 241346 239730
rect 241164 239668 241170 239670
rect 241646 239668 241652 239732
rect 241716 239730 241722 239732
rect 241973 239730 242039 239733
rect 241716 239728 242039 239730
rect 241716 239672 241978 239728
rect 242034 239672 242039 239728
rect 241716 239670 242039 239672
rect 241716 239668 241722 239670
rect 241973 239667 242039 239670
rect 242801 239728 242867 239733
rect 243997 239732 244063 239733
rect 242801 239672 242806 239728
rect 242862 239672 242867 239728
rect 242801 239667 242867 239672
rect 243486 239668 243492 239732
rect 243556 239730 243562 239732
rect 243997 239730 244044 239732
rect 243556 239728 244044 239730
rect 243556 239672 244002 239728
rect 243556 239670 244044 239672
rect 243556 239668 243562 239670
rect 243997 239668 244044 239670
rect 244108 239668 244114 239732
rect 244276 239730 244336 239806
rect 244779 239864 245516 239866
rect 244779 239808 244784 239864
rect 244840 239808 245516 239864
rect 244779 239806 245516 239808
rect 244779 239803 244845 239806
rect 245510 239804 245516 239806
rect 245580 239804 245586 239868
rect 245883 239842 245888 239898
rect 245944 239866 245949 239898
rect 246062 239866 246068 239868
rect 245944 239842 246068 239866
rect 245883 239837 246068 239842
rect 245886 239806 246068 239837
rect 246062 239804 246068 239806
rect 246132 239804 246138 239868
rect 246430 239804 246436 239868
rect 246500 239866 246506 239868
rect 246573 239866 246639 239869
rect 246500 239864 246639 239866
rect 246500 239808 246578 239864
rect 246634 239808 246639 239864
rect 246500 239806 246639 239808
rect 246500 239804 246506 239806
rect 246573 239803 246639 239806
rect 244276 239670 245762 239730
rect 243997 239667 244063 239668
rect 157149 239594 157215 239597
rect 210693 239594 210759 239597
rect 157149 239592 210759 239594
rect 157149 239536 157154 239592
rect 157210 239536 210698 239592
rect 210754 239536 210759 239592
rect 157149 239534 210759 239536
rect 157149 239531 157215 239534
rect 210693 239531 210759 239534
rect 212901 239594 212967 239597
rect 245702 239594 245762 239670
rect 245878 239668 245884 239732
rect 245948 239730 245954 239732
rect 246573 239730 246639 239733
rect 246798 239730 246804 239732
rect 245948 239728 246804 239730
rect 245948 239672 246578 239728
rect 246634 239672 246804 239728
rect 245948 239670 246804 239672
rect 245948 239668 245954 239670
rect 246573 239667 246639 239670
rect 246798 239668 246804 239670
rect 246868 239668 246874 239732
rect 246944 239730 247004 240078
rect 249014 240078 259010 240138
rect 261158 240272 282519 240274
rect 261158 240216 281538 240272
rect 281594 240216 282458 240272
rect 282514 240216 282519 240272
rect 261158 240214 282519 240216
rect 247723 239898 247789 239903
rect 247171 239866 247237 239869
rect 247350 239866 247356 239868
rect 247171 239864 247356 239866
rect 247171 239808 247176 239864
rect 247232 239808 247356 239864
rect 247171 239806 247356 239808
rect 247171 239803 247237 239806
rect 247350 239804 247356 239806
rect 247420 239804 247426 239868
rect 247534 239804 247540 239868
rect 247604 239866 247610 239868
rect 247723 239866 247728 239898
rect 247604 239842 247728 239866
rect 247784 239842 247789 239898
rect 249014 239869 249074 240078
rect 257102 240002 257108 240004
rect 257064 239940 257108 240002
rect 257172 239940 257178 240004
rect 258390 240002 258396 240004
rect 258168 239942 258396 240002
rect 247604 239837 247789 239842
rect 248551 239866 248617 239869
rect 248822 239866 248828 239868
rect 248551 239864 248828 239866
rect 247604 239806 247786 239837
rect 248551 239808 248556 239864
rect 248612 239808 248828 239864
rect 248551 239806 248828 239808
rect 247604 239804 247610 239806
rect 248551 239803 248617 239806
rect 248822 239804 248828 239806
rect 248892 239804 248898 239868
rect 248965 239864 249074 239869
rect 248965 239808 248970 239864
rect 249026 239808 249074 239864
rect 249747 239898 249813 239903
rect 249747 239842 249752 239898
rect 249808 239866 249813 239898
rect 251955 239898 252021 239903
rect 249926 239866 249932 239868
rect 249808 239842 249932 239866
rect 249747 239837 249932 239842
rect 248965 239806 249074 239808
rect 249750 239806 249932 239837
rect 248965 239803 249031 239806
rect 249926 239804 249932 239806
rect 249996 239804 250002 239868
rect 250110 239804 250116 239868
rect 250180 239866 250186 239868
rect 250529 239866 250595 239869
rect 251955 239868 251960 239898
rect 252016 239868 252021 239898
rect 253059 239898 253125 239903
rect 250180 239864 250595 239866
rect 250180 239808 250534 239864
rect 250590 239808 250595 239864
rect 250180 239806 250595 239808
rect 250180 239804 250186 239806
rect 250529 239803 250595 239806
rect 251950 239804 251956 239868
rect 252020 239866 252026 239868
rect 252020 239806 252078 239866
rect 252020 239804 252026 239806
rect 252686 239804 252692 239868
rect 252756 239866 252762 239868
rect 253059 239866 253064 239898
rect 252756 239842 253064 239866
rect 253120 239842 253125 239898
rect 254347 239898 254413 239903
rect 252756 239837 253125 239842
rect 253243 239866 253309 239869
rect 253422 239866 253428 239868
rect 253243 239864 253428 239866
rect 252756 239806 253122 239837
rect 253243 239808 253248 239864
rect 253304 239808 253428 239864
rect 253243 239806 253428 239808
rect 252756 239804 252762 239806
rect 253243 239803 253309 239806
rect 253422 239804 253428 239806
rect 253492 239804 253498 239868
rect 253565 239866 253631 239869
rect 253703 239866 253769 239869
rect 253565 239864 253769 239866
rect 253565 239808 253570 239864
rect 253626 239808 253708 239864
rect 253764 239808 253769 239864
rect 254347 239842 254352 239898
rect 254408 239842 254413 239898
rect 254715 239898 254781 239903
rect 254715 239868 254720 239898
rect 254776 239868 254781 239898
rect 254899 239898 254965 239903
rect 254347 239837 254413 239842
rect 253565 239806 253769 239808
rect 253565 239803 253631 239806
rect 253703 239803 253769 239806
rect 254350 239733 254410 239837
rect 254710 239804 254716 239868
rect 254780 239866 254786 239868
rect 254780 239806 254838 239866
rect 254899 239842 254904 239898
rect 254960 239842 254965 239898
rect 254899 239837 254965 239842
rect 255543 239866 255609 239869
rect 255998 239866 256004 239868
rect 255543 239864 256004 239866
rect 254780 239804 254786 239806
rect 254902 239733 254962 239837
rect 255543 239808 255548 239864
rect 255604 239808 256004 239864
rect 255543 239806 256004 239808
rect 255543 239803 255609 239806
rect 255998 239804 256004 239806
rect 256068 239804 256074 239868
rect 257064 239866 257124 239940
rect 258168 239903 258228 239942
rect 258390 239940 258396 239942
rect 258460 239940 258466 240004
rect 259310 240002 259316 240004
rect 258582 239942 259316 240002
rect 258119 239898 258228 239903
rect 257199 239866 257265 239869
rect 257064 239864 257265 239866
rect 257064 239808 257204 239864
rect 257260 239808 257265 239864
rect 258119 239842 258124 239898
rect 258180 239842 258228 239898
rect 258582 239869 258642 239942
rect 259310 239940 259316 239942
rect 259380 239940 259386 240004
rect 261158 239903 261218 240214
rect 281533 240211 281599 240214
rect 282453 240211 282519 240214
rect 268653 240138 268719 240141
rect 263550 240136 268719 240138
rect 263550 240080 268658 240136
rect 268714 240080 268719 240136
rect 263550 240078 268719 240080
rect 261518 239940 261524 240004
rect 261588 240002 261594 240004
rect 262806 240002 262812 240004
rect 261588 239942 262812 240002
rect 261588 239940 261594 239942
rect 259499 239898 259565 239903
rect 258119 239840 258228 239842
rect 258303 239864 258369 239869
rect 258119 239837 258185 239840
rect 257064 239806 257265 239808
rect 257199 239803 257265 239806
rect 258303 239808 258308 239864
rect 258364 239808 258369 239864
rect 258303 239803 258369 239808
rect 258579 239864 258645 239869
rect 258763 239868 258829 239869
rect 258579 239808 258584 239864
rect 258640 239808 258645 239864
rect 258579 239803 258645 239808
rect 258758 239804 258764 239868
rect 258828 239866 258834 239868
rect 259126 239866 259132 239868
rect 258828 239806 259132 239866
rect 258828 239804 258834 239806
rect 259126 239804 259132 239806
rect 259196 239804 259202 239868
rect 259499 239842 259504 239898
rect 259560 239866 259565 239898
rect 261155 239898 261221 239903
rect 259678 239866 259684 239868
rect 259560 239842 259684 239866
rect 259499 239837 259684 239842
rect 259502 239806 259684 239837
rect 259678 239804 259684 239806
rect 259748 239804 259754 239868
rect 260230 239804 260236 239868
rect 260300 239866 260306 239868
rect 260787 239866 260853 239869
rect 260300 239864 260853 239866
rect 260300 239808 260792 239864
rect 260848 239808 260853 239864
rect 261155 239842 261160 239898
rect 261216 239842 261221 239898
rect 262032 239869 262092 239942
rect 262806 239940 262812 239942
rect 262876 239940 262882 240004
rect 263550 239903 263610 240078
rect 268653 240075 268719 240078
rect 270493 240138 270559 240141
rect 271086 240138 271092 240140
rect 270493 240136 271092 240138
rect 270493 240080 270498 240136
rect 270554 240080 271092 240136
rect 270493 240078 271092 240080
rect 270493 240075 270559 240078
rect 271086 240076 271092 240078
rect 271156 240076 271162 240140
rect 266302 239940 266308 240004
rect 266372 240002 266378 240004
rect 275553 240002 275619 240005
rect 266372 240000 275619 240002
rect 266372 239944 275558 240000
rect 275614 239944 275619 240000
rect 266372 239942 275619 239944
rect 266372 239940 266378 239942
rect 275553 239939 275619 239942
rect 263547 239898 263613 239903
rect 261155 239837 261221 239842
rect 261523 239864 261589 239869
rect 260300 239806 260853 239808
rect 260300 239804 260306 239806
rect 258763 239803 258829 239804
rect 260787 239803 260853 239806
rect 261523 239808 261528 239864
rect 261584 239808 261589 239864
rect 261523 239803 261589 239808
rect 262029 239864 262095 239869
rect 262627 239868 262693 239869
rect 262622 239866 262628 239868
rect 262029 239808 262034 239864
rect 262090 239808 262095 239864
rect 262029 239803 262095 239808
rect 262536 239806 262628 239866
rect 262622 239804 262628 239806
rect 262692 239804 262698 239868
rect 263087 239866 263153 239869
rect 263317 239866 263383 239869
rect 263087 239864 263383 239866
rect 263087 239808 263092 239864
rect 263148 239808 263322 239864
rect 263378 239808 263383 239864
rect 263547 239842 263552 239898
rect 263608 239842 263613 239898
rect 266031 239900 266097 239903
rect 266031 239898 266140 239900
rect 263547 239837 263613 239842
rect 264467 239866 264533 239869
rect 265387 239868 265453 239869
rect 265755 239868 265821 239869
rect 264646 239866 264652 239868
rect 264467 239864 264652 239866
rect 263087 239806 263383 239808
rect 262627 239803 262693 239804
rect 263087 239803 263153 239806
rect 263317 239803 263383 239806
rect 264467 239808 264472 239864
rect 264528 239808 264652 239864
rect 264467 239806 264652 239808
rect 264467 239803 264533 239806
rect 264646 239804 264652 239806
rect 264716 239804 264722 239868
rect 265382 239866 265388 239868
rect 265296 239806 265388 239866
rect 265382 239804 265388 239806
rect 265452 239804 265458 239868
rect 265750 239866 265756 239868
rect 265664 239806 265756 239866
rect 265750 239804 265756 239806
rect 265820 239804 265826 239868
rect 266031 239842 266036 239898
rect 266092 239868 266140 239898
rect 266092 239842 266124 239868
rect 266031 239837 266124 239842
rect 266080 239806 266124 239837
rect 266118 239804 266124 239806
rect 266188 239804 266194 239868
rect 266583 239866 266649 239869
rect 267641 239868 267707 239869
rect 267590 239866 267596 239868
rect 266583 239864 267596 239866
rect 267660 239864 267707 239868
rect 266583 239808 266588 239864
rect 266644 239808 267596 239864
rect 267702 239808 267707 239864
rect 266583 239806 267596 239808
rect 265387 239803 265453 239804
rect 265755 239803 265821 239804
rect 266583 239803 266649 239806
rect 267590 239804 267596 239806
rect 267660 239804 267707 239808
rect 267641 239803 267707 239804
rect 246944 239670 253950 239730
rect 254350 239728 254459 239733
rect 254350 239672 254398 239728
rect 254454 239672 254459 239728
rect 254350 239670 254459 239672
rect 246113 239594 246179 239597
rect 212901 239592 245210 239594
rect 212901 239536 212906 239592
rect 212962 239536 245210 239592
rect 212901 239534 245210 239536
rect 245702 239592 246179 239594
rect 245702 239536 246118 239592
rect 246174 239536 246179 239592
rect 245702 239534 246179 239536
rect 212901 239531 212967 239534
rect 153009 239458 153075 239461
rect 213453 239458 213519 239461
rect 223113 239460 223179 239461
rect 223062 239458 223068 239460
rect 153009 239456 213519 239458
rect 153009 239400 153014 239456
rect 153070 239400 213458 239456
rect 213514 239400 213519 239456
rect 153009 239398 213519 239400
rect 223022 239398 223068 239458
rect 223132 239456 223179 239460
rect 223174 239400 223179 239456
rect 153009 239395 153075 239398
rect 213453 239395 213519 239398
rect 223062 239396 223068 239398
rect 223132 239396 223179 239400
rect 223614 239396 223620 239460
rect 223684 239458 223690 239460
rect 224033 239458 224099 239461
rect 224493 239458 224559 239461
rect 223684 239456 224559 239458
rect 223684 239400 224038 239456
rect 224094 239400 224498 239456
rect 224554 239400 224559 239456
rect 223684 239398 224559 239400
rect 223684 239396 223690 239398
rect 223113 239395 223179 239396
rect 224033 239395 224099 239398
rect 224493 239395 224559 239398
rect 225229 239458 225295 239461
rect 226190 239458 226196 239460
rect 225229 239456 226196 239458
rect 225229 239400 225234 239456
rect 225290 239400 226196 239456
rect 225229 239398 226196 239400
rect 225229 239395 225295 239398
rect 226190 239396 226196 239398
rect 226260 239396 226266 239460
rect 226333 239458 226399 239461
rect 226793 239460 226859 239461
rect 226558 239458 226564 239460
rect 226333 239456 226564 239458
rect 226333 239400 226338 239456
rect 226394 239400 226564 239456
rect 226333 239398 226564 239400
rect 226333 239395 226399 239398
rect 226558 239396 226564 239398
rect 226628 239396 226634 239460
rect 226742 239396 226748 239460
rect 226812 239458 226859 239460
rect 226812 239456 226904 239458
rect 226854 239400 226904 239456
rect 226812 239398 226904 239400
rect 226812 239396 226859 239398
rect 227478 239396 227484 239460
rect 227548 239458 227554 239460
rect 227621 239458 227687 239461
rect 227548 239456 227687 239458
rect 227548 239400 227626 239456
rect 227682 239400 227687 239456
rect 227548 239398 227687 239400
rect 227548 239396 227554 239398
rect 226793 239395 226859 239396
rect 227621 239395 227687 239398
rect 228214 239396 228220 239460
rect 228284 239458 228290 239460
rect 228725 239458 228791 239461
rect 228284 239456 228791 239458
rect 228284 239400 228730 239456
rect 228786 239400 228791 239456
rect 228284 239398 228791 239400
rect 228284 239396 228290 239398
rect 228725 239395 228791 239398
rect 229645 239460 229711 239461
rect 229645 239456 229692 239460
rect 229756 239458 229762 239460
rect 231209 239458 231275 239461
rect 231945 239460 232011 239461
rect 231526 239458 231532 239460
rect 229645 239400 229650 239456
rect 229645 239396 229692 239400
rect 229756 239398 229802 239458
rect 231209 239456 231532 239458
rect 231209 239400 231214 239456
rect 231270 239400 231532 239456
rect 231209 239398 231532 239400
rect 229756 239396 229762 239398
rect 229645 239395 229711 239396
rect 231209 239395 231275 239398
rect 231526 239396 231532 239398
rect 231596 239396 231602 239460
rect 231894 239458 231900 239460
rect 231854 239398 231900 239458
rect 231964 239456 232011 239460
rect 232006 239400 232011 239456
rect 231894 239396 231900 239398
rect 231964 239396 232011 239400
rect 232078 239396 232084 239460
rect 232148 239458 232154 239460
rect 232630 239458 232636 239460
rect 232148 239398 232636 239458
rect 232148 239396 232154 239398
rect 232630 239396 232636 239398
rect 232700 239396 232706 239460
rect 232998 239396 233004 239460
rect 233068 239458 233074 239460
rect 233141 239458 233207 239461
rect 233068 239456 233207 239458
rect 233068 239400 233146 239456
rect 233202 239400 233207 239456
rect 233068 239398 233207 239400
rect 233068 239396 233074 239398
rect 231945 239395 232011 239396
rect 233141 239395 233207 239398
rect 233918 239396 233924 239460
rect 233988 239458 233994 239460
rect 234613 239458 234679 239461
rect 233988 239456 234679 239458
rect 233988 239400 234618 239456
rect 234674 239400 234679 239456
rect 233988 239398 234679 239400
rect 233988 239396 233994 239398
rect 234613 239395 234679 239398
rect 235257 239458 235323 239461
rect 237097 239460 237163 239461
rect 235390 239458 235396 239460
rect 235257 239456 235396 239458
rect 235257 239400 235262 239456
rect 235318 239400 235396 239456
rect 235257 239398 235396 239400
rect 235257 239395 235323 239398
rect 235390 239396 235396 239398
rect 235460 239396 235466 239460
rect 237046 239458 237052 239460
rect 237006 239398 237052 239458
rect 237116 239456 237163 239460
rect 237158 239400 237163 239456
rect 237046 239396 237052 239398
rect 237116 239396 237163 239400
rect 237097 239395 237163 239396
rect 237465 239458 237531 239461
rect 238150 239458 238156 239460
rect 237465 239456 238156 239458
rect 237465 239400 237470 239456
rect 237526 239400 238156 239456
rect 237465 239398 238156 239400
rect 237465 239395 237531 239398
rect 238150 239396 238156 239398
rect 238220 239396 238226 239460
rect 238845 239458 238911 239461
rect 239070 239458 239076 239460
rect 238845 239456 239076 239458
rect 238845 239400 238850 239456
rect 238906 239400 239076 239456
rect 238845 239398 239076 239400
rect 238845 239395 238911 239398
rect 239070 239396 239076 239398
rect 239140 239396 239146 239460
rect 239990 239396 239996 239460
rect 240060 239458 240066 239460
rect 240133 239458 240199 239461
rect 241329 239460 241395 239461
rect 241278 239458 241284 239460
rect 240060 239456 240199 239458
rect 240060 239400 240138 239456
rect 240194 239400 240199 239456
rect 240060 239398 240199 239400
rect 241238 239398 241284 239458
rect 241348 239456 241395 239460
rect 241390 239400 241395 239456
rect 240060 239396 240066 239398
rect 240133 239395 240199 239398
rect 241278 239396 241284 239398
rect 241348 239396 241395 239400
rect 241329 239395 241395 239396
rect 241973 239458 242039 239461
rect 242750 239458 242756 239460
rect 241973 239456 242756 239458
rect 241973 239400 241978 239456
rect 242034 239400 242756 239456
rect 241973 239398 242756 239400
rect 241973 239395 242039 239398
rect 242750 239396 242756 239398
rect 242820 239396 242826 239460
rect 244365 239458 244431 239461
rect 244774 239458 244780 239460
rect 244365 239456 244780 239458
rect 244365 239400 244370 239456
rect 244426 239400 244780 239456
rect 244365 239398 244780 239400
rect 244365 239395 244431 239398
rect 244774 239396 244780 239398
rect 244844 239396 244850 239460
rect 245150 239458 245210 239534
rect 246113 239531 246179 239534
rect 246246 239532 246252 239596
rect 246316 239594 246322 239596
rect 247033 239594 247099 239597
rect 246316 239592 247099 239594
rect 246316 239536 247038 239592
rect 247094 239536 247099 239592
rect 246316 239534 247099 239536
rect 246316 239532 246322 239534
rect 247033 239531 247099 239534
rect 247166 239532 247172 239596
rect 247236 239594 247242 239596
rect 247309 239594 247375 239597
rect 247236 239592 247375 239594
rect 247236 239536 247314 239592
rect 247370 239536 247375 239592
rect 247236 239534 247375 239536
rect 247236 239532 247242 239534
rect 247309 239531 247375 239534
rect 247902 239532 247908 239596
rect 247972 239594 247978 239596
rect 248045 239594 248111 239597
rect 247972 239592 248111 239594
rect 247972 239536 248050 239592
rect 248106 239536 248111 239592
rect 247972 239534 248111 239536
rect 247972 239532 247978 239534
rect 248045 239531 248111 239534
rect 248597 239594 248663 239597
rect 248822 239594 248828 239596
rect 248597 239592 248828 239594
rect 248597 239536 248602 239592
rect 248658 239536 248828 239592
rect 248597 239534 248828 239536
rect 248597 239531 248663 239534
rect 248822 239532 248828 239534
rect 248892 239532 248898 239596
rect 249558 239532 249564 239596
rect 249628 239594 249634 239596
rect 249701 239594 249767 239597
rect 250621 239596 250687 239597
rect 250621 239594 250668 239596
rect 249628 239592 249767 239594
rect 249628 239536 249706 239592
rect 249762 239536 249767 239592
rect 249628 239534 249767 239536
rect 250576 239592 250668 239594
rect 250576 239536 250626 239592
rect 250576 239534 250668 239536
rect 249628 239532 249634 239534
rect 249701 239531 249767 239534
rect 250621 239532 250668 239534
rect 250732 239532 250738 239596
rect 250897 239594 250963 239597
rect 251030 239594 251036 239596
rect 250897 239592 251036 239594
rect 250897 239536 250902 239592
rect 250958 239536 251036 239592
rect 250897 239534 251036 239536
rect 250621 239531 250687 239532
rect 250897 239531 250963 239534
rect 251030 239532 251036 239534
rect 251100 239532 251106 239596
rect 251766 239532 251772 239596
rect 251836 239594 251842 239596
rect 252829 239594 252895 239597
rect 251836 239592 252895 239594
rect 251836 239536 252834 239592
rect 252890 239536 252895 239592
rect 251836 239534 252895 239536
rect 253890 239594 253950 239670
rect 254393 239667 254459 239670
rect 254853 239728 254962 239733
rect 254853 239672 254858 239728
rect 254914 239672 254962 239728
rect 254853 239670 254962 239672
rect 255129 239730 255195 239733
rect 255814 239730 255820 239732
rect 255129 239728 255820 239730
rect 255129 239672 255134 239728
rect 255190 239672 255820 239728
rect 255129 239670 255820 239672
rect 254853 239667 254919 239670
rect 255129 239667 255195 239670
rect 255814 239668 255820 239670
rect 255884 239668 255890 239732
rect 255957 239730 256023 239733
rect 256550 239730 256556 239732
rect 255957 239728 256556 239730
rect 255957 239672 255962 239728
rect 256018 239672 256556 239728
rect 255957 239670 256556 239672
rect 255957 239667 256023 239670
rect 256550 239668 256556 239670
rect 256620 239668 256626 239732
rect 256918 239668 256924 239732
rect 256988 239730 256994 239732
rect 257061 239730 257127 239733
rect 256988 239728 257127 239730
rect 256988 239672 257066 239728
rect 257122 239672 257127 239728
rect 256988 239670 257127 239672
rect 256988 239668 256994 239670
rect 257061 239667 257127 239670
rect 257245 239730 257311 239733
rect 257797 239730 257863 239733
rect 257245 239728 257863 239730
rect 257245 239672 257250 239728
rect 257306 239672 257802 239728
rect 257858 239672 257863 239728
rect 257245 239670 257863 239672
rect 258306 239730 258366 239803
rect 259494 239730 259500 239732
rect 258306 239670 259500 239730
rect 257245 239667 257311 239670
rect 257797 239667 257863 239670
rect 259494 239668 259500 239670
rect 259564 239668 259570 239732
rect 259637 239730 259703 239733
rect 260833 239732 260899 239733
rect 259862 239730 259868 239732
rect 259637 239728 259868 239730
rect 259637 239672 259642 239728
rect 259698 239672 259868 239728
rect 259637 239670 259868 239672
rect 259637 239667 259703 239670
rect 259862 239668 259868 239670
rect 259932 239668 259938 239732
rect 260782 239730 260788 239732
rect 260742 239670 260788 239730
rect 260852 239728 260899 239732
rect 260894 239672 260899 239728
rect 260782 239668 260788 239670
rect 260852 239668 260899 239672
rect 260966 239668 260972 239732
rect 261036 239730 261042 239732
rect 261526 239730 261586 239803
rect 262213 239732 262279 239733
rect 262213 239730 262260 239732
rect 261036 239670 261586 239730
rect 262168 239728 262260 239730
rect 262168 239672 262218 239728
rect 262168 239670 262260 239672
rect 261036 239668 261042 239670
rect 262213 239668 262260 239670
rect 262324 239668 262330 239732
rect 262673 239730 262739 239733
rect 266302 239730 266308 239732
rect 262673 239728 266308 239730
rect 262673 239672 262678 239728
rect 262734 239672 266308 239728
rect 262673 239670 266308 239672
rect 260833 239667 260899 239668
rect 262213 239667 262279 239668
rect 262673 239667 262739 239670
rect 266302 239668 266308 239670
rect 266372 239668 266378 239732
rect 266629 239730 266695 239733
rect 271822 239730 271828 239732
rect 266629 239728 271828 239730
rect 266629 239672 266634 239728
rect 266690 239672 271828 239728
rect 266629 239670 271828 239672
rect 266629 239667 266695 239670
rect 271822 239668 271828 239670
rect 271892 239668 271898 239732
rect 269573 239594 269639 239597
rect 253890 239592 269639 239594
rect 253890 239536 269578 239592
rect 269634 239536 269639 239592
rect 253890 239534 269639 239536
rect 251836 239532 251842 239534
rect 252829 239531 252895 239534
rect 269573 239531 269639 239534
rect 245150 239398 248568 239458
rect 248508 239325 248568 239398
rect 249374 239396 249380 239460
rect 249444 239458 249450 239460
rect 250110 239458 250116 239460
rect 249444 239398 250116 239458
rect 249444 239396 249450 239398
rect 250110 239396 250116 239398
rect 250180 239396 250186 239460
rect 250253 239458 250319 239461
rect 250846 239458 250852 239460
rect 250253 239456 250852 239458
rect 250253 239400 250258 239456
rect 250314 239400 250852 239456
rect 250253 239398 250852 239400
rect 250253 239395 250319 239398
rect 250846 239396 250852 239398
rect 250916 239396 250922 239460
rect 255405 239458 255471 239461
rect 255957 239458 256023 239461
rect 256182 239458 256188 239460
rect 255405 239456 256188 239458
rect 255405 239400 255410 239456
rect 255466 239400 255962 239456
rect 256018 239400 256188 239456
rect 255405 239398 256188 239400
rect 255405 239395 255471 239398
rect 255957 239395 256023 239398
rect 256182 239396 256188 239398
rect 256252 239396 256258 239460
rect 256877 239458 256943 239461
rect 257286 239458 257292 239460
rect 256877 239456 257292 239458
rect 256877 239400 256882 239456
rect 256938 239400 257292 239456
rect 256877 239398 257292 239400
rect 256877 239395 256943 239398
rect 257286 239396 257292 239398
rect 257356 239396 257362 239460
rect 258533 239458 258599 239461
rect 258717 239458 258783 239461
rect 258533 239456 258783 239458
rect 258533 239400 258538 239456
rect 258594 239400 258722 239456
rect 258778 239400 258783 239456
rect 258533 239398 258783 239400
rect 258533 239395 258599 239398
rect 258717 239395 258783 239398
rect 259913 239458 259979 239461
rect 260598 239458 260604 239460
rect 259913 239456 260604 239458
rect 259913 239400 259918 239456
rect 259974 239400 260604 239456
rect 259913 239398 260604 239400
rect 259913 239395 259979 239398
rect 260598 239396 260604 239398
rect 260668 239396 260674 239460
rect 261334 239396 261340 239460
rect 261404 239458 261410 239460
rect 262213 239458 262279 239461
rect 261404 239456 262279 239458
rect 261404 239400 262218 239456
rect 262274 239400 262279 239456
rect 261404 239398 262279 239400
rect 261404 239396 261410 239398
rect 262213 239395 262279 239398
rect 262765 239458 262831 239461
rect 263174 239458 263180 239460
rect 262765 239456 263180 239458
rect 262765 239400 262770 239456
rect 262826 239400 263180 239456
rect 262765 239398 263180 239400
rect 262765 239395 262831 239398
rect 263174 239396 263180 239398
rect 263244 239396 263250 239460
rect 266629 239458 266695 239461
rect 263504 239456 266695 239458
rect 263504 239400 266634 239456
rect 266690 239400 266695 239456
rect 263504 239398 266695 239400
rect 210693 239322 210759 239325
rect 226425 239322 226491 239325
rect 227345 239324 227411 239325
rect 227294 239322 227300 239324
rect 210693 239320 226491 239322
rect 210693 239264 210698 239320
rect 210754 239264 226430 239320
rect 226486 239264 226491 239320
rect 210693 239262 226491 239264
rect 227254 239262 227300 239322
rect 227364 239320 227411 239324
rect 233325 239322 233391 239325
rect 227406 239264 227411 239320
rect 210693 239259 210759 239262
rect 226425 239259 226491 239262
rect 227294 239260 227300 239262
rect 227364 239260 227411 239264
rect 227345 239259 227411 239260
rect 227670 239320 233391 239322
rect 227670 239264 233330 239320
rect 233386 239264 233391 239320
rect 227670 239262 233391 239264
rect 217317 239186 217383 239189
rect 227670 239186 227730 239262
rect 233325 239259 233391 239262
rect 233550 239260 233556 239324
rect 233620 239322 233626 239324
rect 233969 239322 234035 239325
rect 233620 239320 234035 239322
rect 233620 239264 233974 239320
rect 234030 239264 234035 239320
rect 233620 239262 234035 239264
rect 233620 239260 233626 239262
rect 233969 239259 234035 239262
rect 234245 239322 234311 239325
rect 234654 239322 234660 239324
rect 234245 239320 234660 239322
rect 234245 239264 234250 239320
rect 234306 239264 234660 239320
rect 234245 239262 234660 239264
rect 234245 239259 234311 239262
rect 234654 239260 234660 239262
rect 234724 239260 234730 239324
rect 237230 239260 237236 239324
rect 237300 239322 237306 239324
rect 247166 239322 247172 239324
rect 237300 239262 247172 239322
rect 237300 239260 237306 239262
rect 247166 239260 247172 239262
rect 247236 239260 247242 239324
rect 248505 239322 248571 239325
rect 249701 239322 249767 239325
rect 251357 239322 251423 239325
rect 248505 239320 249442 239322
rect 248505 239264 248510 239320
rect 248566 239264 249442 239320
rect 248505 239262 249442 239264
rect 248505 239259 248571 239262
rect 217317 239184 227730 239186
rect 217317 239128 217322 239184
rect 217378 239128 227730 239184
rect 217317 239126 227730 239128
rect 229277 239186 229343 239189
rect 230105 239188 230171 239189
rect 229870 239186 229876 239188
rect 229277 239184 229876 239186
rect 229277 239128 229282 239184
rect 229338 239128 229876 239184
rect 229277 239126 229876 239128
rect 217317 239123 217383 239126
rect 229277 239123 229343 239126
rect 229870 239124 229876 239126
rect 229940 239124 229946 239188
rect 230054 239124 230060 239188
rect 230124 239186 230171 239188
rect 232037 239186 232103 239189
rect 232446 239186 232452 239188
rect 230124 239184 230216 239186
rect 230166 239128 230216 239184
rect 230124 239126 230216 239128
rect 232037 239184 232452 239186
rect 232037 239128 232042 239184
rect 232098 239128 232452 239184
rect 232037 239126 232452 239128
rect 230124 239124 230171 239126
rect 230105 239123 230171 239124
rect 232037 239123 232103 239126
rect 232446 239124 232452 239126
rect 232516 239124 232522 239188
rect 233182 239124 233188 239188
rect 233252 239186 233258 239188
rect 233252 239126 244290 239186
rect 233252 239124 233258 239126
rect 205081 239050 205147 239053
rect 224125 239050 224191 239053
rect 205081 239048 224191 239050
rect 205081 238992 205086 239048
rect 205142 238992 224130 239048
rect 224186 238992 224191 239048
rect 205081 238990 224191 238992
rect 205081 238987 205147 238990
rect 224125 238987 224191 238990
rect 225045 239050 225111 239053
rect 225454 239050 225460 239052
rect 225045 239048 225460 239050
rect 225045 238992 225050 239048
rect 225106 238992 225460 239048
rect 225045 238990 225460 238992
rect 225045 238987 225111 238990
rect 225454 238988 225460 238990
rect 225524 239050 225530 239052
rect 226374 239050 226380 239052
rect 225524 238990 226380 239050
rect 225524 238988 225530 238990
rect 226374 238988 226380 238990
rect 226444 238988 226450 239052
rect 226517 239050 226583 239053
rect 227110 239050 227116 239052
rect 226517 239048 227116 239050
rect 226517 238992 226522 239048
rect 226578 238992 227116 239048
rect 226517 238990 227116 238992
rect 226517 238987 226583 238990
rect 227110 238988 227116 238990
rect 227180 238988 227186 239052
rect 228030 238988 228036 239052
rect 228100 239050 228106 239052
rect 237230 239050 237236 239052
rect 228100 238990 237236 239050
rect 228100 238988 228106 238990
rect 237230 238988 237236 238990
rect 237300 238988 237306 239052
rect 239673 239050 239739 239053
rect 241513 239050 241579 239053
rect 239673 239048 241579 239050
rect 239673 238992 239678 239048
rect 239734 238992 241518 239048
rect 241574 238992 241579 239048
rect 239673 238990 241579 238992
rect 244230 239050 244290 239126
rect 244958 239124 244964 239188
rect 245028 239186 245034 239188
rect 245561 239186 245627 239189
rect 245028 239184 245627 239186
rect 245028 239128 245566 239184
rect 245622 239128 245627 239184
rect 245028 239126 245627 239128
rect 245028 239124 245034 239126
rect 245561 239123 245627 239126
rect 245929 239186 245995 239189
rect 246062 239186 246068 239188
rect 245929 239184 246068 239186
rect 245929 239128 245934 239184
rect 245990 239128 246068 239184
rect 245929 239126 246068 239128
rect 245929 239123 245995 239126
rect 246062 239124 246068 239126
rect 246132 239124 246138 239188
rect 246389 239186 246455 239189
rect 247401 239186 247467 239189
rect 246389 239184 247467 239186
rect 246389 239128 246394 239184
rect 246450 239128 247406 239184
rect 247462 239128 247467 239184
rect 246389 239126 247467 239128
rect 246389 239123 246455 239126
rect 247401 239123 247467 239126
rect 249149 239188 249215 239189
rect 249149 239184 249196 239188
rect 249260 239186 249266 239188
rect 249382 239186 249442 239262
rect 249701 239320 251423 239322
rect 249701 239264 249706 239320
rect 249762 239264 251362 239320
rect 251418 239264 251423 239320
rect 249701 239262 251423 239264
rect 249701 239259 249767 239262
rect 251357 239259 251423 239262
rect 252185 239322 252251 239325
rect 263504 239322 263564 239398
rect 266629 239395 266695 239398
rect 252185 239320 263564 239322
rect 252185 239264 252190 239320
rect 252246 239264 263564 239320
rect 252185 239262 263564 239264
rect 264237 239322 264303 239325
rect 265709 239322 265775 239325
rect 264237 239320 265775 239322
rect 264237 239264 264242 239320
rect 264298 239264 265714 239320
rect 265770 239264 265775 239320
rect 264237 239262 265775 239264
rect 252185 239259 252251 239262
rect 264237 239259 264303 239262
rect 265709 239259 265775 239262
rect 266077 239324 266143 239325
rect 266077 239320 266124 239324
rect 266188 239322 266194 239324
rect 267273 239322 267339 239325
rect 267406 239322 267412 239324
rect 266077 239264 266082 239320
rect 266077 239260 266124 239264
rect 266188 239262 266234 239322
rect 267273 239320 267412 239322
rect 267273 239264 267278 239320
rect 267334 239264 267412 239320
rect 267273 239262 267412 239264
rect 266188 239260 266194 239262
rect 266077 239259 266143 239260
rect 267273 239259 267339 239262
rect 267406 239260 267412 239262
rect 267476 239260 267482 239324
rect 271229 239322 271295 239325
rect 271229 239320 282930 239322
rect 271229 239264 271234 239320
rect 271290 239264 282930 239320
rect 271229 239262 282930 239264
rect 271229 239259 271295 239262
rect 262121 239186 262187 239189
rect 274909 239186 274975 239189
rect 249149 239128 249154 239184
rect 249149 239124 249196 239128
rect 249260 239126 249306 239186
rect 249382 239126 256710 239186
rect 249260 239124 249266 239126
rect 249149 239123 249215 239124
rect 255313 239050 255379 239053
rect 255865 239050 255931 239053
rect 256366 239050 256372 239052
rect 244230 238990 251190 239050
rect 239673 238987 239739 238990
rect 241513 238987 241579 238990
rect 209405 238914 209471 238917
rect 228449 238914 228515 238917
rect 209405 238912 228515 238914
rect 209405 238856 209410 238912
rect 209466 238856 228454 238912
rect 228510 238856 228515 238912
rect 209405 238854 228515 238856
rect 209405 238851 209471 238854
rect 228449 238851 228515 238854
rect 228725 238914 228791 238917
rect 247534 238914 247540 238916
rect 228725 238912 247540 238914
rect 228725 238856 228730 238912
rect 228786 238856 247540 238912
rect 228725 238854 247540 238856
rect 228725 238851 228791 238854
rect 247534 238852 247540 238854
rect 247604 238852 247610 238916
rect 248045 238914 248111 238917
rect 250529 238914 250595 238917
rect 248045 238912 250595 238914
rect 248045 238856 248050 238912
rect 248106 238856 250534 238912
rect 250590 238856 250595 238912
rect 248045 238854 250595 238856
rect 248045 238851 248111 238854
rect 250529 238851 250595 238854
rect 250897 238912 250963 238917
rect 250897 238856 250902 238912
rect 250958 238856 250963 238912
rect 250897 238851 250963 238856
rect 251130 238914 251190 238990
rect 255313 239048 256372 239050
rect 255313 238992 255318 239048
rect 255374 238992 255870 239048
rect 255926 238992 256372 239048
rect 255313 238990 256372 238992
rect 255313 238987 255379 238990
rect 255865 238987 255931 238990
rect 256366 238988 256372 238990
rect 256436 238988 256442 239052
rect 256650 239050 256710 239126
rect 262121 239184 274975 239186
rect 262121 239128 262126 239184
rect 262182 239128 274914 239184
rect 274970 239128 274975 239184
rect 262121 239126 274975 239128
rect 262121 239123 262187 239126
rect 274909 239123 274975 239126
rect 264421 239052 264487 239053
rect 264973 239052 265039 239053
rect 256650 238990 263610 239050
rect 260966 238914 260972 238916
rect 251130 238854 260972 238914
rect 260966 238852 260972 238854
rect 261036 238852 261042 238916
rect 262438 238852 262444 238916
rect 262508 238914 262514 238916
rect 262949 238914 263015 238917
rect 262508 238912 263015 238914
rect 262508 238856 262954 238912
rect 263010 238856 263015 238912
rect 262508 238854 263015 238856
rect 263550 238914 263610 238990
rect 264094 238988 264100 239052
rect 264164 239050 264170 239052
rect 264421 239050 264468 239052
rect 264164 239048 264468 239050
rect 264164 238992 264426 239048
rect 264164 238990 264468 238992
rect 264164 238988 264170 238990
rect 264421 238988 264468 238990
rect 264532 238988 264538 239052
rect 264973 239048 265020 239052
rect 265084 239050 265090 239052
rect 265433 239050 265499 239053
rect 270861 239050 270927 239053
rect 264973 238992 264978 239048
rect 264973 238988 265020 238992
rect 265084 238990 265130 239050
rect 265433 239048 270927 239050
rect 265433 238992 265438 239048
rect 265494 238992 270866 239048
rect 270922 238992 270927 239048
rect 265433 238990 270927 238992
rect 282870 239050 282930 239262
rect 288525 239050 288591 239053
rect 282870 239048 288591 239050
rect 282870 238992 288530 239048
rect 288586 238992 288591 239048
rect 282870 238990 288591 238992
rect 265084 238988 265090 238990
rect 264421 238987 264487 238988
rect 264973 238987 265039 238988
rect 265433 238987 265499 238990
rect 270861 238987 270927 238990
rect 288525 238987 288591 238990
rect 296069 238914 296135 238917
rect 263550 238912 296135 238914
rect 263550 238856 296074 238912
rect 296130 238856 296135 238912
rect 263550 238854 296135 238856
rect 262508 238852 262514 238854
rect 262949 238851 263015 238854
rect 296069 238851 296135 238854
rect 222694 238716 222700 238780
rect 222764 238778 222770 238780
rect 223389 238778 223455 238781
rect 223941 238780 224007 238781
rect 223941 238778 223988 238780
rect 222764 238776 223455 238778
rect 222764 238720 223394 238776
rect 223450 238720 223455 238776
rect 222764 238718 223455 238720
rect 223896 238776 223988 238778
rect 223896 238720 223946 238776
rect 223896 238718 223988 238720
rect 222764 238716 222770 238718
rect 223389 238715 223455 238718
rect 223941 238716 223988 238718
rect 224052 238716 224058 238780
rect 225781 238778 225847 238781
rect 237189 238780 237255 238781
rect 236494 238778 236500 238780
rect 225781 238776 236500 238778
rect 225781 238720 225786 238776
rect 225842 238720 236500 238776
rect 225781 238718 236500 238720
rect 223941 238715 224007 238716
rect 225781 238715 225847 238718
rect 236494 238716 236500 238718
rect 236564 238716 236570 238780
rect 237189 238776 237236 238780
rect 237300 238778 237306 238780
rect 238753 238778 238819 238781
rect 239254 238778 239260 238780
rect 237189 238720 237194 238776
rect 237189 238716 237236 238720
rect 237300 238718 237346 238778
rect 238753 238776 239260 238778
rect 238753 238720 238758 238776
rect 238814 238720 239260 238776
rect 238753 238718 239260 238720
rect 237300 238716 237306 238718
rect 237189 238715 237255 238716
rect 238753 238715 238819 238718
rect 239254 238716 239260 238718
rect 239324 238716 239330 238780
rect 240726 238716 240732 238780
rect 240796 238778 240802 238780
rect 244365 238778 244431 238781
rect 240796 238776 244431 238778
rect 240796 238720 244370 238776
rect 244426 238720 244431 238776
rect 240796 238718 244431 238720
rect 240796 238716 240802 238718
rect 244365 238715 244431 238718
rect 245377 238778 245443 238781
rect 247401 238778 247467 238781
rect 245377 238776 247467 238778
rect 245377 238720 245382 238776
rect 245438 238720 247406 238776
rect 247462 238720 247467 238776
rect 245377 238718 247467 238720
rect 245377 238715 245443 238718
rect 247401 238715 247467 238718
rect 250529 238778 250595 238781
rect 250900 238778 250960 238851
rect 250529 238776 250960 238778
rect 250529 238720 250534 238776
rect 250590 238720 250960 238776
rect 250529 238718 250960 238720
rect 258073 238778 258139 238781
rect 258809 238778 258875 238781
rect 258073 238776 258875 238778
rect 258073 238720 258078 238776
rect 258134 238720 258814 238776
rect 258870 238720 258875 238776
rect 258073 238718 258875 238720
rect 250529 238715 250595 238718
rect 258073 238715 258139 238718
rect 258809 238715 258875 238718
rect 262949 238778 263015 238781
rect 264973 238778 265039 238781
rect 262949 238776 265039 238778
rect 262949 238720 262954 238776
rect 263010 238720 264978 238776
rect 265034 238720 265039 238776
rect 262949 238718 265039 238720
rect 262949 238715 263015 238718
rect 264973 238715 265039 238718
rect 265198 238716 265204 238780
rect 265268 238778 265274 238780
rect 265525 238778 265591 238781
rect 265268 238776 265591 238778
rect 265268 238720 265530 238776
rect 265586 238720 265591 238776
rect 265268 238718 265591 238720
rect 265268 238716 265274 238718
rect 265525 238715 265591 238718
rect 265801 238778 265867 238781
rect 268377 238778 268443 238781
rect 332777 238778 332843 238781
rect 265801 238776 268443 238778
rect 265801 238720 265806 238776
rect 265862 238720 268382 238776
rect 268438 238720 268443 238776
rect 265801 238718 268443 238720
rect 265801 238715 265867 238718
rect 268377 238715 268443 238718
rect 275970 238776 332843 238778
rect 275970 238720 332782 238776
rect 332838 238720 332843 238776
rect 275970 238718 332843 238720
rect 210693 238642 210759 238645
rect 210969 238642 211035 238645
rect 226926 238642 226932 238644
rect 210693 238640 211035 238642
rect 210693 238584 210698 238640
rect 210754 238584 210974 238640
rect 211030 238584 211035 238640
rect 210693 238582 211035 238584
rect 210693 238579 210759 238582
rect 210969 238579 211035 238582
rect 215250 238582 226932 238642
rect 188286 238444 188292 238508
rect 188356 238506 188362 238508
rect 215250 238506 215310 238582
rect 226926 238580 226932 238582
rect 226996 238642 227002 238644
rect 227253 238642 227319 238645
rect 226996 238640 227319 238642
rect 226996 238584 227258 238640
rect 227314 238584 227319 238640
rect 226996 238582 227319 238584
rect 226996 238580 227002 238582
rect 227253 238579 227319 238582
rect 228081 238642 228147 238645
rect 228950 238642 228956 238644
rect 228081 238640 228956 238642
rect 228081 238584 228086 238640
rect 228142 238584 228956 238640
rect 228081 238582 228956 238584
rect 228081 238579 228147 238582
rect 228950 238580 228956 238582
rect 229020 238580 229026 238644
rect 229829 238642 229895 238645
rect 230657 238644 230723 238645
rect 230238 238642 230244 238644
rect 229829 238640 230244 238642
rect 229829 238584 229834 238640
rect 229890 238584 230244 238640
rect 229829 238582 230244 238584
rect 229829 238579 229895 238582
rect 230238 238580 230244 238582
rect 230308 238580 230314 238644
rect 230606 238642 230612 238644
rect 230566 238582 230612 238642
rect 230676 238640 230723 238644
rect 230718 238584 230723 238640
rect 230606 238580 230612 238582
rect 230676 238580 230723 238584
rect 230657 238579 230723 238580
rect 231301 238642 231367 238645
rect 234654 238642 234660 238644
rect 231301 238640 234660 238642
rect 231301 238584 231306 238640
rect 231362 238584 234660 238640
rect 231301 238582 234660 238584
rect 231301 238579 231367 238582
rect 234654 238580 234660 238582
rect 234724 238580 234730 238644
rect 244457 238642 244523 238645
rect 245142 238642 245148 238644
rect 244457 238640 245148 238642
rect 244457 238584 244462 238640
rect 244518 238584 245148 238640
rect 244457 238582 245148 238584
rect 244457 238579 244523 238582
rect 245142 238580 245148 238582
rect 245212 238580 245218 238644
rect 245377 238642 245443 238645
rect 245510 238642 245516 238644
rect 245377 238640 245516 238642
rect 245377 238584 245382 238640
rect 245438 238584 245516 238640
rect 245377 238582 245516 238584
rect 245377 238579 245443 238582
rect 245510 238580 245516 238582
rect 245580 238580 245586 238644
rect 247166 238580 247172 238644
rect 247236 238642 247242 238644
rect 247493 238642 247559 238645
rect 247236 238640 247559 238642
rect 247236 238584 247498 238640
rect 247554 238584 247559 238640
rect 247236 238582 247559 238584
rect 247236 238580 247242 238582
rect 247493 238579 247559 238582
rect 248270 238580 248276 238644
rect 248340 238642 248346 238644
rect 248413 238642 248479 238645
rect 248340 238640 248479 238642
rect 248340 238584 248418 238640
rect 248474 238584 248479 238640
rect 248340 238582 248479 238584
rect 248340 238580 248346 238582
rect 248413 238579 248479 238582
rect 250294 238580 250300 238644
rect 250364 238642 250370 238644
rect 252686 238642 252692 238644
rect 250364 238582 252692 238642
rect 250364 238580 250370 238582
rect 252686 238580 252692 238582
rect 252756 238580 252762 238644
rect 255630 238580 255636 238644
rect 255700 238642 255706 238644
rect 256877 238642 256943 238645
rect 255700 238640 256943 238642
rect 255700 238584 256882 238640
rect 256938 238584 256943 238640
rect 255700 238582 256943 238584
rect 255700 238580 255706 238582
rect 256877 238579 256943 238582
rect 258625 238642 258691 238645
rect 263961 238642 264027 238645
rect 258625 238640 264027 238642
rect 258625 238584 258630 238640
rect 258686 238584 263966 238640
rect 264022 238584 264027 238640
rect 258625 238582 264027 238584
rect 258625 238579 258691 238582
rect 263961 238579 264027 238582
rect 264513 238642 264579 238645
rect 264830 238642 264836 238644
rect 264513 238640 264836 238642
rect 264513 238584 264518 238640
rect 264574 238584 264836 238640
rect 264513 238582 264836 238584
rect 264513 238579 264579 238582
rect 264830 238580 264836 238582
rect 264900 238580 264906 238644
rect 265249 238642 265315 238645
rect 275970 238642 276030 238718
rect 332777 238715 332843 238718
rect 265249 238640 276030 238642
rect 265249 238584 265254 238640
rect 265310 238584 276030 238640
rect 265249 238582 276030 238584
rect 265249 238579 265315 238582
rect 188356 238446 215310 238506
rect 188356 238444 188362 238446
rect 223798 238444 223804 238508
rect 223868 238506 223874 238508
rect 224125 238506 224191 238509
rect 223868 238504 224191 238506
rect 223868 238448 224130 238504
rect 224186 238448 224191 238504
rect 223868 238446 224191 238448
rect 223868 238444 223874 238446
rect 224125 238443 224191 238446
rect 225229 238506 225295 238509
rect 225873 238506 225939 238509
rect 226006 238506 226012 238508
rect 225229 238504 226012 238506
rect 225229 238448 225234 238504
rect 225290 238448 225878 238504
rect 225934 238448 226012 238504
rect 225229 238446 226012 238448
rect 225229 238443 225295 238446
rect 225873 238443 225939 238446
rect 226006 238444 226012 238446
rect 226076 238444 226082 238508
rect 228173 238506 228239 238509
rect 229001 238506 229067 238509
rect 237097 238506 237163 238509
rect 263869 238506 263935 238509
rect 264278 238506 264284 238508
rect 228173 238504 232882 238506
rect 228173 238448 228178 238504
rect 228234 238448 229006 238504
rect 229062 238448 232882 238504
rect 228173 238446 232882 238448
rect 228173 238443 228239 238446
rect 229001 238443 229067 238446
rect 224401 238370 224467 238373
rect 227989 238370 228055 238373
rect 231025 238372 231091 238373
rect 230974 238370 230980 238372
rect 224401 238368 228055 238370
rect 224401 238312 224406 238368
rect 224462 238312 227994 238368
rect 228050 238312 228055 238368
rect 224401 238310 228055 238312
rect 230934 238310 230980 238370
rect 231044 238368 231091 238372
rect 232681 238370 232747 238373
rect 231086 238312 231091 238368
rect 224401 238307 224467 238310
rect 227989 238307 228055 238310
rect 230974 238308 230980 238310
rect 231044 238308 231091 238312
rect 231025 238307 231091 238308
rect 231166 238368 232747 238370
rect 231166 238312 232686 238368
rect 232742 238312 232747 238368
rect 231166 238310 232747 238312
rect 232822 238370 232882 238446
rect 237097 238504 263794 238506
rect 237097 238448 237102 238504
rect 237158 238448 263794 238504
rect 237097 238446 263794 238448
rect 237097 238443 237163 238446
rect 258625 238370 258691 238373
rect 232822 238368 258691 238370
rect 232822 238312 258630 238368
rect 258686 238312 258691 238368
rect 232822 238310 258691 238312
rect 263734 238370 263794 238446
rect 263869 238504 264284 238506
rect 263869 238448 263874 238504
rect 263930 238448 264284 238504
rect 263869 238446 264284 238448
rect 263869 238443 263935 238446
rect 264278 238444 264284 238446
rect 264348 238444 264354 238508
rect 266302 238444 266308 238508
rect 266372 238506 266378 238508
rect 266905 238506 266971 238509
rect 266372 238504 266971 238506
rect 266372 238448 266910 238504
rect 266966 238448 266971 238504
rect 266372 238446 266971 238448
rect 266372 238444 266378 238446
rect 266905 238443 266971 238446
rect 265893 238370 265959 238373
rect 270401 238370 270467 238373
rect 263734 238310 263978 238370
rect 186814 238172 186820 238236
rect 186884 238234 186890 238236
rect 210785 238234 210851 238237
rect 211061 238234 211127 238237
rect 186884 238232 211127 238234
rect 186884 238176 210790 238232
rect 210846 238176 211066 238232
rect 211122 238176 211127 238232
rect 186884 238174 211127 238176
rect 186884 238172 186890 238174
rect 210785 238171 210851 238174
rect 211061 238171 211127 238174
rect 221273 238234 221339 238237
rect 231166 238234 231226 238310
rect 232681 238307 232747 238310
rect 258625 238307 258691 238310
rect 258625 238234 258691 238237
rect 221273 238232 231226 238234
rect 221273 238176 221278 238232
rect 221334 238176 231226 238232
rect 221273 238174 231226 238176
rect 231534 238232 258691 238234
rect 231534 238176 258630 238232
rect 258686 238176 258691 238232
rect 231534 238174 258691 238176
rect 221273 238171 221339 238174
rect 175774 238036 175780 238100
rect 175844 238098 175850 238100
rect 208209 238098 208275 238101
rect 225873 238098 225939 238101
rect 175844 238096 225939 238098
rect 175844 238040 208214 238096
rect 208270 238040 225878 238096
rect 225934 238040 225939 238096
rect 175844 238038 225939 238040
rect 175844 238036 175850 238038
rect 208209 238035 208275 238038
rect 225873 238035 225939 238038
rect 226333 238098 226399 238101
rect 231534 238098 231594 238174
rect 258625 238171 258691 238174
rect 258901 238234 258967 238237
rect 259126 238234 259132 238236
rect 258901 238232 259132 238234
rect 258901 238176 258906 238232
rect 258962 238176 259132 238232
rect 258901 238174 259132 238176
rect 258901 238171 258967 238174
rect 259126 238172 259132 238174
rect 259196 238172 259202 238236
rect 263726 238234 263732 238236
rect 263550 238174 263732 238234
rect 226333 238096 231594 238098
rect 226333 238040 226338 238096
rect 226394 238040 231594 238096
rect 226333 238038 231594 238040
rect 231669 238098 231735 238101
rect 263550 238098 263610 238174
rect 263726 238172 263732 238174
rect 263796 238172 263802 238236
rect 263918 238234 263978 238310
rect 265893 238368 270467 238370
rect 265893 238312 265898 238368
rect 265954 238312 270406 238368
rect 270462 238312 270467 238368
rect 265893 238310 270467 238312
rect 265893 238307 265959 238310
rect 270401 238307 270467 238310
rect 270309 238234 270375 238237
rect 263918 238232 270375 238234
rect 263918 238176 270314 238232
rect 270370 238176 270375 238232
rect 263918 238174 270375 238176
rect 270309 238171 270375 238174
rect 270861 238234 270927 238237
rect 302141 238234 302207 238237
rect 270861 238232 302207 238234
rect 270861 238176 270866 238232
rect 270922 238176 302146 238232
rect 302202 238176 302207 238232
rect 270861 238174 302207 238176
rect 270861 238171 270927 238174
rect 302141 238171 302207 238174
rect 231669 238096 263610 238098
rect 231669 238040 231674 238096
rect 231730 238040 263610 238096
rect 231669 238038 263610 238040
rect 263961 238098 264027 238101
rect 268653 238098 268719 238101
rect 310646 238098 310652 238100
rect 263961 238096 266370 238098
rect 263961 238040 263966 238096
rect 264022 238040 266370 238096
rect 263961 238038 266370 238040
rect 226333 238035 226399 238038
rect 231669 238035 231735 238038
rect 263961 238035 264027 238038
rect 175958 237900 175964 237964
rect 176028 237962 176034 237964
rect 231577 237962 231643 237965
rect 241605 237964 241671 237965
rect 241605 237962 241652 237964
rect 176028 237960 231643 237962
rect 176028 237904 231582 237960
rect 231638 237904 231643 237960
rect 176028 237902 231643 237904
rect 241560 237960 241652 237962
rect 241560 237904 241610 237960
rect 241560 237902 241652 237904
rect 176028 237900 176034 237902
rect 231577 237899 231643 237902
rect 241605 237900 241652 237902
rect 241716 237900 241722 237964
rect 248505 237962 248571 237965
rect 249558 237962 249564 237964
rect 248505 237960 249564 237962
rect 248505 237904 248510 237960
rect 248566 237904 249564 237960
rect 248505 237902 249564 237904
rect 241605 237899 241671 237900
rect 248505 237899 248571 237902
rect 249558 237900 249564 237902
rect 249628 237900 249634 237964
rect 262622 237900 262628 237964
rect 262692 237962 262698 237964
rect 265801 237962 265867 237965
rect 262692 237960 265867 237962
rect 262692 237904 265806 237960
rect 265862 237904 265867 237960
rect 262692 237902 265867 237904
rect 266310 237962 266370 238038
rect 268653 238096 310652 238098
rect 268653 238040 268658 238096
rect 268714 238040 310652 238096
rect 268653 238038 310652 238040
rect 268653 238035 268719 238038
rect 310646 238036 310652 238038
rect 310716 238036 310722 238100
rect 270585 237962 270651 237965
rect 328729 237962 328795 237965
rect 266310 237960 270651 237962
rect 266310 237904 270590 237960
rect 270646 237904 270651 237960
rect 266310 237902 270651 237904
rect 262692 237900 262698 237902
rect 265801 237899 265867 237902
rect 270585 237899 270651 237902
rect 285630 237960 328795 237962
rect 285630 237904 328734 237960
rect 328790 237904 328795 237960
rect 285630 237902 328795 237904
rect 231158 237826 231164 237828
rect 223530 237766 231164 237826
rect 177246 237628 177252 237692
rect 177316 237690 177322 237692
rect 223530 237690 223590 237766
rect 231158 237764 231164 237766
rect 231228 237764 231234 237828
rect 237598 237764 237604 237828
rect 237668 237826 237674 237828
rect 238385 237826 238451 237829
rect 259729 237828 259795 237829
rect 237668 237824 238451 237826
rect 237668 237768 238390 237824
rect 238446 237768 238451 237824
rect 237668 237766 238451 237768
rect 237668 237764 237674 237766
rect 238385 237763 238451 237766
rect 242014 237764 242020 237828
rect 242084 237826 242090 237828
rect 246246 237826 246252 237828
rect 242084 237766 246252 237826
rect 242084 237764 242090 237766
rect 246246 237764 246252 237766
rect 246316 237764 246322 237828
rect 259678 237764 259684 237828
rect 259748 237826 259795 237828
rect 260281 237826 260347 237829
rect 260598 237826 260604 237828
rect 259748 237824 259840 237826
rect 259790 237768 259840 237824
rect 259748 237766 259840 237768
rect 260281 237824 260604 237826
rect 260281 237768 260286 237824
rect 260342 237768 260604 237824
rect 260281 237766 260604 237768
rect 259748 237764 259795 237766
rect 259729 237763 259795 237764
rect 260281 237763 260347 237766
rect 260598 237764 260604 237766
rect 260668 237764 260674 237828
rect 264881 237826 264947 237829
rect 267774 237826 267780 237828
rect 264881 237824 267780 237826
rect 264881 237768 264886 237824
rect 264942 237768 267780 237824
rect 264881 237766 267780 237768
rect 264881 237763 264947 237766
rect 267774 237764 267780 237766
rect 267844 237826 267850 237828
rect 285630 237826 285690 237902
rect 328729 237899 328795 237902
rect 267844 237766 285690 237826
rect 267844 237764 267850 237766
rect 177316 237630 223590 237690
rect 229093 237690 229159 237693
rect 236637 237690 236703 237693
rect 229093 237688 236703 237690
rect 229093 237632 229098 237688
rect 229154 237632 236642 237688
rect 236698 237632 236703 237688
rect 229093 237630 236703 237632
rect 177316 237628 177322 237630
rect 229093 237627 229159 237630
rect 236637 237627 236703 237630
rect 245101 237690 245167 237693
rect 247902 237690 247908 237692
rect 245101 237688 247908 237690
rect 245101 237632 245106 237688
rect 245162 237632 247908 237688
rect 245101 237630 247908 237632
rect 245101 237627 245167 237630
rect 247902 237628 247908 237630
rect 247972 237628 247978 237692
rect 251541 237690 251607 237693
rect 252318 237690 252324 237692
rect 251541 237688 252324 237690
rect 251541 237632 251546 237688
rect 251602 237632 252324 237688
rect 251541 237630 252324 237632
rect 251541 237627 251607 237630
rect 252318 237628 252324 237630
rect 252388 237628 252394 237692
rect 254485 237690 254551 237693
rect 255446 237690 255452 237692
rect 254485 237688 255452 237690
rect 254485 237632 254490 237688
rect 254546 237632 255452 237688
rect 254485 237630 255452 237632
rect 254485 237627 254551 237630
rect 255446 237628 255452 237630
rect 255516 237628 255522 237692
rect 258625 237690 258691 237693
rect 265934 237690 265940 237692
rect 258625 237688 265940 237690
rect 258625 237632 258630 237688
rect 258686 237632 265940 237688
rect 258625 237630 265940 237632
rect 258625 237627 258691 237630
rect 265934 237628 265940 237630
rect 266004 237628 266010 237692
rect 229553 237554 229619 237557
rect 213870 237552 229619 237554
rect 213870 237496 229558 237552
rect 229614 237496 229619 237552
rect 213870 237494 229619 237496
rect 211061 237418 211127 237421
rect 213870 237418 213930 237494
rect 229553 237491 229619 237494
rect 231209 237554 231275 237557
rect 268285 237554 268351 237557
rect 231209 237552 268351 237554
rect 231209 237496 231214 237552
rect 231270 237496 268290 237552
rect 268346 237496 268351 237552
rect 231209 237494 268351 237496
rect 231209 237491 231275 237494
rect 268285 237491 268351 237494
rect 211061 237416 213930 237418
rect 211061 237360 211066 237416
rect 211122 237360 213930 237416
rect 211061 237358 213930 237360
rect 230473 237418 230539 237421
rect 231342 237418 231348 237420
rect 230473 237416 231348 237418
rect 230473 237360 230478 237416
rect 230534 237360 231348 237416
rect 230473 237358 231348 237360
rect 211061 237355 211127 237358
rect 230473 237355 230539 237358
rect 231342 237356 231348 237358
rect 231412 237356 231418 237420
rect 249977 237418 250043 237421
rect 251030 237418 251036 237420
rect 249977 237416 251036 237418
rect 249977 237360 249982 237416
rect 250038 237360 251036 237416
rect 249977 237358 251036 237360
rect 249977 237355 250043 237358
rect 251030 237356 251036 237358
rect 251100 237356 251106 237420
rect 252686 237356 252692 237420
rect 252756 237418 252762 237420
rect 253289 237418 253355 237421
rect 252756 237416 253355 237418
rect 252756 237360 253294 237416
rect 253350 237360 253355 237416
rect 252756 237358 253355 237360
rect 252756 237356 252762 237358
rect 253289 237355 253355 237358
rect 258625 237418 258691 237421
rect 260373 237420 260439 237421
rect 258758 237418 258764 237420
rect 258625 237416 258764 237418
rect 258625 237360 258630 237416
rect 258686 237360 258764 237416
rect 258625 237358 258764 237360
rect 258625 237355 258691 237358
rect 258758 237356 258764 237358
rect 258828 237356 258834 237420
rect 260373 237416 260420 237420
rect 260484 237418 260490 237420
rect 260741 237418 260807 237421
rect 268929 237418 268995 237421
rect 260373 237360 260378 237416
rect 260373 237356 260420 237360
rect 260484 237358 260530 237418
rect 260741 237416 268995 237418
rect 260741 237360 260746 237416
rect 260802 237360 268934 237416
rect 268990 237360 268995 237416
rect 260741 237358 268995 237360
rect 260484 237356 260490 237358
rect 260373 237355 260439 237356
rect 260741 237355 260807 237358
rect 268929 237355 268995 237358
rect 269389 237418 269455 237421
rect 269573 237418 269639 237421
rect 271689 237418 271755 237421
rect 269389 237416 271755 237418
rect 269389 237360 269394 237416
rect 269450 237360 269578 237416
rect 269634 237360 271694 237416
rect 271750 237360 271755 237416
rect 269389 237358 271755 237360
rect 269389 237355 269455 237358
rect 269573 237355 269639 237358
rect 271689 237355 271755 237358
rect 211981 237282 212047 237285
rect 228449 237282 228515 237285
rect 211981 237280 228515 237282
rect 211981 237224 211986 237280
rect 212042 237224 228454 237280
rect 228510 237224 228515 237280
rect 211981 237222 228515 237224
rect 211981 237219 212047 237222
rect 228449 237219 228515 237222
rect 253289 237282 253355 237285
rect 254393 237282 254459 237285
rect 253289 237280 254459 237282
rect 253289 237224 253294 237280
rect 253350 237224 254398 237280
rect 254454 237224 254459 237280
rect 253289 237222 254459 237224
rect 253289 237219 253355 237222
rect 254393 237219 254459 237222
rect 265709 237282 265775 237285
rect 268326 237282 268332 237284
rect 265709 237280 268332 237282
rect 265709 237224 265714 237280
rect 265770 237224 268332 237280
rect 265709 237222 268332 237224
rect 265709 237219 265775 237222
rect 268326 237220 268332 237222
rect 268396 237282 268402 237284
rect 333145 237282 333211 237285
rect 268396 237280 333211 237282
rect 268396 237224 333150 237280
rect 333206 237224 333211 237280
rect 268396 237222 333211 237224
rect 268396 237220 268402 237222
rect 333145 237219 333211 237222
rect 220721 237146 220787 237149
rect 234981 237146 235047 237149
rect 220721 237144 235047 237146
rect 220721 237088 220726 237144
rect 220782 237088 234986 237144
rect 235042 237088 235047 237144
rect 220721 237086 235047 237088
rect 220721 237083 220787 237086
rect 234981 237083 235047 237086
rect 263685 237146 263751 237149
rect 298185 237146 298251 237149
rect 298829 237146 298895 237149
rect 263685 237144 298895 237146
rect 263685 237088 263690 237144
rect 263746 237088 298190 237144
rect 298246 237088 298834 237144
rect 298890 237088 298895 237144
rect 263685 237086 298895 237088
rect 263685 237083 263751 237086
rect 298185 237083 298251 237086
rect 298829 237083 298895 237086
rect 213821 237010 213887 237013
rect 236729 237010 236795 237013
rect 213821 237008 236795 237010
rect 213821 236952 213826 237008
rect 213882 236952 236734 237008
rect 236790 236952 236795 237008
rect 213821 236950 236795 236952
rect 213821 236947 213887 236950
rect 236729 236947 236795 236950
rect 244406 236948 244412 237012
rect 244476 237010 244482 237012
rect 245193 237010 245259 237013
rect 244476 237008 245259 237010
rect 244476 236952 245198 237008
rect 245254 236952 245259 237008
rect 244476 236950 245259 236952
rect 244476 236948 244482 236950
rect 245193 236947 245259 236950
rect 252134 236948 252140 237012
rect 252204 237010 252210 237012
rect 256325 237010 256391 237013
rect 252204 237008 256391 237010
rect 252204 236952 256330 237008
rect 256386 236952 256391 237008
rect 252204 236950 256391 236952
rect 252204 236948 252210 236950
rect 256325 236947 256391 236950
rect 262489 237010 262555 237013
rect 294045 237010 294111 237013
rect 262489 237008 294111 237010
rect 262489 236952 262494 237008
rect 262550 236952 294050 237008
rect 294106 236952 294111 237008
rect 262489 236950 294111 236952
rect 262489 236947 262555 236950
rect 294045 236947 294111 236950
rect 213085 236874 213151 236877
rect 218789 236874 218855 236877
rect 239949 236874 240015 236877
rect 247401 236876 247467 236877
rect 213085 236872 240015 236874
rect 213085 236816 213090 236872
rect 213146 236816 218794 236872
rect 218850 236816 239954 236872
rect 240010 236816 240015 236872
rect 213085 236814 240015 236816
rect 213085 236811 213151 236814
rect 218789 236811 218855 236814
rect 239949 236811 240015 236814
rect 247350 236812 247356 236876
rect 247420 236874 247467 236876
rect 255773 236874 255839 236877
rect 258390 236874 258396 236876
rect 247420 236872 247512 236874
rect 247462 236816 247512 236872
rect 247420 236814 247512 236816
rect 255773 236872 258396 236874
rect 255773 236816 255778 236872
rect 255834 236816 258396 236872
rect 255773 236814 258396 236816
rect 247420 236812 247467 236814
rect 247401 236811 247467 236812
rect 255773 236811 255839 236814
rect 258390 236812 258396 236814
rect 258460 236812 258466 236876
rect 261017 236874 261083 236877
rect 262070 236874 262076 236876
rect 261017 236872 262076 236874
rect 261017 236816 261022 236872
rect 261078 236816 262076 236872
rect 261017 236814 262076 236816
rect 261017 236811 261083 236814
rect 262070 236812 262076 236814
rect 262140 236812 262146 236876
rect 165838 236676 165844 236740
rect 165908 236738 165914 236740
rect 206645 236738 206711 236741
rect 165908 236736 206711 236738
rect 165908 236680 206650 236736
rect 206706 236680 206711 236736
rect 165908 236678 206711 236680
rect 165908 236676 165914 236678
rect 206645 236675 206711 236678
rect 216581 236738 216647 236741
rect 237189 236738 237255 236741
rect 216581 236736 237255 236738
rect 216581 236680 216586 236736
rect 216642 236680 237194 236736
rect 237250 236680 237255 236736
rect 216581 236678 237255 236680
rect 216581 236675 216647 236678
rect 237189 236675 237255 236678
rect 238150 236676 238156 236740
rect 238220 236738 238226 236740
rect 262622 236738 262628 236740
rect 238220 236678 262628 236738
rect 238220 236676 238226 236678
rect 262622 236676 262628 236678
rect 262692 236676 262698 236740
rect 270350 236676 270356 236740
rect 270420 236738 270426 236740
rect 270769 236738 270835 236741
rect 270420 236736 270835 236738
rect 270420 236680 270774 236736
rect 270830 236680 270835 236736
rect 270420 236678 270835 236680
rect 270420 236676 270426 236678
rect 270769 236675 270835 236678
rect 272149 236738 272215 236741
rect 272977 236738 273043 236741
rect 272149 236736 273043 236738
rect 272149 236680 272154 236736
rect 272210 236680 272982 236736
rect 273038 236680 273043 236736
rect 272149 236678 273043 236680
rect 272149 236675 272215 236678
rect 272977 236675 273043 236678
rect 173750 236540 173756 236604
rect 173820 236602 173826 236604
rect 233509 236602 233575 236605
rect 173820 236600 233575 236602
rect 173820 236544 233514 236600
rect 233570 236544 233575 236600
rect 173820 236542 233575 236544
rect 173820 236540 173826 236542
rect 233509 236539 233575 236542
rect 236494 236540 236500 236604
rect 236564 236602 236570 236604
rect 251766 236602 251772 236604
rect 236564 236542 251772 236602
rect 236564 236540 236570 236542
rect 251766 236540 251772 236542
rect 251836 236540 251842 236604
rect 255129 236602 255195 236605
rect 255262 236602 255268 236604
rect 255129 236600 255268 236602
rect 255129 236544 255134 236600
rect 255190 236544 255268 236600
rect 255129 236542 255268 236544
rect 255129 236539 255195 236542
rect 255262 236540 255268 236542
rect 255332 236540 255338 236604
rect 261937 236602 262003 236605
rect 288341 236602 288407 236605
rect 261937 236600 288407 236602
rect 261937 236544 261942 236600
rect 261998 236544 288346 236600
rect 288402 236544 288407 236600
rect 261937 236542 288407 236544
rect 261937 236539 262003 236542
rect 288341 236539 288407 236542
rect 222009 236466 222075 236469
rect 237741 236466 237807 236469
rect 222009 236464 237807 236466
rect 222009 236408 222014 236464
rect 222070 236408 237746 236464
rect 237802 236408 237807 236464
rect 222009 236406 237807 236408
rect 222009 236403 222075 236406
rect 237741 236403 237807 236406
rect 253473 236466 253539 236469
rect 272149 236466 272215 236469
rect 253473 236464 272215 236466
rect 253473 236408 253478 236464
rect 253534 236408 272154 236464
rect 272210 236408 272215 236464
rect 253473 236406 272215 236408
rect 253473 236403 253539 236406
rect 272149 236403 272215 236406
rect 227345 236330 227411 236333
rect 227478 236330 227484 236332
rect 227345 236328 227484 236330
rect 227345 236272 227350 236328
rect 227406 236272 227484 236328
rect 227345 236270 227484 236272
rect 227345 236267 227411 236270
rect 227478 236268 227484 236270
rect 227548 236268 227554 236332
rect 234838 236268 234844 236332
rect 234908 236330 234914 236332
rect 235441 236330 235507 236333
rect 234908 236328 235507 236330
rect 234908 236272 235446 236328
rect 235502 236272 235507 236328
rect 234908 236270 235507 236272
rect 234908 236268 234914 236270
rect 235441 236267 235507 236270
rect 255998 236268 256004 236332
rect 256068 236330 256074 236332
rect 256509 236330 256575 236333
rect 256068 236328 256575 236330
rect 256068 236272 256514 236328
rect 256570 236272 256575 236328
rect 256068 236270 256575 236272
rect 256068 236268 256074 236270
rect 256509 236267 256575 236270
rect 259453 236330 259519 236333
rect 272333 236330 272399 236333
rect 259453 236328 272399 236330
rect 259453 236272 259458 236328
rect 259514 236272 272338 236328
rect 272394 236272 272399 236328
rect 259453 236270 272399 236272
rect 259453 236267 259519 236270
rect 272333 236267 272399 236270
rect 213545 236058 213611 236061
rect 215385 236058 215451 236061
rect 216581 236058 216647 236061
rect 213545 236056 216647 236058
rect 213545 236000 213550 236056
rect 213606 236000 215390 236056
rect 215446 236000 216586 236056
rect 216642 236000 216647 236056
rect 213545 235998 216647 236000
rect 213545 235995 213611 235998
rect 215385 235995 215451 235998
rect 216581 235995 216647 235998
rect 224350 235996 224356 236060
rect 224420 236058 224426 236060
rect 224769 236058 224835 236061
rect 224420 236056 224835 236058
rect 224420 236000 224774 236056
rect 224830 236000 224835 236056
rect 224420 235998 224835 236000
rect 224420 235996 224426 235998
rect 224769 235995 224835 235998
rect 235349 236058 235415 236061
rect 235574 236058 235580 236060
rect 235349 236056 235580 236058
rect 235349 236000 235354 236056
rect 235410 236000 235580 236056
rect 235349 235998 235580 236000
rect 235349 235995 235415 235998
rect 235574 235996 235580 235998
rect 235644 235996 235650 236060
rect 241697 236058 241763 236061
rect 247217 236060 247283 236061
rect 247769 236060 247835 236061
rect 250713 236060 250779 236061
rect 242750 236058 242756 236060
rect 241697 236056 242756 236058
rect 241697 236000 241702 236056
rect 241758 236000 242756 236056
rect 241697 235998 242756 236000
rect 241697 235995 241763 235998
rect 242750 235996 242756 235998
rect 242820 235996 242826 236060
rect 247166 235996 247172 236060
rect 247236 236058 247283 236060
rect 247718 236058 247724 236060
rect 247236 236056 247328 236058
rect 247278 236000 247328 236056
rect 247236 235998 247328 236000
rect 247678 235998 247724 236058
rect 247788 236056 247835 236060
rect 250662 236058 250668 236060
rect 247830 236000 247835 236056
rect 247236 235996 247283 235998
rect 247718 235996 247724 235998
rect 247788 235996 247835 236000
rect 250622 235998 250668 236058
rect 250732 236056 250779 236060
rect 250774 236000 250779 236056
rect 250662 235996 250668 235998
rect 250732 235996 250779 236000
rect 247217 235995 247283 235996
rect 247769 235995 247835 235996
rect 250713 235995 250779 235996
rect 294045 236058 294111 236061
rect 295057 236058 295123 236061
rect 294045 236056 295123 236058
rect 294045 236000 294050 236056
rect 294106 236000 295062 236056
rect 295118 236000 295123 236056
rect 294045 235998 295123 236000
rect 294045 235995 294111 235998
rect 295057 235995 295123 235998
rect 213637 235922 213703 235925
rect 235993 235922 236059 235925
rect 213637 235920 236059 235922
rect 213637 235864 213642 235920
rect 213698 235864 235998 235920
rect 236054 235864 236059 235920
rect 213637 235862 236059 235864
rect 213637 235859 213703 235862
rect 235993 235859 236059 235862
rect 241145 235922 241211 235925
rect 241881 235922 241947 235925
rect 241145 235920 241947 235922
rect 241145 235864 241150 235920
rect 241206 235864 241886 235920
rect 241942 235864 241947 235920
rect 241145 235862 241947 235864
rect 241145 235859 241211 235862
rect 241881 235859 241947 235862
rect 267457 235922 267523 235925
rect 331397 235922 331463 235925
rect 267457 235920 331463 235922
rect 267457 235864 267462 235920
rect 267518 235864 331402 235920
rect 331458 235864 331463 235920
rect 267457 235862 331463 235864
rect 267457 235859 267523 235862
rect 331397 235859 331463 235862
rect 241881 235786 241947 235789
rect 242566 235786 242572 235788
rect 241881 235784 242572 235786
rect 241881 235728 241886 235784
rect 241942 235728 242572 235784
rect 241881 235726 242572 235728
rect 241881 235723 241947 235726
rect 242566 235724 242572 235726
rect 242636 235724 242642 235788
rect 229829 235650 229895 235653
rect 236310 235650 236316 235652
rect 229829 235648 236316 235650
rect 229829 235592 229834 235648
rect 229890 235592 236316 235648
rect 229829 235590 236316 235592
rect 229829 235587 229895 235590
rect 236310 235588 236316 235590
rect 236380 235588 236386 235652
rect 243261 235650 243327 235653
rect 243854 235650 243860 235652
rect 243261 235648 243860 235650
rect 243261 235592 243266 235648
rect 243322 235592 243860 235648
rect 243261 235590 243860 235592
rect 243261 235587 243327 235590
rect 243854 235588 243860 235590
rect 243924 235588 243930 235652
rect 162894 235452 162900 235516
rect 162964 235514 162970 235516
rect 182909 235514 182975 235517
rect 162964 235512 182975 235514
rect 162964 235456 182914 235512
rect 182970 235456 182975 235512
rect 162964 235454 182975 235456
rect 162964 235452 162970 235454
rect 182909 235451 182975 235454
rect 210877 235514 210943 235517
rect 233785 235514 233851 235517
rect 239673 235514 239739 235517
rect 210877 235512 239739 235514
rect 210877 235456 210882 235512
rect 210938 235456 233790 235512
rect 233846 235456 239678 235512
rect 239734 235456 239739 235512
rect 210877 235454 239739 235456
rect 210877 235451 210943 235454
rect 233785 235451 233851 235454
rect 239673 235451 239739 235454
rect 243905 235514 243971 235517
rect 244038 235514 244044 235516
rect 243905 235512 244044 235514
rect 243905 235456 243910 235512
rect 243966 235456 244044 235512
rect 243905 235454 244044 235456
rect 243905 235451 243971 235454
rect 244038 235452 244044 235454
rect 244108 235452 244114 235516
rect 176510 235316 176516 235380
rect 176580 235378 176586 235380
rect 213637 235378 213703 235381
rect 176580 235376 213703 235378
rect 176580 235320 213642 235376
rect 213698 235320 213703 235376
rect 176580 235318 213703 235320
rect 176580 235316 176586 235318
rect 213637 235315 213703 235318
rect 239029 235378 239095 235381
rect 239990 235378 239996 235380
rect 239029 235376 239996 235378
rect 239029 235320 239034 235376
rect 239090 235320 239996 235376
rect 239029 235318 239996 235320
rect 239029 235315 239095 235318
rect 239990 235316 239996 235318
rect 240060 235316 240066 235380
rect 240910 235316 240916 235380
rect 240980 235378 240986 235380
rect 259545 235378 259611 235381
rect 259729 235378 259795 235381
rect 240980 235376 259795 235378
rect 240980 235320 259550 235376
rect 259606 235320 259734 235376
rect 259790 235320 259795 235376
rect 240980 235318 259795 235320
rect 240980 235316 240986 235318
rect 259545 235315 259611 235318
rect 259729 235315 259795 235318
rect 159449 235242 159515 235245
rect 215661 235242 215727 235245
rect 159449 235240 215727 235242
rect 159449 235184 159454 235240
rect 159510 235184 215666 235240
rect 215722 235184 215727 235240
rect 159449 235182 215727 235184
rect 159449 235179 159515 235182
rect 215661 235179 215727 235182
rect 220445 235242 220511 235245
rect 266353 235242 266419 235245
rect 220445 235240 266419 235242
rect 220445 235184 220450 235240
rect 220506 235184 266358 235240
rect 266414 235184 266419 235240
rect 220445 235182 266419 235184
rect 220445 235179 220511 235182
rect 266353 235179 266419 235182
rect 267917 235242 267983 235245
rect 331305 235242 331371 235245
rect 267917 235240 331371 235242
rect 267917 235184 267922 235240
rect 267978 235184 331310 235240
rect 331366 235184 331371 235240
rect 267917 235182 331371 235184
rect 267917 235179 267983 235182
rect 331305 235179 331371 235182
rect 224861 235106 224927 235109
rect 239673 235108 239739 235109
rect 231894 235106 231900 235108
rect 224861 235104 231900 235106
rect 224861 235048 224866 235104
rect 224922 235048 231900 235104
rect 224861 235046 231900 235048
rect 224861 235043 224927 235046
rect 231894 235044 231900 235046
rect 231964 235044 231970 235108
rect 239622 235106 239628 235108
rect 239582 235046 239628 235106
rect 239692 235104 239739 235108
rect 243445 235108 243511 235109
rect 243445 235106 243492 235108
rect 239734 235048 239739 235104
rect 239622 235044 239628 235046
rect 239692 235044 239739 235048
rect 243400 235104 243492 235106
rect 243400 235048 243450 235104
rect 243400 235046 243492 235048
rect 239673 235043 239739 235044
rect 243445 235044 243492 235046
rect 243556 235044 243562 235108
rect 243445 235043 243511 235044
rect 259545 234970 259611 234973
rect 268469 234970 268535 234973
rect 259545 234968 268535 234970
rect 259545 234912 259550 234968
rect 259606 234912 268474 234968
rect 268530 234912 268535 234968
rect 259545 234910 268535 234912
rect 259545 234907 259611 234910
rect 268469 234907 268535 234910
rect 240869 234834 240935 234837
rect 241094 234834 241100 234836
rect 240869 234832 241100 234834
rect 240869 234776 240874 234832
rect 240930 234776 241100 234832
rect 240869 234774 241100 234776
rect 240869 234771 240935 234774
rect 241094 234772 241100 234774
rect 241164 234772 241170 234836
rect 255497 234834 255563 234837
rect 256049 234834 256115 234837
rect 268009 234834 268075 234837
rect 255497 234832 268075 234834
rect 255497 234776 255502 234832
rect 255558 234776 256054 234832
rect 256110 234776 268014 234832
rect 268070 234776 268075 234832
rect 255497 234774 268075 234776
rect 255497 234771 255563 234774
rect 256049 234771 256115 234774
rect 268009 234771 268075 234774
rect 234470 234636 234476 234700
rect 234540 234698 234546 234700
rect 249701 234698 249767 234701
rect 234540 234696 249767 234698
rect 234540 234640 249706 234696
rect 249762 234640 249767 234696
rect 234540 234638 249767 234640
rect 234540 234636 234546 234638
rect 249701 234635 249767 234638
rect 211061 234562 211127 234565
rect 242617 234562 242683 234565
rect 211061 234560 242683 234562
rect 211061 234504 211066 234560
rect 211122 234504 242622 234560
rect 242678 234504 242683 234560
rect 211061 234502 242683 234504
rect 211061 234499 211127 234502
rect 242617 234499 242683 234502
rect 255865 234562 255931 234565
rect 269941 234562 270007 234565
rect 255865 234560 270007 234562
rect 255865 234504 255870 234560
rect 255926 234504 269946 234560
rect 270002 234504 270007 234560
rect 255865 234502 270007 234504
rect 255865 234499 255931 234502
rect 269941 234499 270007 234502
rect 180374 234364 180380 234428
rect 180444 234426 180450 234428
rect 240133 234426 240199 234429
rect 180444 234424 240199 234426
rect 180444 234368 240138 234424
rect 240194 234368 240199 234424
rect 180444 234366 240199 234368
rect 180444 234364 180450 234366
rect 240133 234363 240199 234366
rect 256417 234426 256483 234429
rect 271781 234426 271847 234429
rect 256417 234424 271847 234426
rect 256417 234368 256422 234424
rect 256478 234368 271786 234424
rect 271842 234368 271847 234424
rect 256417 234366 271847 234368
rect 256417 234363 256483 234366
rect 271781 234363 271847 234366
rect 184422 234228 184428 234292
rect 184492 234290 184498 234292
rect 244181 234290 244247 234293
rect 268745 234290 268811 234293
rect 184492 234288 268811 234290
rect 184492 234232 244186 234288
rect 244242 234232 268750 234288
rect 268806 234232 268811 234288
rect 184492 234230 268811 234232
rect 184492 234228 184498 234230
rect 244181 234227 244247 234230
rect 268745 234227 268811 234230
rect 231853 234154 231919 234157
rect 250529 234154 250595 234157
rect 231853 234152 250595 234154
rect 231853 234096 231858 234152
rect 231914 234096 250534 234152
rect 250590 234096 250595 234152
rect 231853 234094 250595 234096
rect 231853 234091 231919 234094
rect 250529 234091 250595 234094
rect 252001 234154 252067 234157
rect 252185 234154 252251 234157
rect 312629 234154 312695 234157
rect 252001 234152 312695 234154
rect 252001 234096 252006 234152
rect 252062 234096 252190 234152
rect 252246 234096 312634 234152
rect 312690 234096 312695 234152
rect 252001 234094 312695 234096
rect 252001 234091 252067 234094
rect 252185 234091 252251 234094
rect 312629 234091 312695 234094
rect 181478 233956 181484 234020
rect 181548 234018 181554 234020
rect 239213 234018 239279 234021
rect 181548 234016 239279 234018
rect 181548 233960 239218 234016
rect 239274 233960 239279 234016
rect 181548 233958 239279 233960
rect 181548 233956 181554 233958
rect 239213 233955 239279 233958
rect 270125 234018 270191 234021
rect 278681 234018 278747 234021
rect 270125 234016 278747 234018
rect 270125 233960 270130 234016
rect 270186 233960 278686 234016
rect 278742 233960 278747 234016
rect 270125 233958 278747 233960
rect 270125 233955 270191 233958
rect 278681 233955 278747 233958
rect 180558 233820 180564 233884
rect 180628 233882 180634 233884
rect 240358 233882 240364 233884
rect 180628 233822 240364 233882
rect 180628 233820 180634 233822
rect 240358 233820 240364 233822
rect 240428 233820 240434 233884
rect 258257 233882 258323 233885
rect 287513 233882 287579 233885
rect 258257 233880 287579 233882
rect 258257 233824 258262 233880
rect 258318 233824 287518 233880
rect 287574 233824 287579 233880
rect 258257 233822 287579 233824
rect 258257 233819 258323 233822
rect 287513 233819 287579 233822
rect 182582 233684 182588 233748
rect 182652 233746 182658 233748
rect 210233 233746 210299 233749
rect 211061 233746 211127 233749
rect 182652 233744 211127 233746
rect 182652 233688 210238 233744
rect 210294 233688 211066 233744
rect 211122 233688 211127 233744
rect 182652 233686 211127 233688
rect 182652 233684 182658 233686
rect 210233 233683 210299 233686
rect 211061 233683 211127 233686
rect 263869 233746 263935 233749
rect 311525 233746 311591 233749
rect 263869 233744 311591 233746
rect 263869 233688 263874 233744
rect 263930 233688 311530 233744
rect 311586 233688 311591 233744
rect 263869 233686 311591 233688
rect 263869 233683 263935 233686
rect 311525 233683 311591 233686
rect 173566 233548 173572 233612
rect 173636 233610 173642 233612
rect 232814 233610 232820 233612
rect 173636 233550 232820 233610
rect 173636 233548 173642 233550
rect 232814 233548 232820 233550
rect 232884 233548 232890 233612
rect 258574 233548 258580 233612
rect 258644 233610 258650 233612
rect 261569 233610 261635 233613
rect 258644 233608 261635 233610
rect 258644 233552 261574 233608
rect 261630 233552 261635 233608
rect 258644 233550 261635 233552
rect 258644 233548 258650 233550
rect 261569 233547 261635 233550
rect 173014 233412 173020 233476
rect 173084 233474 173090 233476
rect 232262 233474 232268 233476
rect 173084 233414 232268 233474
rect 173084 233412 173090 233414
rect 232262 233412 232268 233414
rect 232332 233412 232338 233476
rect 257102 233412 257108 233476
rect 257172 233474 257178 233476
rect 257705 233474 257771 233477
rect 257172 233472 257771 233474
rect 257172 233416 257710 233472
rect 257766 233416 257771 233472
rect 257172 233414 257771 233416
rect 257172 233412 257178 233414
rect 257705 233411 257771 233414
rect 165470 233140 165476 233204
rect 165540 233202 165546 233204
rect 205541 233202 205607 233205
rect 229134 233202 229140 233204
rect 165540 233200 205607 233202
rect 165540 233144 205546 233200
rect 205602 233144 205607 233200
rect 165540 233142 205607 233144
rect 165540 233140 165546 233142
rect 205541 233139 205607 233142
rect 209730 233142 229140 233202
rect 154389 233066 154455 233069
rect 208117 233066 208183 233069
rect 209730 233066 209790 233142
rect 229134 233140 229140 233142
rect 229204 233140 229210 233204
rect 154389 233064 209790 233066
rect 154389 233008 154394 233064
rect 154450 233008 208122 233064
rect 208178 233008 209790 233064
rect 154389 233006 209790 233008
rect 252553 233066 252619 233069
rect 252686 233066 252692 233068
rect 252553 233064 252692 233066
rect 252553 233008 252558 233064
rect 252614 233008 252692 233064
rect 252553 233006 252692 233008
rect 154389 233003 154455 233006
rect 208117 233003 208183 233006
rect 252553 233003 252619 233006
rect 252686 233004 252692 233006
rect 252756 233004 252762 233068
rect 263133 233066 263199 233069
rect 334065 233066 334131 233069
rect 263133 233064 334131 233066
rect 263133 233008 263138 233064
rect 263194 233008 334070 233064
rect 334126 233008 334131 233064
rect 263133 233006 334131 233008
rect 263133 233003 263199 233006
rect 334065 233003 334131 233006
rect 191598 232868 191604 232932
rect 191668 232930 191674 232932
rect 251081 232930 251147 232933
rect 268653 232930 268719 232933
rect 191668 232928 268719 232930
rect 191668 232872 251086 232928
rect 251142 232872 268658 232928
rect 268714 232872 268719 232928
rect 191668 232870 268719 232872
rect 191668 232868 191674 232870
rect 251081 232867 251147 232870
rect 268653 232867 268719 232870
rect 174302 232732 174308 232796
rect 174372 232794 174378 232796
rect 234429 232794 234495 232797
rect 174372 232792 234495 232794
rect 174372 232736 234434 232792
rect 234490 232736 234495 232792
rect 174372 232734 234495 232736
rect 174372 232732 174378 232734
rect 234429 232731 234495 232734
rect 236085 232794 236151 232797
rect 237230 232794 237236 232796
rect 236085 232792 237236 232794
rect 236085 232736 236090 232792
rect 236146 232736 237236 232792
rect 236085 232734 237236 232736
rect 236085 232731 236151 232734
rect 237230 232732 237236 232734
rect 237300 232794 237306 232796
rect 274449 232794 274515 232797
rect 237300 232792 274515 232794
rect 237300 232736 274454 232792
rect 274510 232736 274515 232792
rect 237300 232734 274515 232736
rect 237300 232732 237306 232734
rect 274449 232731 274515 232734
rect 175038 232596 175044 232660
rect 175108 232658 175114 232660
rect 233877 232658 233943 232661
rect 175108 232656 233943 232658
rect 175108 232600 233882 232656
rect 233938 232600 233943 232656
rect 175108 232598 233943 232600
rect 175108 232596 175114 232598
rect 233877 232595 233943 232598
rect 251950 232596 251956 232660
rect 252020 232658 252026 232660
rect 343633 232658 343699 232661
rect 252020 232656 343699 232658
rect 252020 232600 343638 232656
rect 343694 232600 343699 232656
rect 252020 232598 343699 232600
rect 252020 232596 252026 232598
rect 343633 232595 343699 232598
rect 163814 232460 163820 232524
rect 163884 232522 163890 232524
rect 192477 232522 192543 232525
rect 163884 232520 192543 232522
rect 163884 232464 192482 232520
rect 192538 232464 192543 232520
rect 163884 232462 192543 232464
rect 163884 232460 163890 232462
rect 192477 232459 192543 232462
rect 193070 232460 193076 232524
rect 193140 232522 193146 232524
rect 252001 232522 252067 232525
rect 193140 232520 252067 232522
rect 193140 232464 252006 232520
rect 252062 232464 252067 232520
rect 193140 232462 252067 232464
rect 193140 232460 193146 232462
rect 252001 232459 252067 232462
rect 164734 232324 164740 232388
rect 164804 232386 164810 232388
rect 194317 232386 194383 232389
rect 164804 232384 194383 232386
rect 164804 232328 194322 232384
rect 194378 232328 194383 232384
rect 164804 232326 194383 232328
rect 164804 232324 164810 232326
rect 194317 232323 194383 232326
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 194358 231916 194364 231980
rect 194428 231978 194434 231980
rect 253381 231978 253447 231981
rect 253657 231978 253723 231981
rect 194428 231976 253723 231978
rect 194428 231920 253386 231976
rect 253442 231920 253662 231976
rect 253718 231920 253723 231976
rect 194428 231918 253723 231920
rect 194428 231916 194434 231918
rect 253381 231915 253447 231918
rect 253657 231915 253723 231918
rect 172278 231780 172284 231844
rect 172348 231842 172354 231844
rect 228817 231842 228883 231845
rect 230841 231844 230907 231845
rect 172348 231840 228883 231842
rect 172348 231784 228822 231840
rect 228878 231784 228883 231840
rect 172348 231782 228883 231784
rect 172348 231780 172354 231782
rect 228817 231779 228883 231782
rect 230790 231780 230796 231844
rect 230860 231842 230907 231844
rect 237925 231844 237991 231845
rect 230860 231840 230952 231842
rect 230902 231784 230952 231840
rect 230860 231782 230952 231784
rect 237925 231840 237972 231844
rect 238036 231842 238042 231844
rect 270677 231842 270743 231845
rect 237925 231784 237930 231840
rect 230860 231780 230907 231782
rect 230841 231779 230907 231780
rect 237925 231780 237972 231784
rect 238036 231782 238082 231842
rect 248370 231840 270743 231842
rect 248370 231784 270682 231840
rect 270738 231784 270743 231840
rect 248370 231782 270743 231784
rect 238036 231780 238042 231782
rect 237925 231779 237991 231780
rect 174670 231644 174676 231708
rect 174740 231706 174746 231708
rect 234286 231706 234292 231708
rect 174740 231646 234292 231706
rect 174740 231644 174746 231646
rect 234286 231644 234292 231646
rect 234356 231644 234362 231708
rect 166390 231508 166396 231572
rect 166460 231570 166466 231572
rect 226241 231570 226307 231573
rect 166460 231568 226307 231570
rect 166460 231512 226246 231568
rect 226302 231512 226307 231568
rect 166460 231510 226307 231512
rect 166460 231508 166466 231510
rect 226241 231507 226307 231510
rect 168230 231372 168236 231436
rect 168300 231434 168306 231436
rect 227713 231434 227779 231437
rect 168300 231432 227779 231434
rect 168300 231376 227718 231432
rect 227774 231376 227779 231432
rect 168300 231374 227779 231376
rect 168300 231372 168306 231374
rect 227713 231371 227779 231374
rect 166574 231236 166580 231300
rect 166644 231298 166650 231300
rect 226333 231298 226399 231301
rect 166644 231296 226399 231298
rect 166644 231240 226338 231296
rect 226394 231240 226399 231296
rect 166644 231238 226399 231240
rect 166644 231236 166650 231238
rect 226333 231235 226399 231238
rect 229001 231298 229067 231301
rect 239857 231298 239923 231301
rect 248370 231298 248430 231782
rect 270677 231779 270743 231782
rect 254485 231706 254551 231709
rect 258165 231706 258231 231709
rect 317454 231706 317460 231708
rect 254485 231704 317460 231706
rect 254485 231648 254490 231704
rect 254546 231648 258170 231704
rect 258226 231648 317460 231704
rect 254485 231646 317460 231648
rect 254485 231643 254551 231646
rect 258165 231643 258231 231646
rect 317454 231644 317460 231646
rect 317524 231644 317530 231708
rect 261753 231570 261819 231573
rect 296621 231570 296687 231573
rect 261753 231568 296687 231570
rect 261753 231512 261758 231568
rect 261814 231512 296626 231568
rect 296682 231512 296687 231568
rect 261753 231510 296687 231512
rect 261753 231507 261819 231510
rect 296621 231507 296687 231510
rect 277301 231434 277367 231437
rect 229001 231296 248430 231298
rect 229001 231240 229006 231296
rect 229062 231240 239862 231296
rect 239918 231240 248430 231296
rect 229001 231238 248430 231240
rect 253890 231432 277367 231434
rect 253890 231376 277306 231432
rect 277362 231376 277367 231432
rect 253890 231374 277367 231376
rect 229001 231235 229067 231238
rect 239857 231235 239923 231238
rect 165654 231100 165660 231164
rect 165724 231162 165730 231164
rect 226517 231162 226583 231165
rect 165724 231160 226583 231162
rect 165724 231104 226522 231160
rect 226578 231104 226583 231160
rect 165724 231102 226583 231104
rect 165724 231100 165730 231102
rect 226517 231099 226583 231102
rect 234061 231162 234127 231165
rect 250662 231162 250668 231164
rect 234061 231160 250668 231162
rect 234061 231104 234066 231160
rect 234122 231104 250668 231160
rect 234061 231102 250668 231104
rect 234061 231099 234127 231102
rect 250662 231100 250668 231102
rect 250732 231162 250738 231164
rect 253890 231162 253950 231374
rect 277301 231371 277367 231374
rect 267089 231298 267155 231301
rect 268561 231298 268627 231301
rect 327574 231298 327580 231300
rect 267089 231296 327580 231298
rect 267089 231240 267094 231296
rect 267150 231240 268566 231296
rect 268622 231240 327580 231296
rect 267089 231238 327580 231240
rect 267089 231235 267155 231238
rect 268561 231235 268627 231238
rect 327574 231236 327580 231238
rect 327644 231236 327650 231300
rect 250732 231102 253950 231162
rect 250732 231100 250738 231102
rect 176142 230964 176148 231028
rect 176212 231026 176218 231028
rect 227437 231026 227503 231029
rect 176212 231024 227503 231026
rect 176212 230968 227442 231024
rect 227498 230968 227503 231024
rect 176212 230966 227503 230968
rect 176212 230964 176218 230966
rect 227437 230963 227503 230966
rect 253841 230482 253907 230485
rect 264237 230482 264303 230485
rect 328821 230482 328887 230485
rect 253841 230480 253950 230482
rect 253841 230424 253846 230480
rect 253902 230424 253950 230480
rect 253841 230419 253950 230424
rect 264237 230480 328887 230482
rect 264237 230424 264242 230480
rect 264298 230424 328826 230480
rect 328882 230424 328887 230480
rect 264237 230422 328887 230424
rect 264237 230419 264303 230422
rect 328821 230419 328887 230422
rect 253890 230346 253950 230419
rect 255262 230346 255268 230348
rect 253890 230286 255268 230346
rect 255262 230284 255268 230286
rect 255332 230346 255338 230348
rect 283005 230346 283071 230349
rect 255332 230344 283071 230346
rect 255332 230288 283010 230344
rect 283066 230288 283071 230344
rect 255332 230286 283071 230288
rect 255332 230284 255338 230286
rect 283005 230283 283071 230286
rect 184606 230148 184612 230212
rect 184676 230210 184682 230212
rect 244457 230210 244523 230213
rect 184676 230208 244523 230210
rect 184676 230152 244462 230208
rect 244518 230152 244523 230208
rect 184676 230150 244523 230152
rect 184676 230148 184682 230150
rect 244457 230147 244523 230150
rect 264145 230210 264211 230213
rect 271270 230210 271276 230212
rect 264145 230208 271276 230210
rect 264145 230152 264150 230208
rect 264206 230152 271276 230208
rect 264145 230150 271276 230152
rect 264145 230147 264211 230150
rect 271270 230148 271276 230150
rect 271340 230148 271346 230212
rect 181294 230012 181300 230076
rect 181364 230074 181370 230076
rect 241973 230074 242039 230077
rect 181364 230072 242039 230074
rect 181364 230016 241978 230072
rect 242034 230016 242039 230072
rect 181364 230014 242039 230016
rect 181364 230012 181370 230014
rect 241973 230011 242039 230014
rect 248689 230074 248755 230077
rect 249006 230074 249012 230076
rect 248689 230072 249012 230074
rect 248689 230016 248694 230072
rect 248750 230016 249012 230072
rect 248689 230014 249012 230016
rect 248689 230011 248755 230014
rect 249006 230012 249012 230014
rect 249076 230012 249082 230076
rect 168782 229876 168788 229940
rect 168852 229938 168858 229940
rect 229553 229938 229619 229941
rect 168852 229936 229619 229938
rect 168852 229880 229558 229936
rect 229614 229880 229619 229936
rect 168852 229878 229619 229880
rect 168852 229876 168858 229878
rect 229553 229875 229619 229878
rect 255129 229938 255195 229941
rect 287697 229938 287763 229941
rect 327165 229938 327231 229941
rect 255129 229936 327231 229938
rect 255129 229880 255134 229936
rect 255190 229880 287702 229936
rect 287758 229880 327170 229936
rect 327226 229880 327231 229936
rect 255129 229878 327231 229880
rect 255129 229875 255195 229878
rect 287697 229875 287763 229878
rect 327165 229875 327231 229878
rect 168046 229740 168052 229804
rect 168116 229802 168122 229804
rect 228265 229802 228331 229805
rect 168116 229800 228331 229802
rect 168116 229744 228270 229800
rect 228326 229744 228331 229800
rect 168116 229742 228331 229744
rect 168116 229740 168122 229742
rect 228265 229739 228331 229742
rect 261477 229802 261543 229805
rect 290641 229802 290707 229805
rect 331213 229802 331279 229805
rect 261477 229800 331279 229802
rect 261477 229744 261482 229800
rect 261538 229744 290646 229800
rect 290702 229744 331218 229800
rect 331274 229744 331279 229800
rect 261477 229742 331279 229744
rect 261477 229739 261543 229742
rect 290641 229739 290707 229742
rect 331213 229739 331279 229742
rect 266721 228986 266787 228989
rect 266997 228986 267063 228989
rect 338246 228986 338252 228988
rect 266721 228984 338252 228986
rect 266721 228928 266726 228984
rect 266782 228928 267002 228984
rect 267058 228928 338252 228984
rect 266721 228926 338252 228928
rect 266721 228923 266787 228926
rect 266997 228923 267063 228926
rect 338246 228924 338252 228926
rect 338316 228924 338322 228988
rect 265709 228850 265775 228853
rect 330334 228850 330340 228852
rect 265709 228848 330340 228850
rect 265709 228792 265714 228848
rect 265770 228792 330340 228848
rect 265709 228790 330340 228792
rect 265709 228787 265775 228790
rect 330334 228788 330340 228790
rect 330404 228788 330410 228852
rect 246389 228714 246455 228717
rect 251173 228714 251239 228717
rect 310513 228714 310579 228717
rect 246389 228712 310579 228714
rect 246389 228656 246394 228712
rect 246450 228656 251178 228712
rect 251234 228656 310518 228712
rect 310574 228656 310579 228712
rect 246389 228654 310579 228656
rect 246389 228651 246455 228654
rect 251173 228651 251239 228654
rect 310513 228651 310579 228654
rect 181110 228516 181116 228580
rect 181180 228578 181186 228580
rect 240542 228578 240548 228580
rect 181180 228518 240548 228578
rect 181180 228516 181186 228518
rect 240542 228516 240548 228518
rect 240612 228516 240618 228580
rect 249742 228516 249748 228580
rect 249812 228578 249818 228580
rect 251030 228578 251036 228580
rect 249812 228518 251036 228578
rect 249812 228516 249818 228518
rect 251030 228516 251036 228518
rect 251100 228578 251106 228580
rect 309174 228578 309180 228580
rect 251100 228518 309180 228578
rect 251100 228516 251106 228518
rect 309174 228516 309180 228518
rect 309244 228516 309250 228580
rect 150249 228442 150315 228445
rect 225454 228442 225460 228444
rect 150249 228440 225460 228442
rect 150249 228384 150254 228440
rect 150310 228384 225460 228440
rect 150249 228382 225460 228384
rect 150249 228379 150315 228382
rect 225454 228380 225460 228382
rect 225524 228380 225530 228444
rect 292021 228442 292087 228445
rect 238710 228440 292087 228442
rect 238710 228384 292026 228440
rect 292082 228384 292087 228440
rect 238710 228382 292087 228384
rect 158345 228306 158411 228309
rect 235574 228306 235580 228308
rect 158345 228304 235580 228306
rect 158345 228248 158350 228304
rect 158406 228248 235580 228304
rect 158345 228246 235580 228248
rect 158345 228243 158411 228246
rect 235574 228244 235580 228246
rect 235644 228306 235650 228308
rect 238710 228306 238770 228382
rect 292021 228379 292087 228382
rect 235644 228246 238770 228306
rect 235644 228244 235650 228246
rect -960 227884 480 228124
rect 259126 227564 259132 227628
rect 259196 227626 259202 227628
rect 333973 227626 334039 227629
rect 259196 227624 334039 227626
rect 259196 227568 333978 227624
rect 334034 227568 334039 227624
rect 259196 227566 334039 227568
rect 259196 227564 259202 227566
rect 333973 227563 334039 227566
rect 236821 227490 236887 227493
rect 264697 227490 264763 227493
rect 236821 227488 264763 227490
rect 236821 227432 236826 227488
rect 236882 227432 264702 227488
rect 264758 227432 264763 227488
rect 236821 227430 264763 227432
rect 236821 227427 236887 227430
rect 264697 227427 264763 227430
rect 267181 227490 267247 227493
rect 330518 227490 330524 227492
rect 267181 227488 330524 227490
rect 267181 227432 267186 227488
rect 267242 227432 330524 227488
rect 267181 227430 330524 227432
rect 267181 227427 267247 227430
rect 330518 227428 330524 227430
rect 330588 227428 330594 227492
rect 248045 227354 248111 227357
rect 248270 227354 248276 227356
rect 248045 227352 248276 227354
rect 248045 227296 248050 227352
rect 248106 227296 248276 227352
rect 248045 227294 248276 227296
rect 248045 227291 248111 227294
rect 248270 227292 248276 227294
rect 248340 227354 248346 227356
rect 308489 227354 308555 227357
rect 248340 227352 308555 227354
rect 248340 227296 308494 227352
rect 308550 227296 308555 227352
rect 248340 227294 308555 227296
rect 248340 227292 248346 227294
rect 308489 227291 308555 227294
rect 264605 227218 264671 227221
rect 296345 227218 296411 227221
rect 264605 227216 296411 227218
rect 264605 227160 264610 227216
rect 264666 227160 296350 227216
rect 296406 227160 296411 227216
rect 264605 227158 296411 227160
rect 264605 227155 264671 227158
rect 296345 227155 296411 227158
rect 221641 227082 221707 227085
rect 249742 227082 249748 227084
rect 221641 227080 249748 227082
rect 221641 227024 221646 227080
rect 221702 227024 249748 227080
rect 221641 227022 249748 227024
rect 221641 227019 221707 227022
rect 249742 227020 249748 227022
rect 249812 227020 249818 227084
rect 183134 226884 183140 226948
rect 183204 226946 183210 226948
rect 243445 226946 243511 226949
rect 183204 226944 243511 226946
rect 183204 226888 243450 226944
rect 243506 226888 243511 226944
rect 183204 226886 243511 226888
rect 183204 226884 183210 226886
rect 243445 226883 243511 226886
rect 259085 226404 259151 226405
rect 259085 226400 259132 226404
rect 259196 226402 259202 226404
rect 259085 226344 259090 226400
rect 259085 226340 259132 226344
rect 259196 226342 259242 226402
rect 259196 226340 259202 226342
rect 259085 226339 259151 226340
rect 227253 226266 227319 226269
rect 232773 226266 232839 226269
rect 269757 226266 269823 226269
rect 227253 226264 269823 226266
rect 227253 226208 227258 226264
rect 227314 226208 232778 226264
rect 232834 226208 269762 226264
rect 269818 226208 269823 226264
rect 227253 226206 269823 226208
rect 227253 226203 227319 226206
rect 232773 226203 232839 226206
rect 269757 226203 269823 226206
rect 247217 226130 247283 226133
rect 306414 226130 306420 226132
rect 247217 226128 306420 226130
rect 247217 226072 247222 226128
rect 247278 226072 306420 226128
rect 247217 226070 306420 226072
rect 247217 226067 247283 226070
rect 306414 226068 306420 226070
rect 306484 226068 306490 226132
rect 254894 225932 254900 225996
rect 254964 225994 254970 225996
rect 258717 225994 258783 225997
rect 254964 225992 258783 225994
rect 254964 225936 258722 225992
rect 258778 225936 258783 225992
rect 254964 225934 258783 225936
rect 254964 225932 254970 225934
rect 258717 225931 258783 225934
rect 261702 225932 261708 225996
rect 261772 225994 261778 225996
rect 312537 225994 312603 225997
rect 261772 225992 312603 225994
rect 261772 225936 312542 225992
rect 312598 225936 312603 225992
rect 261772 225934 312603 225936
rect 261772 225932 261778 225934
rect 312537 225931 312603 225934
rect 260414 225796 260420 225860
rect 260484 225858 260490 225860
rect 327809 225858 327875 225861
rect 260484 225856 327875 225858
rect 260484 225800 327814 225856
rect 327870 225800 327875 225856
rect 260484 225798 327875 225800
rect 260484 225796 260490 225798
rect 327809 225795 327875 225798
rect 197118 225660 197124 225724
rect 197188 225722 197194 225724
rect 255630 225722 255636 225724
rect 197188 225662 255636 225722
rect 197188 225660 197194 225662
rect 255630 225660 255636 225662
rect 255700 225660 255706 225724
rect 188838 225524 188844 225588
rect 188908 225586 188914 225588
rect 248045 225586 248111 225589
rect 188908 225584 248111 225586
rect 188908 225528 248050 225584
rect 248106 225528 248111 225584
rect 188908 225526 248111 225528
rect 188908 225524 188914 225526
rect 248045 225523 248111 225526
rect 209681 224906 209747 224909
rect 224677 224906 224743 224909
rect 209681 224904 224743 224906
rect 209681 224848 209686 224904
rect 209742 224848 224682 224904
rect 224738 224848 224743 224904
rect 209681 224846 224743 224848
rect 209681 224843 209790 224846
rect 224677 224843 224743 224846
rect 234337 224906 234403 224909
rect 234470 224906 234476 224908
rect 234337 224904 234476 224906
rect 234337 224848 234342 224904
rect 234398 224848 234476 224904
rect 234337 224846 234476 224848
rect 234337 224843 234403 224846
rect 234470 224844 234476 224846
rect 234540 224906 234546 224908
rect 311341 224906 311407 224909
rect 234540 224904 311407 224906
rect 234540 224848 311346 224904
rect 311402 224848 311407 224904
rect 234540 224846 311407 224848
rect 234540 224844 234546 224846
rect 311341 224843 311407 224846
rect 167678 224300 167684 224364
rect 167748 224362 167754 224364
rect 209730 224362 209790 224843
rect 253381 224770 253447 224773
rect 313958 224770 313964 224772
rect 253381 224768 313964 224770
rect 253381 224712 253386 224768
rect 253442 224712 313964 224768
rect 253381 224710 313964 224712
rect 253381 224707 253447 224710
rect 313958 224708 313964 224710
rect 314028 224708 314034 224772
rect 316769 224634 316835 224637
rect 167748 224302 209790 224362
rect 258030 224632 316835 224634
rect 258030 224576 316774 224632
rect 316830 224576 316835 224632
rect 258030 224574 316835 224576
rect 167748 224300 167754 224302
rect 169334 224164 169340 224228
rect 169404 224226 169410 224228
rect 228081 224226 228147 224229
rect 169404 224224 228147 224226
rect 169404 224168 228086 224224
rect 228142 224168 228147 224224
rect 169404 224166 228147 224168
rect 169404 224164 169410 224166
rect 228081 224163 228147 224166
rect 228541 224226 228607 224229
rect 256969 224226 257035 224229
rect 258030 224226 258090 224574
rect 316769 224571 316835 224574
rect 228541 224224 258090 224226
rect 228541 224168 228546 224224
rect 228602 224168 256974 224224
rect 257030 224168 258090 224224
rect 228541 224166 258090 224168
rect 228541 224163 228607 224166
rect 256969 224163 257035 224166
rect 262078 223622 263610 223682
rect 260373 223546 260439 223549
rect 260598 223546 260604 223548
rect 260373 223544 260604 223546
rect 260373 223488 260378 223544
rect 260434 223488 260604 223544
rect 260373 223486 260604 223488
rect 260373 223483 260439 223486
rect 260598 223484 260604 223486
rect 260668 223546 260674 223548
rect 262078 223546 262138 223622
rect 260668 223486 262138 223546
rect 262213 223546 262279 223549
rect 263317 223546 263383 223549
rect 262213 223544 263383 223546
rect 262213 223488 262218 223544
rect 262274 223488 263322 223544
rect 263378 223488 263383 223544
rect 262213 223486 263383 223488
rect 263550 223546 263610 223622
rect 339493 223546 339559 223549
rect 263550 223544 339559 223546
rect 263550 223488 339498 223544
rect 339554 223488 339559 223544
rect 263550 223486 339559 223488
rect 260668 223484 260674 223486
rect 262213 223483 262279 223486
rect 263317 223483 263383 223486
rect 339493 223483 339559 223486
rect 252134 223348 252140 223412
rect 252204 223410 252210 223412
rect 252502 223410 252508 223412
rect 252204 223350 252508 223410
rect 252204 223348 252210 223350
rect 252502 223348 252508 223350
rect 252572 223410 252578 223412
rect 317413 223410 317479 223413
rect 252572 223408 317479 223410
rect 252572 223352 317418 223408
rect 317474 223352 317479 223408
rect 252572 223350 317479 223352
rect 252572 223348 252578 223350
rect 317413 223347 317479 223350
rect 263133 223274 263199 223277
rect 263358 223274 263364 223276
rect 263133 223272 263364 223274
rect 263133 223216 263138 223272
rect 263194 223216 263364 223272
rect 263133 223214 263364 223216
rect 263133 223211 263199 223214
rect 263358 223212 263364 223214
rect 263428 223274 263434 223276
rect 328453 223274 328519 223277
rect 263428 223272 328519 223274
rect 263428 223216 328458 223272
rect 328514 223216 328519 223272
rect 263428 223214 328519 223216
rect 263428 223212 263434 223214
rect 328453 223211 328519 223214
rect 263317 223138 263383 223141
rect 321502 223138 321508 223140
rect 263317 223136 321508 223138
rect 263317 223080 263322 223136
rect 263378 223080 321508 223136
rect 263317 223078 321508 223080
rect 263317 223075 263383 223078
rect 321502 223076 321508 223078
rect 321572 223076 321578 223140
rect 224217 223002 224283 223005
rect 235390 223002 235396 223004
rect 224217 223000 235396 223002
rect 224217 222944 224222 223000
rect 224278 222944 235396 223000
rect 224217 222942 235396 222944
rect 224217 222939 224283 222942
rect 235390 222940 235396 222942
rect 235460 223002 235466 223004
rect 289353 223002 289419 223005
rect 235460 223000 289419 223002
rect 235460 222944 289358 223000
rect 289414 222944 289419 223000
rect 235460 222942 289419 222944
rect 235460 222940 235466 222942
rect 289353 222939 289419 222942
rect 209589 222866 209655 222869
rect 214189 222866 214255 222869
rect 234838 222866 234844 222868
rect 209589 222864 234844 222866
rect 209589 222808 209594 222864
rect 209650 222808 214194 222864
rect 214250 222808 234844 222864
rect 209589 222806 234844 222808
rect 209589 222803 209655 222806
rect 214189 222803 214255 222806
rect 234838 222804 234844 222806
rect 234908 222804 234914 222868
rect 247769 222866 247835 222869
rect 252502 222866 252508 222868
rect 247769 222864 252508 222866
rect 247769 222808 247774 222864
rect 247830 222808 252508 222864
rect 247769 222806 252508 222808
rect 247769 222803 247835 222806
rect 252502 222804 252508 222806
rect 252572 222804 252578 222868
rect 298921 222866 298987 222869
rect 252878 222864 298987 222866
rect 252878 222808 298926 222864
rect 298982 222808 298987 222864
rect 252878 222806 298987 222808
rect 252502 222668 252508 222732
rect 252572 222730 252578 222732
rect 252878 222730 252938 222806
rect 298921 222803 298987 222806
rect 285397 222730 285463 222733
rect 252572 222670 252938 222730
rect 258030 222728 285463 222730
rect 258030 222672 285402 222728
rect 285458 222672 285463 222728
rect 258030 222670 285463 222672
rect 252572 222668 252578 222670
rect 249006 222532 249012 222596
rect 249076 222594 249082 222596
rect 249742 222594 249748 222596
rect 249076 222534 249748 222594
rect 249076 222532 249082 222534
rect 249742 222532 249748 222534
rect 249812 222594 249818 222596
rect 258030 222594 258090 222670
rect 285397 222667 285463 222670
rect 249812 222534 258090 222594
rect 249812 222532 249818 222534
rect 253473 222188 253539 222189
rect 253422 222124 253428 222188
rect 253492 222186 253539 222188
rect 339585 222186 339651 222189
rect 253492 222184 339651 222186
rect 253534 222128 339590 222184
rect 339646 222128 339651 222184
rect 253492 222126 339651 222128
rect 253492 222124 253539 222126
rect 253473 222123 253539 222124
rect 339585 222123 339651 222126
rect 258390 221988 258396 222052
rect 258460 222050 258466 222052
rect 259126 222050 259132 222052
rect 258460 221990 259132 222050
rect 258460 221988 258466 221990
rect 259126 221988 259132 221990
rect 259196 222050 259202 222052
rect 315573 222050 315639 222053
rect 259196 222048 315639 222050
rect 259196 221992 315578 222048
rect 315634 221992 315639 222048
rect 259196 221990 315639 221992
rect 259196 221988 259202 221990
rect 315573 221987 315639 221990
rect 249374 221852 249380 221916
rect 249444 221914 249450 221916
rect 286777 221914 286843 221917
rect 249444 221912 286843 221914
rect 249444 221856 286782 221912
rect 286838 221856 286843 221912
rect 249444 221854 286843 221856
rect 249444 221852 249450 221854
rect 286777 221851 286843 221854
rect 231209 221778 231275 221781
rect 252502 221778 252508 221780
rect 231209 221776 252508 221778
rect 231209 221720 231214 221776
rect 231270 221720 252508 221776
rect 231209 221718 252508 221720
rect 231209 221715 231275 221718
rect 252502 221716 252508 221718
rect 252572 221716 252578 221780
rect 257102 221716 257108 221780
rect 257172 221778 257178 221780
rect 257521 221778 257587 221781
rect 289445 221778 289511 221781
rect 257172 221776 289511 221778
rect 257172 221720 257526 221776
rect 257582 221720 289450 221776
rect 289506 221720 289511 221776
rect 257172 221718 289511 221720
rect 257172 221716 257178 221718
rect 257521 221715 257587 221718
rect 289445 221715 289511 221718
rect 224309 221642 224375 221645
rect 249742 221642 249748 221644
rect 224309 221640 249748 221642
rect 224309 221584 224314 221640
rect 224370 221584 249748 221640
rect 224309 221582 249748 221584
rect 224309 221579 224375 221582
rect 249742 221580 249748 221582
rect 249812 221580 249818 221644
rect 173198 221444 173204 221508
rect 173268 221506 173274 221508
rect 233785 221506 233851 221509
rect 173268 221504 233851 221506
rect 173268 221448 233790 221504
rect 233846 221448 233851 221504
rect 173268 221446 233851 221448
rect 173268 221444 173274 221446
rect 233785 221443 233851 221446
rect 251817 221098 251883 221101
rect 259126 221098 259132 221100
rect 251817 221096 259132 221098
rect 251817 221040 251822 221096
rect 251878 221040 259132 221096
rect 251817 221038 259132 221040
rect 251817 221035 251883 221038
rect 259126 221036 259132 221038
rect 259196 221036 259202 221100
rect 249190 220962 249196 220964
rect 249068 220902 249196 220962
rect 249190 220900 249196 220902
rect 249260 220962 249266 220964
rect 249260 220902 249810 220962
rect 249260 220900 249266 220902
rect 178534 220764 178540 220828
rect 178604 220826 178610 220828
rect 237465 220826 237531 220829
rect 249198 220826 249258 220900
rect 178604 220824 237531 220826
rect 178604 220768 237470 220824
rect 237526 220768 237531 220824
rect 178604 220766 237531 220768
rect 178604 220764 178610 220766
rect 237465 220763 237531 220766
rect 238710 220766 249258 220826
rect 249425 220826 249491 220829
rect 249558 220826 249564 220828
rect 249425 220824 249564 220826
rect 249425 220768 249430 220824
rect 249486 220768 249564 220824
rect 249425 220766 249564 220768
rect 223573 220690 223639 220693
rect 224350 220690 224356 220692
rect 223573 220688 224356 220690
rect 223573 220632 223578 220688
rect 223634 220632 224356 220688
rect 223573 220630 224356 220632
rect 223573 220627 223639 220630
rect 224350 220628 224356 220630
rect 224420 220628 224426 220692
rect 225965 220690 226031 220693
rect 238710 220690 238770 220766
rect 249425 220763 249491 220766
rect 249558 220764 249564 220766
rect 249628 220764 249634 220828
rect 249750 220826 249810 220902
rect 340873 220826 340939 220829
rect 249750 220824 340939 220826
rect 249750 220768 340878 220824
rect 340934 220768 340939 220824
rect 249750 220766 340939 220768
rect 225965 220688 238770 220690
rect 225965 220632 225970 220688
rect 226026 220632 238770 220688
rect 225965 220630 238770 220632
rect 249566 220690 249626 220764
rect 340873 220763 340939 220766
rect 309726 220690 309732 220692
rect 249566 220630 309732 220690
rect 225965 220627 226031 220630
rect 309726 220628 309732 220630
rect 309796 220628 309802 220692
rect 246982 220492 246988 220556
rect 247052 220554 247058 220556
rect 247718 220554 247724 220556
rect 247052 220494 247724 220554
rect 247052 220492 247058 220494
rect 247718 220492 247724 220494
rect 247788 220554 247794 220556
rect 307702 220554 307708 220556
rect 247788 220494 307708 220554
rect 247788 220492 247794 220494
rect 307702 220492 307708 220494
rect 307772 220492 307778 220556
rect 235349 220418 235415 220421
rect 252277 220418 252343 220421
rect 310830 220418 310836 220420
rect 235349 220416 310836 220418
rect 235349 220360 235354 220416
rect 235410 220360 252282 220416
rect 252338 220360 310836 220416
rect 235349 220358 310836 220360
rect 235349 220355 235415 220358
rect 252277 220355 252343 220358
rect 310830 220356 310836 220358
rect 310900 220356 310906 220420
rect 169150 220220 169156 220284
rect 169220 220282 169226 220284
rect 228449 220282 228515 220285
rect 169220 220280 228515 220282
rect 169220 220224 228454 220280
rect 228510 220224 228515 220280
rect 169220 220222 228515 220224
rect 169220 220220 169226 220222
rect 228449 220219 228515 220222
rect 229921 220282 229987 220285
rect 246982 220282 246988 220284
rect 229921 220280 246988 220282
rect 229921 220224 229926 220280
rect 229982 220224 246988 220280
rect 229921 220222 246988 220224
rect 229921 220219 229987 220222
rect 246982 220220 246988 220222
rect 247052 220220 247058 220284
rect 256509 220282 256575 220285
rect 314694 220282 314700 220284
rect 256509 220280 314700 220282
rect 256509 220224 256514 220280
rect 256570 220224 314700 220280
rect 256509 220222 314700 220224
rect 256509 220219 256575 220222
rect 314694 220220 314700 220222
rect 314764 220220 314770 220284
rect 163630 220084 163636 220148
rect 163700 220146 163706 220148
rect 223665 220146 223731 220149
rect 163700 220144 223731 220146
rect 163700 220088 223670 220144
rect 223726 220088 223731 220144
rect 163700 220086 223731 220088
rect 163700 220084 163706 220086
rect 223665 220083 223731 220086
rect 239489 220146 239555 220149
rect 255446 220146 255452 220148
rect 239489 220144 255452 220146
rect 239489 220088 239494 220144
rect 239550 220088 255452 220144
rect 239489 220086 255452 220088
rect 239489 220083 239555 220086
rect 255446 220084 255452 220086
rect 255516 220146 255522 220148
rect 313774 220146 313780 220148
rect 255516 220086 313780 220146
rect 255516 220084 255522 220086
rect 313774 220084 313780 220086
rect 313844 220084 313850 220148
rect 254117 220010 254183 220013
rect 291694 220010 291700 220012
rect 254117 220008 291700 220010
rect 254117 219952 254122 220008
rect 254178 219952 291700 220008
rect 254117 219950 291700 219952
rect 254117 219947 254183 219950
rect 291694 219948 291700 219950
rect 291764 219948 291770 220012
rect 206737 219330 206803 219333
rect 224585 219330 224651 219333
rect 206737 219328 224651 219330
rect 206737 219272 206742 219328
rect 206798 219272 224590 219328
rect 224646 219272 224651 219328
rect 206737 219270 224651 219272
rect 206737 219267 206803 219270
rect 224585 219267 224651 219270
rect 242198 219268 242204 219332
rect 242268 219330 242274 219332
rect 301446 219330 301452 219332
rect 242268 219270 301452 219330
rect 242268 219268 242274 219270
rect 301446 219268 301452 219270
rect 301516 219268 301522 219332
rect 243854 219132 243860 219196
rect 243924 219194 243930 219196
rect 302918 219194 302924 219196
rect 243924 219134 302924 219194
rect 243924 219132 243930 219134
rect 302918 219132 302924 219134
rect 302988 219132 302994 219196
rect 182950 218996 182956 219060
rect 183020 219058 183026 219060
rect 242249 219058 242315 219061
rect 183020 219056 242315 219058
rect 183020 219000 242254 219056
rect 242310 219000 242315 219056
rect 183020 218998 242315 219000
rect 183020 218996 183026 218998
rect 242249 218995 242315 218998
rect 244038 218996 244044 219060
rect 244108 219058 244114 219060
rect 302734 219058 302740 219060
rect 244108 218998 302740 219058
rect 244108 218996 244114 218998
rect 302734 218996 302740 218998
rect 302804 218996 302810 219060
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 165102 218860 165108 218924
rect 165172 218922 165178 218924
rect 206737 218922 206803 218925
rect 165172 218920 206803 218922
rect 165172 218864 206742 218920
rect 206798 218864 206803 218920
rect 165172 218862 206803 218864
rect 165172 218860 165178 218862
rect 206737 218859 206803 218862
rect 237966 218860 237972 218924
rect 238036 218922 238042 218924
rect 296846 218922 296852 218924
rect 238036 218862 296852 218922
rect 238036 218860 238042 218862
rect 296846 218860 296852 218862
rect 296916 218860 296922 218924
rect 583520 218908 584960 218998
rect 167862 218724 167868 218788
rect 167932 218786 167938 218788
rect 227621 218786 227687 218789
rect 167932 218784 227687 218786
rect 167932 218728 227626 218784
rect 227682 218728 227687 218784
rect 167932 218726 227687 218728
rect 167932 218724 167938 218726
rect 227621 218723 227687 218726
rect 242249 218786 242315 218789
rect 299606 218786 299612 218788
rect 242249 218784 299612 218786
rect 242249 218728 242254 218784
rect 242310 218728 299612 218784
rect 242249 218726 299612 218728
rect 242249 218723 242315 218726
rect 299606 218724 299612 218726
rect 299676 218724 299682 218788
rect 164918 218588 164924 218652
rect 164988 218650 164994 218652
rect 225413 218650 225479 218653
rect 164988 218648 225479 218650
rect 164988 218592 225418 218648
rect 225474 218592 225479 218648
rect 164988 218590 225479 218592
rect 164988 218588 164994 218590
rect 225413 218587 225479 218590
rect 239990 218588 239996 218652
rect 240060 218650 240066 218652
rect 296161 218650 296227 218653
rect 240060 218648 296227 218650
rect 240060 218592 296166 218648
rect 296222 218592 296227 218648
rect 240060 218590 296227 218592
rect 240060 218588 240066 218590
rect 296161 218587 296227 218590
rect 243997 218244 244063 218245
rect 243997 218240 244044 218244
rect 244108 218242 244114 218244
rect 243997 218184 244002 218240
rect 243997 218180 244044 218184
rect 244108 218182 244154 218242
rect 244108 218180 244114 218182
rect 243997 218179 244063 218180
rect 239949 218108 240015 218109
rect 243813 218108 243879 218109
rect 239949 218104 239996 218108
rect 240060 218106 240066 218108
rect 239949 218048 239954 218104
rect 239949 218044 239996 218048
rect 240060 218046 240106 218106
rect 243813 218104 243860 218108
rect 243924 218106 243930 218108
rect 243813 218048 243818 218104
rect 240060 218044 240066 218046
rect 243813 218044 243860 218048
rect 243924 218046 243970 218106
rect 243924 218044 243930 218046
rect 239949 218043 240015 218044
rect 243813 218043 243879 218044
rect 229645 217970 229711 217973
rect 230381 217970 230447 217973
rect 288433 217970 288499 217973
rect 229645 217968 288499 217970
rect 229645 217912 229650 217968
rect 229706 217912 230386 217968
rect 230442 217912 288438 217968
rect 288494 217912 288499 217968
rect 229645 217910 288499 217912
rect 229645 217907 229711 217910
rect 230381 217907 230447 217910
rect 288433 217907 288499 217910
rect 170990 217772 170996 217836
rect 171060 217834 171066 217836
rect 230841 217834 230907 217837
rect 284937 217834 285003 217837
rect 171060 217832 285003 217834
rect 171060 217776 230846 217832
rect 230902 217776 284942 217832
rect 284998 217776 285003 217832
rect 171060 217774 285003 217776
rect 171060 217772 171066 217774
rect 230841 217771 230907 217774
rect 284937 217771 285003 217774
rect 168966 217636 168972 217700
rect 169036 217698 169042 217700
rect 229645 217698 229711 217701
rect 169036 217696 229711 217698
rect 169036 217640 229650 217696
rect 229706 217640 229711 217696
rect 169036 217638 229711 217640
rect 169036 217636 169042 217638
rect 229645 217635 229711 217638
rect 171726 217500 171732 217564
rect 171796 217562 171802 217564
rect 231945 217562 232011 217565
rect 171796 217560 232011 217562
rect 171796 217504 231950 217560
rect 232006 217504 232011 217560
rect 171796 217502 232011 217504
rect 171796 217500 171802 217502
rect 231945 217499 232011 217502
rect 170622 217364 170628 217428
rect 170692 217426 170698 217428
rect 231393 217426 231459 217429
rect 170692 217424 231459 217426
rect 170692 217368 231398 217424
rect 231454 217368 231459 217424
rect 170692 217366 231459 217368
rect 170692 217364 170698 217366
rect 231393 217363 231459 217366
rect 171910 217228 171916 217292
rect 171980 217290 171986 217292
rect 233049 217290 233115 217293
rect 171980 217288 233115 217290
rect 171980 217232 233054 217288
rect 233110 217232 233115 217288
rect 171980 217230 233115 217232
rect 171980 217228 171986 217230
rect 233049 217227 233115 217230
rect 172094 217092 172100 217156
rect 172164 217154 172170 217156
rect 230473 217154 230539 217157
rect 172164 217152 230539 217154
rect 172164 217096 230478 217152
rect 230534 217096 230539 217152
rect 172164 217094 230539 217096
rect 172164 217092 172170 217094
rect 230473 217091 230539 217094
rect 170806 216956 170812 217020
rect 170876 217018 170882 217020
rect 229277 217018 229343 217021
rect 170876 217016 229343 217018
rect 170876 216960 229282 217016
rect 229338 216960 229343 217016
rect 170876 216958 229343 216960
rect 170876 216956 170882 216958
rect 229277 216955 229343 216958
rect 259361 216610 259427 216613
rect 318926 216610 318932 216612
rect 259361 216608 318932 216610
rect 259361 216552 259366 216608
rect 259422 216552 318932 216608
rect 259361 216550 318932 216552
rect 259361 216547 259427 216550
rect 318926 216548 318932 216550
rect 318996 216548 319002 216612
rect 230974 216412 230980 216476
rect 231044 216474 231050 216476
rect 290733 216474 290799 216477
rect 231044 216472 290799 216474
rect 231044 216416 290738 216472
rect 290794 216416 290799 216472
rect 231044 216414 290799 216416
rect 231044 216412 231050 216414
rect 290733 216411 290799 216414
rect 259310 216276 259316 216340
rect 259380 216338 259386 216340
rect 290549 216338 290615 216341
rect 259380 216336 290615 216338
rect 259380 216280 290554 216336
rect 290610 216280 290615 216336
rect 259380 216278 290615 216280
rect 259380 216276 259386 216278
rect 290549 216275 290615 216278
rect 258073 215522 258139 215525
rect 259361 215522 259427 215525
rect 258073 215520 259427 215522
rect 258073 215464 258078 215520
rect 258134 215464 259366 215520
rect 259422 215464 259427 215520
rect 258073 215462 259427 215464
rect 258073 215459 258139 215462
rect 259361 215459 259427 215462
rect 258809 215386 258875 215389
rect 259310 215386 259316 215388
rect 258809 215384 259316 215386
rect 258809 215328 258814 215384
rect 258870 215328 259316 215384
rect 258809 215326 259316 215328
rect 258809 215323 258875 215326
rect 259310 215324 259316 215326
rect 259380 215324 259386 215388
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 196934 214916 196940 214980
rect 197004 214978 197010 214980
rect 255814 214978 255820 214980
rect 197004 214918 255820 214978
rect 197004 214916 197010 214918
rect 255814 214916 255820 214918
rect 255884 214916 255890 214980
rect 195646 214780 195652 214844
rect 195716 214842 195722 214844
rect 255129 214842 255195 214845
rect 195716 214840 255195 214842
rect 195716 214784 255134 214840
rect 255190 214784 255195 214840
rect 195716 214782 255195 214784
rect 195716 214780 195722 214782
rect 255129 214779 255195 214782
rect 195830 214644 195836 214708
rect 195900 214706 195906 214708
rect 255313 214706 255379 214709
rect 195900 214704 255379 214706
rect 195900 214648 255318 214704
rect 255374 214648 255379 214704
rect 195900 214646 255379 214648
rect 195900 214644 195906 214646
rect 255313 214643 255379 214646
rect 170438 214508 170444 214572
rect 170508 214570 170514 214572
rect 230197 214570 230263 214573
rect 170508 214568 230263 214570
rect 170508 214512 230202 214568
rect 230258 214512 230263 214568
rect 170508 214510 230263 214512
rect 170508 214508 170514 214510
rect 230197 214507 230263 214510
rect 179086 213828 179092 213892
rect 179156 213890 179162 213892
rect 237373 213890 237439 213893
rect 179156 213888 237439 213890
rect 179156 213832 237378 213888
rect 237434 213832 237439 213888
rect 179156 213830 237439 213832
rect 179156 213828 179162 213830
rect 237373 213827 237439 213830
rect 178902 213692 178908 213756
rect 178972 213754 178978 213756
rect 238477 213754 238543 213757
rect 178972 213752 238543 213754
rect 178972 213696 238482 213752
rect 238538 213696 238543 213752
rect 178972 213694 238543 213696
rect 178972 213692 178978 213694
rect 238477 213691 238543 213694
rect 185158 213556 185164 213620
rect 185228 213618 185234 213620
rect 244406 213618 244412 213620
rect 185228 213558 244412 213618
rect 185228 213556 185234 213558
rect 244406 213556 244412 213558
rect 244476 213556 244482 213620
rect 180190 213420 180196 213484
rect 180260 213482 180266 213484
rect 239438 213482 239444 213484
rect 180260 213422 239444 213482
rect 180260 213420 180266 213422
rect 239438 213420 239444 213422
rect 239508 213420 239514 213484
rect 182766 213284 182772 213348
rect 182836 213346 182842 213348
rect 243813 213346 243879 213349
rect 182836 213344 243879 213346
rect 182836 213288 243818 213344
rect 243874 213288 243879 213344
rect 182836 213286 243879 213288
rect 182836 213284 182842 213286
rect 243813 213283 243879 213286
rect 174486 213148 174492 213212
rect 174556 213210 174562 213212
rect 234981 213210 235047 213213
rect 174556 213208 235047 213210
rect 174556 213152 234986 213208
rect 235042 213152 235047 213208
rect 174556 213150 235047 213152
rect 174556 213148 174562 213150
rect 234981 213147 235047 213150
rect 180006 213012 180012 213076
rect 180076 213074 180082 213076
rect 238845 213074 238911 213077
rect 180076 213072 238911 213074
rect 180076 213016 238850 213072
rect 238906 213016 238911 213072
rect 180076 213014 238911 213016
rect 180076 213012 180082 213014
rect 238845 213011 238911 213014
rect 164325 212122 164391 212125
rect 166901 212122 166967 212125
rect 203190 212122 203196 212124
rect 164325 212120 203196 212122
rect 164325 212064 164330 212120
rect 164386 212064 166906 212120
rect 166962 212064 203196 212120
rect 164325 212062 203196 212064
rect 164325 212059 164391 212062
rect 166901 212059 166967 212062
rect 203190 212060 203196 212062
rect 203260 212060 203266 212124
rect 180926 211924 180932 211988
rect 180996 211986 181002 211988
rect 239949 211986 240015 211989
rect 180996 211984 240015 211986
rect 180996 211928 239954 211984
rect 240010 211928 240015 211984
rect 180996 211926 240015 211928
rect 180996 211924 181002 211926
rect 239949 211923 240015 211926
rect 178718 211788 178724 211852
rect 178788 211850 178794 211852
rect 238753 211850 238819 211853
rect 178788 211848 238819 211850
rect 178788 211792 238758 211848
rect 238814 211792 238819 211848
rect 178788 211790 238819 211792
rect 178788 211788 178794 211790
rect 238753 211787 238819 211790
rect 198406 210428 198412 210492
rect 198476 210490 198482 210492
rect 257521 210490 257587 210493
rect 198476 210488 257587 210490
rect 198476 210432 257526 210488
rect 257582 210432 257587 210488
rect 198476 210430 257587 210432
rect 198476 210428 198482 210430
rect 257521 210427 257587 210430
rect 190310 210292 190316 210356
rect 190380 210354 190386 210356
rect 249425 210354 249491 210357
rect 190380 210352 249491 210354
rect 190380 210296 249430 210352
rect 249486 210296 249491 210352
rect 190380 210294 249491 210296
rect 190380 210292 190386 210294
rect 249425 210291 249491 210294
rect 182541 210082 182607 210085
rect 182541 210080 182650 210082
rect 182541 210024 182546 210080
rect 182602 210024 182650 210080
rect 182541 210019 182650 210024
rect 198038 210020 198044 210084
rect 198108 210082 198114 210084
rect 198641 210082 198707 210085
rect 198108 210080 198707 210082
rect 198108 210024 198646 210080
rect 198702 210024 198707 210080
rect 198108 210022 198707 210024
rect 198108 210020 198114 210022
rect 198641 210019 198707 210022
rect 169753 209946 169819 209949
rect 170397 209946 170463 209949
rect 169753 209944 170463 209946
rect 169753 209888 169758 209944
rect 169814 209888 170402 209944
rect 170458 209888 170463 209944
rect 169753 209886 170463 209888
rect 169753 209883 169819 209886
rect 170397 209883 170463 209886
rect 182590 209674 182650 210019
rect 199326 209748 199332 209812
rect 199396 209810 199402 209812
rect 199929 209810 199995 209813
rect 199396 209808 199995 209810
rect 199396 209752 199934 209808
rect 199990 209752 199995 209808
rect 199396 209750 199995 209752
rect 199396 209748 199402 209750
rect 199929 209747 199995 209750
rect 218513 209674 218579 209677
rect 182590 209672 218579 209674
rect 182590 209616 218518 209672
rect 218574 209616 218579 209672
rect 182590 209614 218579 209616
rect 218513 209611 218579 209614
rect 163446 209476 163452 209540
rect 163516 209538 163522 209540
rect 164141 209538 164207 209541
rect 163516 209536 164207 209538
rect 163516 209480 164146 209536
rect 164202 209480 164207 209536
rect 163516 209478 164207 209480
rect 163516 209476 163522 209478
rect 164141 209475 164207 209478
rect 184054 209476 184060 209540
rect 184124 209538 184130 209540
rect 184841 209538 184907 209541
rect 189533 209540 189599 209541
rect 189533 209538 189580 209540
rect 184124 209536 184907 209538
rect 184124 209480 184846 209536
rect 184902 209480 184907 209536
rect 184124 209478 184907 209480
rect 189488 209536 189580 209538
rect 189488 209480 189538 209536
rect 189488 209478 189580 209480
rect 184124 209476 184130 209478
rect 184841 209475 184907 209478
rect 189533 209476 189580 209478
rect 189644 209476 189650 209540
rect 193806 209476 193812 209540
rect 193876 209538 193882 209540
rect 194409 209538 194475 209541
rect 193876 209536 194475 209538
rect 193876 209480 194414 209536
rect 194470 209480 194475 209536
rect 193876 209478 194475 209480
rect 193876 209476 193882 209478
rect 189533 209475 189599 209476
rect 194409 209475 194475 209478
rect 195462 209476 195468 209540
rect 195532 209538 195538 209540
rect 195881 209538 195947 209541
rect 195532 209536 195947 209538
rect 195532 209480 195886 209536
rect 195942 209480 195947 209536
rect 195532 209478 195947 209480
rect 195532 209476 195538 209478
rect 195881 209475 195947 209478
rect 197854 209476 197860 209540
rect 197924 209538 197930 209540
rect 198457 209538 198523 209541
rect 199193 209540 199259 209541
rect 199142 209538 199148 209540
rect 197924 209536 198523 209538
rect 197924 209480 198462 209536
rect 198518 209480 198523 209536
rect 197924 209478 198523 209480
rect 199102 209478 199148 209538
rect 199212 209536 199259 209540
rect 199837 209540 199903 209541
rect 199837 209538 199884 209540
rect 199254 209480 199259 209536
rect 197924 209476 197930 209478
rect 198457 209475 198523 209478
rect 199142 209476 199148 209478
rect 199212 209476 199259 209480
rect 199792 209536 199884 209538
rect 199792 209480 199842 209536
rect 199792 209478 199884 209480
rect 199193 209475 199259 209476
rect 199837 209476 199884 209478
rect 199948 209476 199954 209540
rect 204253 209538 204319 209541
rect 204253 209536 204362 209538
rect 204253 209480 204258 209536
rect 204314 209480 204362 209536
rect 199837 209475 199903 209476
rect 204253 209475 204362 209480
rect 204302 209266 204362 209475
rect 205541 209266 205607 209269
rect 195930 209264 205607 209266
rect 195930 209208 205546 209264
rect 205602 209208 205607 209264
rect 195930 209206 205607 209208
rect 146937 209130 147003 209133
rect 195930 209130 195990 209206
rect 205541 209203 205607 209206
rect 146937 209128 195990 209130
rect 146937 209072 146942 209128
rect 146998 209072 195990 209128
rect 146937 209070 195990 209072
rect 218513 209130 218579 209133
rect 580717 209130 580783 209133
rect 218513 209128 580783 209130
rect 218513 209072 218518 209128
rect 218574 209072 580722 209128
rect 580778 209072 580783 209128
rect 218513 209070 580783 209072
rect 146937 209067 147003 209070
rect 218513 209067 218579 209070
rect 580717 209067 580783 209070
rect 189574 208932 189580 208996
rect 189644 208994 189650 208996
rect 580533 208994 580599 208997
rect 189644 208992 580599 208994
rect 189644 208936 580538 208992
rect 580594 208936 580599 208992
rect 189644 208934 580599 208936
rect 189644 208932 189650 208934
rect 580533 208931 580599 208934
rect 201350 207572 201356 207636
rect 201420 207634 201426 207636
rect 260373 207634 260439 207637
rect 201420 207632 260439 207634
rect 201420 207576 260378 207632
rect 260434 207576 260439 207632
rect 201420 207574 260439 207576
rect 201420 207572 201426 207574
rect 260373 207571 260439 207574
rect 203190 206212 203196 206276
rect 203260 206274 203266 206276
rect 580349 206274 580415 206277
rect 203260 206272 580415 206274
rect 203260 206216 580354 206272
rect 580410 206216 580415 206272
rect 203260 206214 580415 206216
rect 203260 206212 203266 206214
rect 580349 206211 580415 206214
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 583520 205580 584960 205670
rect 208894 204852 208900 204916
rect 208964 204914 208970 204916
rect 267181 204914 267247 204917
rect 208964 204912 267247 204914
rect 208964 204856 267186 204912
rect 267242 204856 267247 204912
rect 208964 204854 267247 204856
rect 208964 204852 208970 204854
rect 267181 204851 267247 204854
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 207841 188322 207907 188325
rect 231301 188322 231367 188325
rect 207841 188320 231367 188322
rect 207841 188264 207846 188320
rect 207902 188264 231306 188320
rect 231362 188264 231367 188320
rect 207841 188262 231367 188264
rect 207841 188259 207907 188262
rect 231301 188259 231367 188262
rect 207933 184242 207999 184245
rect 223941 184242 224007 184245
rect 207933 184240 224007 184242
rect 207933 184184 207938 184240
rect 207994 184184 223946 184240
rect 224002 184184 224007 184240
rect 207933 184182 224007 184184
rect 207933 184179 207999 184182
rect 223941 184179 224007 184182
rect 207790 182820 207796 182884
rect 207860 182882 207866 182884
rect 267457 182882 267523 182885
rect 207860 182880 267523 182882
rect 207860 182824 267462 182880
rect 267518 182824 267523 182880
rect 207860 182822 267523 182824
rect 207860 182820 207866 182822
rect 267457 182819 267523 182822
rect 205766 179964 205772 180028
rect 205836 180026 205842 180028
rect 265709 180026 265775 180029
rect 205836 180024 265775 180026
rect 205836 179968 265714 180024
rect 265770 179968 265775 180024
rect 205836 179966 265775 179968
rect 205836 179964 205842 179966
rect 265709 179963 265775 179966
rect 580441 179210 580507 179213
rect 583520 179210 584960 179300
rect 580441 179208 584960 179210
rect 580441 179152 580446 179208
rect 580502 179152 584960 179208
rect 580441 179150 584960 179152
rect 580441 179147 580507 179150
rect 583520 179060 584960 179150
rect 208025 176082 208091 176085
rect 261477 176082 261543 176085
rect 208025 176080 261543 176082
rect -960 175796 480 176036
rect 208025 176024 208030 176080
rect 208086 176024 261482 176080
rect 261538 176024 261543 176080
rect 208025 176022 261543 176024
rect 208025 176019 208091 176022
rect 261477 176019 261543 176022
rect 205950 175884 205956 175948
rect 206020 175946 206026 175948
rect 266302 175946 266308 175948
rect 206020 175886 266308 175946
rect 206020 175884 206026 175886
rect 266302 175884 266308 175886
rect 266372 175884 266378 175948
rect 207473 174586 207539 174589
rect 266721 174586 266787 174589
rect 207473 174584 266787 174586
rect 207473 174528 207478 174584
rect 207534 174528 266726 174584
rect 266782 174528 266787 174584
rect 207473 174526 266787 174528
rect 207473 174523 207539 174526
rect 266721 174523 266787 174526
rect 207974 171668 207980 171732
rect 208044 171730 208050 171732
rect 267089 171730 267155 171733
rect 208044 171728 267155 171730
rect 208044 171672 267094 171728
rect 267150 171672 267155 171728
rect 208044 171670 267155 171672
rect 208044 171668 208050 171670
rect 267089 171667 267155 171670
rect 204846 170308 204852 170372
rect 204916 170370 204922 170372
rect 263685 170370 263751 170373
rect 204916 170368 263751 170370
rect 204916 170312 263690 170368
rect 263746 170312 263751 170368
rect 204916 170310 263751 170312
rect 204916 170308 204922 170310
rect 263685 170307 263751 170310
rect 208025 169010 208091 169013
rect 224953 169010 225019 169013
rect 208025 169008 225019 169010
rect 208025 168952 208030 169008
rect 208086 168952 224958 169008
rect 225014 168952 225019 169008
rect 208025 168950 225019 168952
rect 208025 168947 208091 168950
rect 224953 168947 225019 168950
rect 204662 167588 204668 167652
rect 204732 167650 204738 167652
rect 263593 167650 263659 167653
rect 204732 167648 263659 167650
rect 204732 167592 263598 167648
rect 263654 167592 263659 167648
rect 204732 167590 263659 167592
rect 204732 167588 204738 167590
rect 263593 167587 263659 167590
rect 206134 166228 206140 166292
rect 206204 166290 206210 166292
rect 266077 166290 266143 166293
rect 206204 166288 266143 166290
rect 206204 166232 266082 166288
rect 266138 166232 266143 166288
rect 206204 166230 266143 166232
rect 206204 166228 206210 166230
rect 266077 166227 266143 166230
rect 580717 165882 580783 165885
rect 583520 165882 584960 165972
rect 580717 165880 584960 165882
rect 580717 165824 580722 165880
rect 580778 165824 584960 165880
rect 580717 165822 584960 165824
rect 580717 165819 580783 165822
rect 583520 165732 584960 165822
rect 205398 165004 205404 165068
rect 205468 165066 205474 165068
rect 265065 165066 265131 165069
rect 205468 165064 265131 165066
rect 205468 165008 265070 165064
rect 265126 165008 265131 165064
rect 205468 165006 265131 165008
rect 205468 165004 205474 165006
rect 265065 165003 265131 165006
rect 204110 164868 204116 164932
rect 204180 164930 204186 164932
rect 264421 164930 264487 164933
rect 204180 164928 264487 164930
rect 204180 164872 264426 164928
rect 264482 164872 264487 164928
rect 204180 164870 264487 164872
rect 204180 164868 204186 164870
rect 264421 164867 264487 164870
rect 208853 164794 208919 164797
rect 209773 164794 209839 164797
rect 208853 164792 209839 164794
rect 208853 164736 208858 164792
rect 208914 164736 209778 164792
rect 209834 164736 209839 164792
rect 208853 164734 209839 164736
rect 208853 164731 208919 164734
rect 209773 164731 209839 164734
rect 203558 163508 203564 163572
rect 203628 163570 203634 163572
rect 256233 163570 256299 163573
rect 203628 163568 256299 163570
rect 203628 163512 256238 163568
rect 256294 163512 256299 163568
rect 203628 163510 256299 163512
rect 203628 163508 203634 163510
rect 256233 163507 256299 163510
rect 205214 163372 205220 163436
rect 205284 163434 205290 163436
rect 265893 163434 265959 163437
rect 205284 163432 265959 163434
rect 205284 163376 265898 163432
rect 265954 163376 265959 163432
rect 205284 163374 265959 163376
rect 205284 163372 205290 163374
rect 265893 163371 265959 163374
rect -960 162890 480 162980
rect 3693 162890 3759 162893
rect -960 162888 3759 162890
rect -960 162832 3698 162888
rect 3754 162832 3759 162888
rect -960 162830 3759 162832
rect -960 162740 480 162830
rect 3693 162827 3759 162830
rect 203374 162284 203380 162348
rect 203444 162346 203450 162348
rect 247769 162346 247835 162349
rect 203444 162344 247835 162346
rect 203444 162288 247774 162344
rect 247830 162288 247835 162344
rect 203444 162286 247835 162288
rect 203444 162284 203450 162286
rect 247769 162283 247835 162286
rect 203190 162148 203196 162212
rect 203260 162210 203266 162212
rect 258993 162210 259059 162213
rect 203260 162208 259059 162210
rect 203260 162152 258998 162208
rect 259054 162152 259059 162208
rect 203260 162150 259059 162152
rect 203260 162148 203266 162150
rect 258993 162147 259059 162150
rect 206870 162012 206876 162076
rect 206940 162074 206946 162076
rect 267641 162074 267707 162077
rect 206940 162072 267707 162074
rect 206940 162016 267646 162072
rect 267702 162016 267707 162072
rect 206940 162014 267707 162016
rect 206940 162012 206946 162014
rect 267641 162011 267707 162014
rect 202638 161876 202644 161940
rect 202708 161938 202714 161940
rect 263133 161938 263199 161941
rect 202708 161936 263199 161938
rect 202708 161880 263138 161936
rect 263194 161880 263199 161936
rect 202708 161878 263199 161880
rect 202708 161876 202714 161878
rect 263133 161875 263199 161878
rect 265617 161394 265683 161397
rect 207982 161392 265683 161394
rect 207982 161336 265622 161392
rect 265678 161336 265683 161392
rect 207982 161334 265683 161336
rect 203558 161258 203564 161260
rect 195930 161198 203564 161258
rect 169518 160652 169524 160716
rect 169588 160714 169594 160716
rect 186814 160714 186820 160716
rect 169588 160654 186820 160714
rect 169588 160652 169594 160654
rect 186814 160652 186820 160654
rect 186884 160652 186890 160716
rect 159725 160442 159791 160445
rect 163998 160442 164004 160444
rect 159725 160440 164004 160442
rect 159725 160384 159730 160440
rect 159786 160384 164004 160440
rect 159725 160382 164004 160384
rect 159725 160379 159791 160382
rect 163998 160380 164004 160382
rect 164068 160380 164074 160444
rect 155401 160306 155467 160309
rect 162710 160306 162716 160308
rect 155401 160304 162716 160306
rect 155401 160248 155406 160304
rect 155462 160248 162716 160304
rect 155401 160246 162716 160248
rect 155401 160243 155467 160246
rect 162710 160244 162716 160246
rect 162780 160244 162786 160308
rect 171358 160244 171364 160308
rect 171428 160306 171434 160308
rect 172278 160306 172284 160308
rect 171428 160246 172284 160306
rect 171428 160244 171434 160246
rect 172278 160244 172284 160246
rect 172348 160244 172354 160308
rect 151169 160170 151235 160173
rect 151537 160170 151603 160173
rect 175958 160170 175964 160172
rect 151169 160168 164434 160170
rect 151169 160112 151174 160168
rect 151230 160112 151542 160168
rect 151598 160112 164434 160168
rect 151169 160110 164434 160112
rect 151169 160107 151235 160110
rect 151537 160107 151603 160110
rect 163129 159930 163195 159935
rect 162710 159836 162716 159900
rect 162780 159898 162786 159900
rect 162945 159898 163011 159901
rect 162780 159896 163011 159898
rect 162780 159840 162950 159896
rect 163006 159840 163011 159896
rect 163129 159874 163134 159930
rect 163190 159898 163195 159930
rect 163446 159898 163452 159900
rect 163190 159874 163452 159898
rect 163129 159869 163452 159874
rect 162780 159838 163011 159840
rect 163132 159838 163452 159869
rect 162780 159836 162786 159838
rect 162945 159835 163011 159838
rect 163446 159836 163452 159838
rect 163516 159836 163522 159900
rect 163589 159898 163655 159901
rect 164049 159900 164115 159901
rect 163814 159898 163820 159900
rect 163589 159896 163820 159898
rect 163589 159840 163594 159896
rect 163650 159840 163820 159896
rect 163589 159838 163820 159840
rect 163589 159835 163655 159838
rect 163814 159836 163820 159838
rect 163884 159836 163890 159900
rect 163998 159836 164004 159900
rect 164068 159898 164115 159900
rect 164374 159898 164434 160110
rect 168422 160110 169586 160170
rect 165654 159972 165660 160036
rect 165724 160034 165730 160036
rect 168422 160034 168482 160110
rect 169334 160034 169340 160036
rect 165724 159974 166826 160034
rect 165724 159972 165730 159974
rect 166766 159901 166826 159974
rect 166950 159974 168482 160034
rect 168606 159974 169340 160034
rect 164509 159898 164575 159901
rect 164068 159896 164160 159898
rect 164110 159840 164160 159896
rect 164068 159838 164160 159840
rect 164374 159896 164575 159898
rect 164374 159840 164514 159896
rect 164570 159840 164575 159896
rect 164374 159838 164575 159840
rect 164068 159836 164115 159838
rect 164049 159835 164115 159836
rect 164509 159835 164575 159838
rect 164734 159836 164740 159900
rect 164804 159898 164810 159900
rect 165429 159898 165495 159901
rect 164804 159896 165495 159898
rect 164804 159840 165434 159896
rect 165490 159840 165495 159896
rect 164804 159838 165495 159840
rect 164804 159836 164810 159838
rect 165429 159835 165495 159838
rect 165613 159898 165679 159901
rect 166533 159900 166599 159901
rect 165838 159898 165844 159900
rect 165613 159896 165844 159898
rect 165613 159840 165618 159896
rect 165674 159840 165844 159896
rect 165613 159838 165844 159840
rect 165613 159835 165679 159838
rect 165838 159836 165844 159838
rect 165908 159836 165914 159900
rect 166533 159898 166580 159900
rect 166488 159896 166580 159898
rect 166488 159840 166538 159896
rect 166488 159838 166580 159840
rect 166533 159836 166580 159838
rect 166644 159836 166650 159900
rect 166766 159896 166875 159901
rect 166766 159840 166814 159896
rect 166870 159840 166875 159896
rect 166766 159838 166875 159840
rect 166533 159835 166599 159836
rect 166809 159835 166875 159838
rect 166950 159765 167010 159974
rect 167637 159898 167703 159901
rect 167862 159898 167868 159900
rect 167637 159896 167868 159898
rect 167637 159840 167642 159896
rect 167698 159840 167868 159896
rect 167637 159838 167868 159840
rect 167637 159835 167703 159838
rect 167862 159836 167868 159838
rect 167932 159836 167938 159900
rect 168046 159836 168052 159900
rect 168116 159898 168122 159900
rect 168189 159898 168255 159901
rect 168116 159896 168255 159898
rect 168116 159840 168194 159896
rect 168250 159840 168255 159896
rect 168116 159838 168255 159840
rect 168116 159836 168122 159838
rect 168189 159835 168255 159838
rect 168465 159898 168531 159901
rect 168606 159898 168666 159974
rect 169334 159972 169340 159974
rect 169404 159972 169410 160036
rect 169526 160034 169586 160110
rect 171550 160110 175964 160170
rect 169526 159974 169954 160034
rect 168465 159896 168666 159898
rect 168465 159840 168470 159896
rect 168526 159840 168666 159896
rect 168465 159838 168666 159840
rect 169017 159898 169083 159901
rect 169569 159900 169635 159901
rect 169150 159898 169156 159900
rect 169017 159896 169156 159898
rect 169017 159840 169022 159896
rect 169078 159840 169156 159896
rect 169017 159838 169156 159840
rect 168465 159835 168531 159838
rect 169017 159835 169083 159838
rect 169150 159836 169156 159838
rect 169220 159836 169226 159900
rect 169518 159836 169524 159900
rect 169588 159898 169635 159900
rect 169588 159896 169680 159898
rect 169630 159840 169680 159896
rect 169588 159838 169680 159840
rect 169588 159836 169635 159838
rect 169569 159835 169635 159836
rect 162853 159764 162919 159765
rect 162853 159760 162900 159764
rect 162964 159762 162970 159764
rect 162853 159704 162858 159760
rect 162853 159700 162900 159704
rect 162964 159702 163010 159762
rect 162964 159700 162970 159702
rect 163630 159700 163636 159764
rect 163700 159762 163706 159764
rect 163865 159762 163931 159765
rect 163700 159760 163931 159762
rect 163700 159704 163870 159760
rect 163926 159704 163931 159760
rect 163700 159702 163931 159704
rect 163700 159700 163706 159702
rect 162853 159699 162919 159700
rect 163865 159699 163931 159702
rect 164233 159762 164299 159765
rect 164550 159762 164556 159764
rect 164233 159760 164556 159762
rect 164233 159704 164238 159760
rect 164294 159704 164556 159760
rect 164233 159702 164556 159704
rect 164233 159699 164299 159702
rect 164550 159700 164556 159702
rect 164620 159762 164626 159764
rect 165470 159762 165476 159764
rect 164620 159702 165476 159762
rect 164620 159700 164626 159702
rect 165470 159700 165476 159702
rect 165540 159700 165546 159764
rect 166257 159762 166323 159765
rect 166390 159762 166396 159764
rect 166257 159760 166396 159762
rect 166257 159704 166262 159760
rect 166318 159704 166396 159760
rect 166257 159702 166396 159704
rect 166257 159699 166323 159702
rect 166390 159700 166396 159702
rect 166460 159700 166466 159764
rect 166901 159760 167010 159765
rect 166901 159704 166906 159760
rect 166962 159704 167010 159760
rect 166901 159702 167010 159704
rect 167913 159762 167979 159765
rect 168230 159762 168236 159764
rect 167913 159760 168236 159762
rect 167913 159704 167918 159760
rect 167974 159704 168236 159760
rect 167913 159702 168236 159704
rect 166901 159699 166967 159702
rect 167913 159699 167979 159702
rect 168230 159700 168236 159702
rect 168300 159700 168306 159764
rect 168833 159762 168899 159765
rect 168422 159760 168899 159762
rect 168422 159704 168838 159760
rect 168894 159704 168899 159760
rect 168422 159702 168899 159704
rect 155677 159626 155743 159629
rect 167821 159626 167887 159629
rect 168422 159626 168482 159702
rect 168833 159699 168899 159702
rect 168966 159700 168972 159764
rect 169036 159762 169042 159764
rect 169477 159762 169543 159765
rect 169036 159760 169543 159762
rect 169036 159704 169482 159760
rect 169538 159704 169543 159760
rect 169036 159702 169543 159704
rect 169036 159700 169042 159702
rect 169477 159699 169543 159702
rect 155677 159624 167887 159626
rect 155677 159568 155682 159624
rect 155738 159568 167826 159624
rect 167882 159568 167887 159624
rect 155677 159566 167887 159568
rect 155677 159563 155743 159566
rect 167821 159563 167887 159566
rect 168054 159566 168482 159626
rect 152825 159490 152891 159493
rect 168054 159490 168114 159566
rect 168782 159564 168788 159628
rect 168852 159626 168858 159628
rect 169293 159626 169359 159629
rect 168852 159624 169359 159626
rect 168852 159568 169298 159624
rect 169354 159568 169359 159624
rect 168852 159566 169359 159568
rect 168852 159564 168858 159566
rect 169293 159563 169359 159566
rect 152825 159488 168114 159490
rect 152825 159432 152830 159488
rect 152886 159432 168114 159488
rect 152825 159430 168114 159432
rect 169894 159490 169954 159974
rect 171041 159930 171107 159935
rect 170305 159900 170371 159901
rect 170254 159836 170260 159900
rect 170324 159898 170371 159900
rect 170806 159898 170812 159900
rect 170324 159896 170812 159898
rect 170366 159840 170812 159896
rect 170324 159838 170812 159840
rect 170324 159836 170371 159838
rect 170806 159836 170812 159838
rect 170876 159836 170882 159900
rect 171041 159874 171046 159930
rect 171102 159898 171107 159930
rect 171550 159901 171610 160110
rect 175958 160108 175964 160110
rect 176028 160108 176034 160172
rect 195930 160170 195990 161198
rect 203558 161196 203564 161198
rect 203628 161196 203634 161260
rect 207749 161258 207815 161261
rect 207982 161258 208042 161334
rect 265617 161331 265683 161334
rect 207749 161256 208042 161258
rect 207749 161200 207754 161256
rect 207810 161200 208042 161256
rect 207749 161198 208042 161200
rect 210233 161258 210299 161261
rect 264237 161258 264303 161261
rect 210233 161256 264303 161258
rect 210233 161200 210238 161256
rect 210294 161200 264242 161256
rect 264298 161200 264303 161256
rect 210233 161198 264303 161200
rect 207749 161195 207815 161198
rect 210233 161195 210299 161198
rect 264237 161195 264303 161198
rect 198774 161060 198780 161124
rect 198844 161122 198850 161124
rect 259085 161122 259151 161125
rect 198844 161120 259151 161122
rect 198844 161064 259090 161120
rect 259146 161064 259151 161120
rect 198844 161062 259151 161064
rect 198844 161060 198850 161062
rect 259085 161059 259151 161062
rect 198038 160924 198044 160988
rect 198108 160986 198114 160988
rect 258901 160986 258967 160989
rect 198108 160984 258967 160986
rect 198108 160928 258906 160984
rect 258962 160928 258967 160984
rect 198108 160926 258967 160928
rect 198108 160924 198114 160926
rect 258901 160923 258967 160926
rect 269205 160850 269271 160853
rect 202646 160848 269271 160850
rect 202646 160792 269210 160848
rect 269266 160792 269271 160848
rect 202646 160790 269271 160792
rect 195470 160110 195990 160170
rect 171501 159900 171610 159901
rect 171961 159930 172027 159935
rect 171174 159898 171180 159900
rect 171102 159874 171180 159898
rect 171041 159869 171180 159874
rect 171044 159838 171180 159869
rect 171174 159836 171180 159838
rect 171244 159836 171250 159900
rect 171501 159898 171548 159900
rect 171456 159896 171548 159898
rect 171456 159840 171506 159896
rect 171456 159838 171548 159840
rect 171501 159836 171548 159838
rect 171612 159836 171618 159900
rect 171726 159836 171732 159900
rect 171796 159898 171802 159900
rect 171961 159898 171966 159930
rect 171796 159874 171966 159898
rect 172022 159874 172027 159930
rect 174537 159930 174603 159935
rect 171796 159869 172027 159874
rect 172605 159900 172671 159901
rect 172605 159896 172652 159900
rect 172716 159898 172722 159900
rect 172881 159898 172947 159901
rect 173014 159898 173020 159900
rect 171796 159838 172024 159869
rect 172605 159840 172610 159896
rect 171796 159836 171802 159838
rect 172605 159836 172652 159840
rect 172716 159838 172762 159898
rect 172838 159896 173020 159898
rect 172838 159840 172886 159896
rect 172942 159840 173020 159896
rect 172838 159838 173020 159840
rect 172716 159836 172722 159838
rect 170305 159835 170371 159836
rect 171501 159835 171567 159836
rect 172605 159835 172671 159836
rect 172838 159835 172947 159838
rect 173014 159836 173020 159838
rect 173084 159836 173090 159900
rect 173198 159836 173204 159900
rect 173268 159898 173274 159900
rect 173433 159898 173499 159901
rect 173709 159900 173775 159901
rect 174261 159900 174327 159901
rect 173709 159898 173756 159900
rect 173268 159896 173499 159898
rect 173268 159840 173438 159896
rect 173494 159840 173499 159896
rect 173268 159838 173499 159840
rect 173664 159896 173756 159898
rect 173664 159840 173714 159896
rect 173664 159838 173756 159840
rect 173268 159836 173274 159838
rect 173433 159835 173499 159838
rect 173709 159836 173756 159838
rect 173820 159836 173826 159900
rect 174261 159898 174308 159900
rect 174216 159896 174308 159898
rect 174216 159840 174266 159896
rect 174216 159838 174308 159840
rect 174261 159836 174308 159838
rect 174372 159836 174378 159900
rect 174537 159874 174542 159930
rect 174598 159898 174603 159930
rect 174997 159932 175063 159935
rect 174997 159930 175106 159932
rect 174670 159898 174676 159900
rect 174598 159874 174676 159898
rect 174537 159869 174676 159874
rect 174540 159838 174676 159869
rect 174670 159836 174676 159838
rect 174740 159836 174746 159900
rect 174997 159874 175002 159930
rect 175058 159898 175106 159930
rect 195470 159901 195530 160110
rect 198774 160108 198780 160172
rect 198844 160108 198850 160172
rect 202646 160170 202706 160790
rect 269205 160787 269271 160790
rect 277485 160714 277551 160717
rect 201542 160110 202706 160170
rect 202830 160712 277551 160714
rect 202830 160656 277490 160712
rect 277546 160656 277551 160712
rect 202830 160654 277551 160656
rect 198782 159901 198842 160108
rect 175222 159898 175228 159900
rect 175058 159874 175228 159898
rect 174997 159869 175228 159874
rect 175046 159838 175228 159869
rect 175222 159836 175228 159838
rect 175292 159836 175298 159900
rect 175917 159898 175983 159901
rect 176510 159898 176516 159900
rect 175917 159896 176516 159898
rect 175917 159840 175922 159896
rect 175978 159840 176516 159896
rect 175917 159838 176516 159840
rect 173709 159835 173775 159836
rect 174261 159835 174327 159836
rect 175917 159835 175983 159838
rect 176510 159836 176516 159838
rect 176580 159836 176586 159900
rect 178125 159898 178191 159901
rect 178902 159898 178908 159900
rect 178125 159896 178908 159898
rect 178125 159840 178130 159896
rect 178186 159840 178908 159896
rect 178125 159838 178908 159840
rect 178125 159835 178191 159838
rect 178902 159836 178908 159838
rect 178972 159836 178978 159900
rect 180057 159898 180123 159901
rect 180609 159900 180675 159901
rect 180374 159898 180380 159900
rect 180057 159896 180380 159898
rect 180057 159840 180062 159896
rect 180118 159840 180380 159896
rect 180057 159838 180380 159840
rect 180057 159835 180123 159838
rect 180374 159836 180380 159838
rect 180444 159836 180450 159900
rect 180558 159898 180564 159900
rect 180518 159838 180564 159898
rect 180628 159896 180675 159900
rect 180670 159840 180675 159896
rect 180558 159836 180564 159838
rect 180628 159836 180675 159840
rect 180609 159835 180675 159836
rect 181161 159898 181227 159901
rect 182541 159900 182607 159901
rect 181478 159898 181484 159900
rect 181161 159896 181484 159898
rect 181161 159840 181166 159896
rect 181222 159840 181484 159896
rect 181161 159838 181484 159840
rect 181161 159835 181227 159838
rect 181478 159836 181484 159838
rect 181548 159836 181554 159900
rect 182541 159898 182588 159900
rect 182496 159896 182588 159898
rect 182496 159840 182546 159896
rect 182496 159838 182588 159840
rect 182541 159836 182588 159838
rect 182652 159836 182658 159900
rect 183134 159836 183140 159900
rect 183204 159898 183210 159900
rect 183369 159898 183435 159901
rect 183204 159896 183435 159898
rect 183204 159840 183374 159896
rect 183430 159840 183435 159896
rect 183204 159838 183435 159840
rect 183204 159836 183210 159838
rect 182541 159835 182607 159836
rect 183369 159835 183435 159838
rect 183921 159898 183987 159901
rect 184054 159898 184060 159900
rect 183921 159896 184060 159898
rect 183921 159840 183926 159896
rect 183982 159840 184060 159896
rect 183921 159838 184060 159840
rect 183921 159835 183987 159838
rect 184054 159836 184060 159838
rect 184124 159836 184130 159900
rect 184473 159898 184539 159901
rect 184606 159898 184612 159900
rect 184473 159896 184612 159898
rect 184473 159840 184478 159896
rect 184534 159840 184612 159896
rect 184473 159838 184612 159840
rect 184473 159835 184539 159838
rect 184606 159836 184612 159838
rect 184676 159836 184682 159900
rect 185158 159836 185164 159900
rect 185228 159898 185234 159900
rect 185301 159898 185367 159901
rect 185228 159896 185367 159898
rect 185228 159840 185306 159896
rect 185362 159840 185367 159896
rect 185228 159838 185367 159840
rect 185228 159836 185234 159838
rect 185301 159835 185367 159838
rect 188337 159898 188403 159901
rect 188470 159898 188476 159900
rect 188337 159896 188476 159898
rect 188337 159840 188342 159896
rect 188398 159840 188476 159896
rect 188337 159838 188476 159840
rect 188337 159835 188403 159838
rect 188470 159836 188476 159838
rect 188540 159898 188546 159900
rect 188838 159898 188844 159900
rect 188540 159838 188844 159898
rect 188540 159836 188546 159838
rect 188838 159836 188844 159838
rect 188908 159836 188914 159900
rect 189717 159898 189783 159901
rect 190310 159898 190316 159900
rect 189717 159896 190316 159898
rect 189717 159840 189722 159896
rect 189778 159840 190316 159896
rect 189717 159838 190316 159840
rect 189717 159835 189783 159838
rect 190310 159836 190316 159838
rect 190380 159836 190386 159900
rect 191097 159896 191163 159901
rect 191097 159840 191102 159896
rect 191158 159840 191163 159896
rect 191097 159835 191163 159840
rect 192201 159898 192267 159901
rect 193581 159900 193647 159901
rect 193070 159898 193076 159900
rect 192201 159896 193076 159898
rect 192201 159840 192206 159896
rect 192262 159840 193076 159896
rect 192201 159838 193076 159840
rect 192201 159835 192267 159838
rect 193070 159836 193076 159838
rect 193140 159836 193146 159900
rect 193581 159898 193628 159900
rect 193536 159896 193628 159898
rect 193536 159840 193586 159896
rect 193536 159838 193628 159840
rect 193581 159836 193628 159838
rect 193692 159836 193698 159900
rect 193857 159898 193923 159901
rect 195237 159900 195303 159901
rect 194358 159898 194364 159900
rect 193857 159896 194364 159898
rect 193857 159840 193862 159896
rect 193918 159840 194364 159896
rect 193857 159838 194364 159840
rect 193581 159835 193647 159836
rect 193857 159835 193923 159838
rect 194358 159836 194364 159838
rect 194428 159836 194434 159900
rect 195237 159898 195284 159900
rect 195192 159896 195284 159898
rect 195192 159840 195242 159896
rect 195192 159838 195284 159840
rect 195237 159836 195284 159838
rect 195348 159836 195354 159900
rect 195470 159896 195579 159901
rect 195789 159900 195855 159901
rect 195789 159898 195836 159900
rect 195470 159840 195518 159896
rect 195574 159840 195579 159896
rect 195470 159838 195579 159840
rect 195744 159896 195836 159898
rect 195744 159840 195794 159896
rect 195744 159838 195836 159840
rect 195237 159835 195303 159836
rect 195513 159835 195579 159838
rect 195789 159836 195836 159838
rect 195900 159836 195906 159900
rect 196617 159898 196683 159901
rect 197118 159898 197124 159900
rect 196617 159896 197124 159898
rect 196617 159840 196622 159896
rect 196678 159840 197124 159896
rect 196617 159838 197124 159840
rect 195789 159835 195855 159836
rect 196617 159835 196683 159838
rect 197118 159836 197124 159838
rect 197188 159836 197194 159900
rect 197854 159836 197860 159900
rect 197924 159898 197930 159900
rect 197997 159898 198063 159901
rect 197924 159896 198063 159898
rect 197924 159840 198002 159896
rect 198058 159840 198063 159896
rect 197924 159838 198063 159840
rect 197924 159836 197930 159838
rect 197997 159835 198063 159838
rect 198222 159836 198228 159900
rect 198292 159898 198298 159900
rect 198549 159898 198615 159901
rect 198292 159896 198615 159898
rect 198292 159840 198554 159896
rect 198610 159840 198615 159896
rect 198292 159838 198615 159840
rect 198782 159896 198891 159901
rect 199101 159900 199167 159901
rect 199101 159898 199148 159900
rect 198782 159840 198830 159896
rect 198886 159840 198891 159896
rect 198782 159838 198891 159840
rect 199056 159896 199148 159898
rect 199056 159840 199106 159896
rect 199056 159838 199148 159840
rect 198292 159836 198298 159838
rect 198549 159835 198615 159838
rect 198825 159835 198891 159838
rect 199101 159836 199148 159838
rect 199212 159836 199218 159900
rect 199377 159898 199443 159901
rect 199878 159898 199884 159900
rect 199377 159896 199884 159898
rect 199377 159840 199382 159896
rect 199438 159840 199884 159896
rect 199377 159838 199884 159840
rect 199101 159835 199167 159836
rect 199377 159835 199443 159838
rect 199878 159836 199884 159838
rect 199948 159836 199954 159900
rect 200205 159898 200271 159901
rect 200982 159898 200988 159900
rect 200205 159896 200988 159898
rect 200205 159840 200210 159896
rect 200266 159840 200988 159896
rect 200205 159838 200988 159840
rect 200205 159835 200271 159838
rect 200982 159836 200988 159838
rect 201052 159898 201058 159900
rect 201350 159898 201356 159900
rect 201052 159838 201356 159898
rect 201052 159836 201058 159838
rect 201350 159836 201356 159838
rect 201420 159836 201426 159900
rect 170673 159764 170739 159765
rect 170070 159700 170076 159764
rect 170140 159762 170146 159764
rect 170622 159762 170628 159764
rect 170140 159702 170628 159762
rect 170692 159760 170739 159764
rect 170734 159704 170739 159760
rect 170140 159700 170146 159702
rect 170622 159700 170628 159702
rect 170692 159700 170739 159704
rect 170673 159699 170739 159700
rect 171133 159762 171199 159765
rect 171358 159762 171364 159764
rect 171133 159760 171364 159762
rect 171133 159704 171138 159760
rect 171194 159704 171364 159760
rect 171133 159702 171364 159704
rect 171133 159699 171199 159702
rect 171358 159700 171364 159702
rect 171428 159700 171434 159764
rect 171910 159700 171916 159764
rect 171980 159762 171986 159764
rect 172053 159762 172119 159765
rect 171980 159760 172119 159762
rect 171980 159704 172058 159760
rect 172114 159704 172119 159760
rect 171980 159702 172119 159704
rect 171980 159700 171986 159702
rect 172053 159699 172119 159702
rect 172697 159762 172763 159765
rect 172838 159762 172898 159835
rect 172697 159760 172898 159762
rect 172697 159704 172702 159760
rect 172758 159704 172898 159760
rect 172697 159702 172898 159704
rect 173157 159762 173223 159765
rect 173566 159762 173572 159764
rect 173157 159760 173572 159762
rect 173157 159704 173162 159760
rect 173218 159704 173572 159760
rect 173157 159702 173572 159704
rect 172697 159699 172763 159702
rect 173157 159699 173223 159702
rect 173566 159700 173572 159702
rect 173636 159700 173642 159764
rect 174486 159700 174492 159764
rect 174556 159762 174562 159764
rect 174813 159762 174879 159765
rect 175089 159762 175155 159765
rect 176377 159764 176443 159765
rect 174556 159760 175155 159762
rect 174556 159704 174818 159760
rect 174874 159704 175094 159760
rect 175150 159704 175155 159760
rect 174556 159702 175155 159704
rect 174556 159700 174562 159702
rect 174813 159699 174879 159702
rect 175089 159699 175155 159702
rect 176326 159700 176332 159764
rect 176396 159762 176443 159764
rect 176396 159760 176488 159762
rect 176438 159704 176488 159760
rect 176396 159702 176488 159704
rect 176396 159700 176443 159702
rect 178534 159700 178540 159764
rect 178604 159762 178610 159764
rect 178677 159762 178743 159765
rect 178604 159760 178743 159762
rect 178604 159704 178682 159760
rect 178738 159704 178743 159760
rect 178604 159702 178743 159704
rect 178604 159700 178610 159702
rect 176377 159699 176443 159700
rect 178677 159699 178743 159702
rect 178953 159762 179019 159765
rect 180926 159762 180932 159764
rect 178953 159760 180932 159762
rect 178953 159704 178958 159760
rect 179014 159704 180932 159760
rect 178953 159702 180932 159704
rect 178953 159699 179019 159702
rect 180926 159700 180932 159702
rect 180996 159700 181002 159764
rect 182541 159762 182607 159765
rect 182766 159762 182772 159764
rect 182541 159760 182772 159762
rect 182541 159704 182546 159760
rect 182602 159704 182772 159760
rect 182541 159702 182772 159704
rect 182541 159699 182607 159702
rect 182766 159700 182772 159702
rect 182836 159700 182842 159764
rect 184197 159762 184263 159765
rect 184422 159762 184428 159764
rect 184197 159760 184428 159762
rect 184197 159704 184202 159760
rect 184258 159704 184428 159760
rect 184197 159702 184428 159704
rect 184197 159699 184263 159702
rect 184422 159700 184428 159702
rect 184492 159700 184498 159764
rect 191100 159762 191160 159835
rect 191598 159762 191604 159764
rect 191100 159702 191604 159762
rect 191598 159700 191604 159702
rect 191668 159762 191674 159764
rect 191741 159762 191807 159765
rect 191668 159760 191807 159762
rect 191668 159704 191746 159760
rect 191802 159704 191807 159760
rect 191668 159702 191807 159704
rect 191668 159700 191674 159702
rect 191741 159699 191807 159702
rect 194961 159762 195027 159765
rect 196341 159764 196407 159765
rect 195646 159762 195652 159764
rect 194961 159760 195652 159762
rect 194961 159704 194966 159760
rect 195022 159704 195652 159760
rect 194961 159702 195652 159704
rect 194961 159699 195027 159702
rect 195646 159700 195652 159702
rect 195716 159700 195722 159764
rect 196341 159762 196388 159764
rect 196260 159760 196388 159762
rect 196452 159762 196458 159764
rect 196934 159762 196940 159764
rect 196260 159704 196346 159760
rect 196260 159702 196388 159704
rect 196341 159700 196388 159702
rect 196452 159702 196940 159762
rect 196452 159700 196458 159702
rect 196934 159700 196940 159702
rect 197004 159700 197010 159764
rect 197721 159762 197787 159765
rect 198406 159762 198412 159764
rect 197721 159760 198412 159762
rect 197721 159704 197726 159760
rect 197782 159704 198412 159760
rect 197721 159702 198412 159704
rect 196341 159699 196407 159700
rect 197721 159699 197787 159702
rect 198406 159700 198412 159702
rect 198476 159700 198482 159764
rect 199326 159700 199332 159764
rect 199396 159762 199402 159764
rect 199653 159762 199719 159765
rect 199396 159760 199719 159762
rect 199396 159704 199658 159760
rect 199714 159704 199719 159760
rect 199396 159702 199719 159704
rect 199396 159700 199402 159702
rect 199653 159699 199719 159702
rect 201217 159762 201283 159765
rect 201542 159762 201602 160110
rect 202830 159901 202890 160654
rect 277485 160651 277551 160654
rect 230105 160578 230171 160581
rect 215250 160576 230171 160578
rect 215250 160520 230110 160576
rect 230166 160520 230171 160576
rect 215250 160518 230171 160520
rect 208945 160442 209011 160445
rect 205360 160440 209011 160442
rect 205360 160384 208950 160440
rect 209006 160384 209011 160440
rect 205360 160382 209011 160384
rect 203558 160306 203564 160308
rect 203244 160246 203564 160306
rect 203244 159935 203304 160246
rect 203558 160244 203564 160246
rect 203628 160306 203634 160308
rect 205360 160306 205420 160382
rect 208945 160379 209011 160382
rect 210233 160306 210299 160309
rect 203628 160246 205420 160306
rect 206326 160304 210299 160306
rect 206326 160248 210238 160304
rect 210294 160248 210299 160304
rect 206326 160246 210299 160248
rect 203628 160244 203634 160246
rect 206326 160170 206386 160246
rect 210233 160243 210299 160246
rect 215250 160170 215310 160518
rect 230105 160515 230171 160518
rect 204302 160110 206386 160170
rect 207062 160110 215310 160170
rect 203241 159930 203307 159935
rect 202830 159896 202939 159901
rect 202830 159840 202878 159896
rect 202934 159840 202939 159896
rect 203241 159874 203246 159930
rect 203302 159874 203307 159930
rect 204302 159901 204362 160110
rect 204069 159900 204135 159901
rect 204069 159898 204116 159900
rect 203241 159869 203307 159874
rect 204024 159896 204116 159898
rect 202830 159838 202939 159840
rect 204024 159840 204074 159896
rect 204024 159838 204116 159840
rect 202873 159835 202939 159838
rect 204069 159836 204116 159838
rect 204180 159836 204186 159900
rect 204253 159896 204362 159901
rect 204253 159840 204258 159896
rect 204314 159840 204362 159896
rect 204253 159838 204362 159840
rect 204069 159835 204135 159836
rect 204253 159835 204319 159838
rect 204662 159836 204668 159900
rect 204732 159898 204738 159900
rect 204897 159898 204963 159901
rect 205173 159900 205239 159901
rect 205449 159900 205515 159901
rect 205173 159898 205220 159900
rect 204732 159896 204963 159898
rect 204732 159840 204902 159896
rect 204958 159840 204963 159896
rect 204732 159838 204963 159840
rect 205128 159896 205220 159898
rect 205128 159840 205178 159896
rect 205128 159838 205220 159840
rect 204732 159836 204738 159838
rect 204897 159835 204963 159838
rect 205173 159836 205220 159838
rect 205284 159836 205290 159900
rect 205398 159836 205404 159900
rect 205468 159898 205515 159900
rect 205468 159896 205560 159898
rect 205510 159840 205560 159896
rect 205468 159838 205560 159840
rect 205468 159836 205515 159838
rect 205766 159836 205772 159900
rect 205836 159898 205842 159900
rect 206277 159898 206343 159901
rect 205836 159896 206343 159898
rect 205836 159840 206282 159896
rect 206338 159840 206343 159896
rect 205836 159838 206343 159840
rect 205836 159836 205842 159838
rect 205173 159835 205239 159836
rect 205449 159835 205515 159836
rect 206277 159835 206343 159838
rect 207062 159765 207122 160110
rect 207289 159898 207355 159901
rect 207974 159898 207980 159900
rect 207289 159896 207980 159898
rect 207289 159840 207294 159896
rect 207350 159840 207980 159896
rect 207289 159838 207980 159840
rect 207289 159835 207355 159838
rect 207974 159836 207980 159838
rect 208044 159836 208050 159900
rect 202413 159764 202479 159765
rect 202689 159764 202755 159765
rect 202413 159762 202460 159764
rect 201217 159760 201602 159762
rect 201217 159704 201222 159760
rect 201278 159704 201602 159760
rect 201217 159702 201602 159704
rect 202368 159760 202460 159762
rect 202368 159704 202418 159760
rect 202368 159702 202460 159704
rect 201217 159699 201283 159702
rect 202413 159700 202460 159702
rect 202524 159700 202530 159764
rect 202638 159700 202644 159764
rect 202708 159762 202755 159764
rect 204621 159762 204687 159765
rect 204846 159762 204852 159764
rect 202708 159760 202800 159762
rect 202750 159704 202800 159760
rect 202708 159702 202800 159704
rect 204621 159760 204852 159762
rect 204621 159704 204626 159760
rect 204682 159704 204852 159760
rect 204621 159702 204852 159704
rect 202708 159700 202755 159702
rect 202413 159699 202479 159700
rect 202689 159699 202755 159700
rect 204621 159699 204687 159702
rect 204846 159700 204852 159702
rect 204916 159700 204922 159764
rect 205950 159700 205956 159764
rect 206020 159762 206026 159764
rect 206829 159762 206895 159765
rect 206020 159760 206895 159762
rect 206020 159704 206834 159760
rect 206890 159704 206895 159760
rect 206020 159702 206895 159704
rect 206020 159700 206026 159702
rect 206829 159699 206895 159702
rect 207013 159760 207122 159765
rect 207013 159704 207018 159760
rect 207074 159704 207122 159760
rect 207013 159702 207122 159704
rect 207381 159762 207447 159765
rect 207790 159762 207796 159764
rect 207381 159760 207796 159762
rect 207381 159704 207386 159760
rect 207442 159704 207796 159760
rect 207381 159702 207796 159704
rect 207013 159699 207079 159702
rect 207381 159699 207447 159702
rect 207790 159700 207796 159702
rect 207860 159700 207866 159764
rect 170121 159626 170187 159629
rect 170438 159626 170444 159628
rect 170121 159624 170444 159626
rect 170121 159568 170126 159624
rect 170182 159568 170444 159624
rect 170121 159566 170444 159568
rect 170121 159563 170187 159566
rect 170438 159564 170444 159566
rect 170508 159564 170514 159628
rect 171685 159626 171751 159629
rect 172094 159626 172100 159628
rect 171685 159624 172100 159626
rect 171685 159568 171690 159624
rect 171746 159568 172100 159624
rect 171685 159566 172100 159568
rect 171685 159563 171751 159566
rect 172094 159564 172100 159566
rect 172164 159564 172170 159628
rect 173985 159626 174051 159629
rect 174721 159626 174787 159629
rect 175038 159626 175044 159628
rect 173985 159624 175044 159626
rect 173985 159568 173990 159624
rect 174046 159568 174726 159624
rect 174782 159568 175044 159624
rect 173985 159566 175044 159568
rect 173985 159563 174051 159566
rect 174721 159563 174787 159566
rect 175038 159564 175044 159566
rect 175108 159564 175114 159628
rect 180885 159626 180951 159629
rect 181110 159626 181116 159628
rect 180885 159624 181116 159626
rect 180885 159568 180890 159624
rect 180946 159568 181116 159624
rect 180885 159566 181116 159568
rect 180885 159563 180951 159566
rect 181110 159564 181116 159566
rect 181180 159564 181186 159628
rect 198038 159564 198044 159628
rect 198108 159626 198114 159628
rect 198181 159626 198247 159629
rect 198108 159624 198247 159626
rect 198108 159568 198186 159624
rect 198242 159568 198247 159624
rect 198108 159566 198247 159568
rect 198108 159564 198114 159566
rect 198181 159563 198247 159566
rect 198457 159626 198523 159629
rect 249149 159626 249215 159629
rect 198457 159624 249215 159626
rect 198457 159568 198462 159624
rect 198518 159568 249154 159624
rect 249210 159568 249215 159624
rect 198457 159566 249215 159568
rect 198457 159563 198523 159566
rect 249149 159563 249215 159566
rect 175774 159490 175780 159492
rect 169894 159430 175780 159490
rect 152825 159427 152891 159430
rect 175774 159428 175780 159430
rect 175844 159428 175850 159492
rect 177246 159490 177252 159492
rect 176610 159430 177252 159490
rect 156873 159354 156939 159357
rect 165613 159354 165679 159357
rect 156873 159352 165679 159354
rect 156873 159296 156878 159352
rect 156934 159296 165618 159352
rect 165674 159296 165679 159352
rect 156873 159294 165679 159296
rect 156873 159291 156939 159294
rect 165613 159291 165679 159294
rect 170949 159356 171015 159357
rect 170949 159352 170996 159356
rect 171060 159354 171066 159356
rect 171593 159354 171659 159357
rect 176610 159354 176670 159430
rect 177246 159428 177252 159430
rect 177316 159428 177322 159492
rect 187417 159490 187483 159493
rect 227662 159490 227668 159492
rect 187417 159488 227668 159490
rect 187417 159432 187422 159488
rect 187478 159432 227668 159488
rect 187417 159430 227668 159432
rect 187417 159427 187483 159430
rect 227662 159428 227668 159430
rect 227732 159428 227738 159492
rect 170949 159296 170954 159352
rect 170949 159292 170996 159296
rect 171060 159294 171106 159354
rect 171593 159352 176670 159354
rect 171593 159296 171598 159352
rect 171654 159296 176670 159352
rect 171593 159294 176670 159296
rect 200941 159354 201007 159357
rect 260097 159354 260163 159357
rect 200941 159352 260163 159354
rect 200941 159296 200946 159352
rect 201002 159296 260102 159352
rect 260158 159296 260163 159352
rect 200941 159294 260163 159296
rect 171060 159292 171066 159294
rect 170949 159291 171015 159292
rect 171593 159291 171659 159294
rect 200941 159291 201007 159294
rect 260097 159291 260163 159294
rect 159449 159218 159515 159221
rect 167821 159218 167887 159221
rect 171501 159218 171567 159221
rect 159449 159216 167746 159218
rect 159449 159160 159454 159216
rect 159510 159160 167746 159216
rect 159449 159158 167746 159160
rect 159449 159155 159515 159158
rect 149145 159082 149211 159085
rect 150249 159082 150315 159085
rect 165061 159082 165127 159085
rect 149145 159080 165127 159082
rect 149145 159024 149150 159080
rect 149206 159024 150254 159080
rect 150310 159024 165066 159080
rect 165122 159024 165127 159080
rect 149145 159022 165127 159024
rect 149145 159019 149211 159022
rect 150249 159019 150315 159022
rect 165061 159019 165127 159022
rect 165889 159082 165955 159085
rect 166901 159082 166967 159085
rect 165889 159080 166967 159082
rect 165889 159024 165894 159080
rect 165950 159024 166906 159080
rect 166962 159024 166967 159080
rect 165889 159022 166967 159024
rect 167686 159082 167746 159158
rect 167821 159216 171567 159218
rect 167821 159160 167826 159216
rect 167882 159160 171506 159216
rect 171562 159160 171567 159216
rect 167821 159158 171567 159160
rect 167821 159155 167887 159158
rect 171501 159155 171567 159158
rect 172462 159156 172468 159220
rect 172532 159218 172538 159220
rect 172881 159218 172947 159221
rect 172532 159216 172947 159218
rect 172532 159160 172886 159216
rect 172942 159160 172947 159216
rect 172532 159158 172947 159160
rect 172532 159156 172538 159158
rect 172881 159155 172947 159158
rect 173985 159218 174051 159221
rect 176101 159218 176167 159221
rect 173985 159216 176167 159218
rect 173985 159160 173990 159216
rect 174046 159160 176106 159216
rect 176162 159160 176167 159216
rect 173985 159158 176167 159160
rect 173985 159155 174051 159158
rect 176101 159155 176167 159158
rect 197077 159218 197143 159221
rect 203374 159218 203380 159220
rect 197077 159216 203380 159218
rect 197077 159160 197082 159216
rect 197138 159160 203380 159216
rect 197077 159158 203380 159160
rect 197077 159155 197143 159158
rect 203374 159156 203380 159158
rect 203444 159156 203450 159220
rect 206001 159218 206067 159221
rect 206134 159218 206140 159220
rect 206001 159216 206140 159218
rect 206001 159160 206006 159216
rect 206062 159160 206140 159216
rect 206001 159158 206140 159160
rect 206001 159155 206067 159158
rect 206134 159156 206140 159158
rect 206204 159156 206210 159220
rect 206737 159218 206803 159221
rect 266997 159218 267063 159221
rect 206737 159216 267063 159218
rect 206737 159160 206742 159216
rect 206798 159160 267002 159216
rect 267058 159160 267063 159216
rect 206737 159158 267063 159160
rect 206737 159155 206803 159158
rect 266997 159155 267063 159158
rect 174169 159082 174235 159085
rect 167686 159080 174235 159082
rect 167686 159024 174174 159080
rect 174230 159024 174235 159080
rect 167686 159022 174235 159024
rect 165889 159019 165955 159022
rect 166901 159019 166967 159022
rect 174169 159019 174235 159022
rect 192518 159020 192524 159084
rect 192588 159082 192594 159084
rect 193029 159082 193095 159085
rect 192588 159080 193095 159082
rect 192588 159024 193034 159080
rect 193090 159024 193095 159080
rect 192588 159022 193095 159024
rect 192588 159020 192594 159022
rect 193029 159019 193095 159022
rect 202321 159082 202387 159085
rect 263041 159082 263107 159085
rect 202321 159080 263107 159082
rect 202321 159024 202326 159080
rect 202382 159024 263046 159080
rect 263102 159024 263107 159080
rect 202321 159022 263107 159024
rect 202321 159019 202387 159022
rect 263041 159019 263107 159022
rect 154021 158946 154087 158949
rect 166809 158946 166875 158949
rect 154021 158944 166875 158946
rect 154021 158888 154026 158944
rect 154082 158888 166814 158944
rect 166870 158888 166875 158944
rect 154021 158886 166875 158888
rect 154021 158883 154087 158886
rect 166809 158883 166875 158886
rect 169753 158946 169819 158949
rect 171501 158948 171567 158949
rect 170070 158946 170076 158948
rect 169753 158944 170076 158946
rect 169753 158888 169758 158944
rect 169814 158888 170076 158944
rect 169753 158886 170076 158888
rect 169753 158883 169819 158886
rect 170070 158884 170076 158886
rect 170140 158884 170146 158948
rect 171501 158944 171548 158948
rect 171612 158946 171618 158948
rect 198917 158946 198983 158949
rect 199142 158946 199148 158948
rect 171501 158888 171506 158944
rect 171501 158884 171548 158888
rect 171612 158886 171658 158946
rect 198917 158944 199148 158946
rect 198917 158888 198922 158944
rect 198978 158888 199148 158944
rect 198917 158886 199148 158888
rect 171612 158884 171618 158886
rect 171501 158883 171567 158884
rect 198917 158883 198983 158886
rect 199142 158884 199148 158886
rect 199212 158946 199218 158948
rect 200941 158946 201007 158949
rect 199212 158944 201007 158946
rect 199212 158888 200946 158944
rect 201002 158888 201007 158944
rect 199212 158886 201007 158888
rect 199212 158884 199218 158886
rect 200941 158883 201007 158886
rect 203977 158946 204043 158949
rect 268009 158946 268075 158949
rect 203977 158944 268075 158946
rect 203977 158888 203982 158944
rect 204038 158888 268014 158944
rect 268070 158888 268075 158944
rect 203977 158886 268075 158888
rect 203977 158883 204043 158886
rect 268009 158883 268075 158886
rect 155309 158810 155375 158813
rect 155677 158810 155743 158813
rect 155309 158808 155743 158810
rect 155309 158752 155314 158808
rect 155370 158752 155682 158808
rect 155738 158752 155743 158808
rect 155309 158750 155743 158752
rect 155309 158747 155375 158750
rect 155677 158747 155743 158750
rect 155861 158810 155927 158813
rect 168005 158810 168071 158813
rect 188286 158810 188292 158812
rect 155861 158808 168071 158810
rect 155861 158752 155866 158808
rect 155922 158752 168010 158808
rect 168066 158752 168071 158808
rect 155861 158750 168071 158752
rect 155861 158747 155927 158750
rect 168005 158747 168071 158750
rect 168238 158750 188292 158810
rect 158713 158674 158779 158677
rect 159909 158674 159975 158677
rect 158713 158672 159975 158674
rect 158713 158616 158718 158672
rect 158774 158616 159914 158672
rect 159970 158616 159975 158672
rect 158713 158614 159975 158616
rect 158713 158611 158779 158614
rect 159909 158611 159975 158614
rect 160093 158674 160159 158677
rect 161105 158674 161171 158677
rect 160093 158672 161171 158674
rect 160093 158616 160098 158672
rect 160154 158616 161110 158672
rect 161166 158616 161171 158672
rect 160093 158614 161171 158616
rect 160093 158611 160159 158614
rect 161105 158611 161171 158614
rect 163313 158674 163379 158677
rect 164233 158676 164299 158677
rect 164785 158676 164851 158677
rect 163446 158674 163452 158676
rect 163313 158672 163452 158674
rect 163313 158616 163318 158672
rect 163374 158616 163452 158672
rect 163313 158614 163452 158616
rect 163313 158611 163379 158614
rect 163446 158612 163452 158614
rect 163516 158612 163522 158676
rect 164182 158674 164188 158676
rect 164142 158614 164188 158674
rect 164252 158672 164299 158676
rect 164294 158616 164299 158672
rect 164182 158612 164188 158614
rect 164252 158612 164299 158616
rect 164734 158612 164740 158676
rect 164804 158674 164851 158676
rect 165153 158674 165219 158677
rect 165705 158676 165771 158677
rect 166073 158676 166139 158677
rect 165286 158674 165292 158676
rect 164804 158672 164896 158674
rect 164846 158616 164896 158672
rect 164804 158614 164896 158616
rect 165153 158672 165292 158674
rect 165153 158616 165158 158672
rect 165214 158616 165292 158672
rect 165153 158614 165292 158616
rect 164804 158612 164851 158614
rect 164233 158611 164299 158612
rect 164785 158611 164851 158612
rect 165153 158611 165219 158614
rect 165286 158612 165292 158614
rect 165356 158612 165362 158676
rect 165654 158612 165660 158676
rect 165724 158674 165771 158676
rect 166022 158674 166028 158676
rect 165724 158672 165816 158674
rect 165766 158616 165816 158672
rect 165724 158614 165816 158616
rect 165946 158614 166028 158674
rect 166092 158674 166139 158676
rect 167678 158674 167684 158676
rect 166092 158672 167684 158674
rect 166134 158616 167684 158672
rect 165724 158612 165771 158614
rect 166022 158612 166028 158614
rect 166092 158614 167684 158616
rect 166092 158612 166139 158614
rect 167678 158612 167684 158614
rect 167748 158612 167754 158676
rect 167821 158674 167887 158677
rect 168238 158674 168298 158750
rect 188286 158748 188292 158750
rect 188356 158748 188362 158812
rect 192385 158810 192451 158813
rect 192342 158808 192451 158810
rect 192342 158752 192390 158808
rect 192446 158752 192451 158808
rect 192342 158747 192451 158752
rect 203977 158810 204043 158813
rect 205909 158810 205975 158813
rect 270861 158810 270927 158813
rect 203977 158808 204178 158810
rect 203977 158752 203982 158808
rect 204038 158752 204178 158808
rect 203977 158750 204178 158752
rect 203977 158747 204043 158750
rect 167821 158672 168298 158674
rect 167821 158616 167826 158672
rect 167882 158616 168298 158672
rect 167821 158614 168298 158616
rect 165705 158611 165771 158612
rect 166073 158611 166139 158612
rect 167821 158611 167887 158614
rect 168414 158612 168420 158676
rect 168484 158674 168490 158676
rect 168649 158674 168715 158677
rect 168484 158672 168715 158674
rect 168484 158616 168654 158672
rect 168710 158616 168715 158672
rect 168484 158614 168715 158616
rect 168484 158612 168490 158614
rect 168649 158611 168715 158614
rect 168966 158612 168972 158676
rect 169036 158674 169042 158676
rect 169385 158674 169451 158677
rect 169036 158672 169451 158674
rect 169036 158616 169390 158672
rect 169446 158616 169451 158672
rect 169036 158614 169451 158616
rect 169036 158612 169042 158614
rect 169385 158611 169451 158614
rect 169845 158674 169911 158677
rect 170254 158674 170260 158676
rect 169845 158672 170260 158674
rect 169845 158616 169850 158672
rect 169906 158616 170260 158672
rect 169845 158614 170260 158616
rect 169845 158611 169911 158614
rect 170254 158612 170260 158614
rect 170324 158612 170330 158676
rect 171726 158612 171732 158676
rect 171796 158674 171802 158676
rect 171869 158674 171935 158677
rect 172329 158676 172395 158677
rect 172278 158674 172284 158676
rect 171796 158672 171935 158674
rect 171796 158616 171874 158672
rect 171930 158616 171935 158672
rect 171796 158614 171935 158616
rect 172238 158614 172284 158674
rect 172348 158672 172395 158676
rect 172390 158616 172395 158672
rect 171796 158612 171802 158614
rect 171869 158611 171935 158614
rect 172278 158612 172284 158614
rect 172348 158612 172395 158616
rect 172329 158611 172395 158612
rect 173065 158674 173131 158677
rect 173198 158674 173204 158676
rect 173065 158672 173204 158674
rect 173065 158616 173070 158672
rect 173126 158616 173204 158672
rect 173065 158614 173204 158616
rect 173065 158611 173131 158614
rect 173198 158612 173204 158614
rect 173268 158612 173274 158676
rect 173893 158674 173959 158677
rect 175038 158674 175044 158676
rect 173893 158672 175044 158674
rect 173893 158616 173898 158672
rect 173954 158616 175044 158672
rect 173893 158614 175044 158616
rect 173893 158611 173959 158614
rect 175038 158612 175044 158614
rect 175108 158612 175114 158676
rect 175406 158612 175412 158676
rect 175476 158674 175482 158676
rect 175641 158674 175707 158677
rect 175476 158672 175707 158674
rect 175476 158616 175646 158672
rect 175702 158616 175707 158672
rect 175476 158614 175707 158616
rect 175476 158612 175482 158614
rect 175641 158611 175707 158614
rect 176009 158674 176075 158677
rect 176326 158674 176332 158676
rect 176009 158672 176332 158674
rect 176009 158616 176014 158672
rect 176070 158616 176332 158672
rect 176009 158614 176332 158616
rect 176009 158611 176075 158614
rect 176326 158612 176332 158614
rect 176396 158612 176402 158676
rect 178718 158612 178724 158676
rect 178788 158674 178794 158676
rect 179229 158674 179295 158677
rect 178788 158672 179295 158674
rect 178788 158616 179234 158672
rect 179290 158616 179295 158672
rect 178788 158614 179295 158616
rect 178788 158612 178794 158614
rect 179229 158611 179295 158614
rect 179781 158674 179847 158677
rect 180190 158674 180196 158676
rect 179781 158672 180196 158674
rect 179781 158616 179786 158672
rect 179842 158616 180196 158672
rect 179781 158614 180196 158616
rect 179781 158611 179847 158614
rect 180190 158612 180196 158614
rect 180260 158612 180266 158676
rect 181294 158612 181300 158676
rect 181364 158674 181370 158676
rect 181989 158674 182055 158677
rect 181364 158672 182055 158674
rect 181364 158616 181994 158672
rect 182050 158616 182055 158672
rect 181364 158614 182055 158616
rect 181364 158612 181370 158614
rect 181989 158611 182055 158614
rect 182265 158674 182331 158677
rect 182950 158674 182956 158676
rect 182265 158672 182956 158674
rect 182265 158616 182270 158672
rect 182326 158616 182956 158672
rect 182265 158614 182956 158616
rect 182265 158611 182331 158614
rect 182950 158612 182956 158614
rect 183020 158612 183026 158676
rect 186313 158674 186379 158677
rect 187233 158676 187299 158677
rect 186998 158674 187004 158676
rect 186313 158672 187004 158674
rect 186313 158616 186318 158672
rect 186374 158616 187004 158672
rect 186313 158614 187004 158616
rect 186313 158611 186379 158614
rect 186998 158612 187004 158614
rect 187068 158612 187074 158676
rect 187182 158674 187188 158676
rect 187142 158614 187188 158674
rect 187252 158672 187299 158676
rect 187294 158616 187299 158672
rect 187182 158612 187188 158614
rect 187252 158612 187299 158616
rect 187233 158611 187299 158612
rect 187509 158676 187575 158677
rect 187509 158672 187556 158676
rect 187620 158674 187626 158676
rect 187785 158674 187851 158677
rect 188613 158676 188679 158677
rect 188889 158676 188955 158677
rect 188286 158674 188292 158676
rect 187509 158616 187514 158672
rect 187509 158612 187556 158616
rect 187620 158614 187666 158674
rect 187785 158672 188292 158674
rect 187785 158616 187790 158672
rect 187846 158616 188292 158672
rect 187785 158614 188292 158616
rect 187620 158612 187626 158614
rect 187509 158611 187575 158612
rect 187785 158611 187851 158614
rect 188286 158612 188292 158614
rect 188356 158612 188362 158676
rect 188613 158672 188660 158676
rect 188724 158674 188730 158676
rect 188613 158616 188618 158672
rect 188613 158612 188660 158616
rect 188724 158614 188770 158674
rect 188724 158612 188730 158614
rect 188838 158612 188844 158676
rect 188908 158674 188955 158676
rect 189165 158674 189231 158677
rect 189993 158676 190059 158677
rect 189574 158674 189580 158676
rect 188908 158672 189000 158674
rect 188950 158616 189000 158672
rect 188908 158614 189000 158616
rect 189165 158672 189580 158674
rect 189165 158616 189170 158672
rect 189226 158616 189580 158672
rect 189165 158614 189580 158616
rect 188908 158612 188955 158614
rect 188613 158611 188679 158612
rect 188889 158611 188955 158612
rect 189165 158611 189231 158614
rect 189574 158612 189580 158614
rect 189644 158612 189650 158676
rect 189942 158674 189948 158676
rect 189902 158614 189948 158674
rect 190012 158672 190059 158676
rect 190054 158616 190059 158672
rect 189942 158612 189948 158614
rect 190012 158612 190059 158616
rect 189993 158611 190059 158612
rect 190269 158676 190335 158677
rect 190269 158672 190316 158676
rect 190380 158674 190386 158676
rect 190637 158674 190703 158677
rect 191230 158674 191236 158676
rect 190269 158616 190274 158672
rect 190269 158612 190316 158616
rect 190380 158614 190426 158674
rect 190637 158672 191236 158674
rect 190637 158616 190642 158672
rect 190698 158616 191236 158672
rect 190637 158614 191236 158616
rect 190380 158612 190386 158614
rect 190269 158611 190335 158612
rect 190637 158611 190703 158614
rect 191230 158612 191236 158614
rect 191300 158612 191306 158676
rect 150433 158538 150499 158541
rect 151629 158538 151695 158541
rect 150433 158536 168482 158538
rect 150433 158480 150438 158536
rect 150494 158480 151634 158536
rect 151690 158480 168482 158536
rect 150433 158478 168482 158480
rect 150433 158475 150499 158478
rect 151629 158475 151695 158478
rect 164693 158402 164759 158405
rect 165102 158402 165108 158404
rect 164693 158400 165108 158402
rect 164693 158344 164698 158400
rect 164754 158344 165108 158400
rect 164693 158342 165108 158344
rect 164693 158339 164759 158342
rect 165102 158340 165108 158342
rect 165172 158340 165178 158404
rect 168281 158402 168347 158405
rect 166214 158400 168347 158402
rect 166214 158344 168286 158400
rect 168342 158344 168347 158400
rect 166214 158342 168347 158344
rect 168422 158402 168482 158478
rect 168598 158476 168604 158540
rect 168668 158538 168674 158540
rect 169109 158538 169175 158541
rect 168668 158536 169175 158538
rect 168668 158480 169114 158536
rect 169170 158480 169175 158536
rect 168668 158478 169175 158480
rect 168668 158476 168674 158478
rect 169109 158475 169175 158478
rect 171593 158538 171659 158541
rect 172145 158540 172211 158541
rect 171910 158538 171916 158540
rect 171593 158536 171916 158538
rect 171593 158480 171598 158536
rect 171654 158480 171916 158536
rect 171593 158478 171916 158480
rect 171593 158475 171659 158478
rect 171910 158476 171916 158478
rect 171980 158476 171986 158540
rect 172094 158476 172100 158540
rect 172164 158538 172211 158540
rect 172164 158536 172256 158538
rect 172206 158480 172256 158536
rect 172164 158478 172256 158480
rect 172164 158476 172211 158478
rect 174670 158476 174676 158540
rect 174740 158538 174746 158540
rect 174813 158538 174879 158541
rect 174740 158536 174879 158538
rect 174740 158480 174818 158536
rect 174874 158480 174879 158536
rect 174740 158478 174879 158480
rect 174740 158476 174746 158478
rect 172145 158475 172211 158476
rect 174813 158475 174879 158478
rect 174997 158538 175063 158541
rect 175222 158538 175228 158540
rect 174997 158536 175228 158538
rect 174997 158480 175002 158536
rect 175058 158480 175228 158536
rect 174997 158478 175228 158480
rect 174997 158475 175063 158478
rect 175222 158476 175228 158478
rect 175292 158476 175298 158540
rect 175365 158538 175431 158541
rect 176510 158538 176516 158540
rect 175365 158536 176516 158538
rect 175365 158480 175370 158536
rect 175426 158480 176516 158536
rect 175365 158478 176516 158480
rect 175365 158475 175431 158478
rect 176510 158476 176516 158478
rect 176580 158476 176586 158540
rect 186681 158538 186747 158541
rect 187366 158538 187372 158540
rect 186681 158536 187372 158538
rect 186681 158480 186686 158536
rect 186742 158480 187372 158536
rect 186681 158478 187372 158480
rect 186681 158475 186747 158478
rect 187366 158476 187372 158478
rect 187436 158476 187442 158540
rect 191046 158476 191052 158540
rect 191116 158538 191122 158540
rect 191373 158538 191439 158541
rect 191116 158536 191439 158538
rect 191116 158480 191378 158536
rect 191434 158480 191439 158536
rect 191116 158478 191439 158480
rect 191116 158476 191122 158478
rect 191373 158475 191439 158478
rect 192017 158538 192083 158541
rect 192342 158538 192402 158747
rect 192753 158674 192819 158677
rect 194133 158676 194199 158677
rect 194409 158676 194475 158677
rect 193070 158674 193076 158676
rect 192753 158672 193076 158674
rect 192753 158616 192758 158672
rect 192814 158616 193076 158672
rect 192753 158614 193076 158616
rect 192753 158611 192819 158614
rect 193070 158612 193076 158614
rect 193140 158612 193146 158676
rect 194133 158674 194180 158676
rect 194088 158672 194180 158674
rect 194088 158616 194138 158672
rect 194088 158614 194180 158616
rect 194133 158612 194180 158614
rect 194244 158612 194250 158676
rect 194358 158674 194364 158676
rect 194318 158614 194364 158674
rect 194428 158672 194475 158676
rect 194470 158616 194475 158672
rect 194358 158612 194364 158614
rect 194428 158612 194475 158616
rect 195278 158612 195284 158676
rect 195348 158674 195354 158676
rect 195513 158674 195579 158677
rect 195348 158672 195579 158674
rect 195348 158616 195518 158672
rect 195574 158616 195579 158672
rect 195348 158614 195579 158616
rect 195348 158612 195354 158614
rect 194133 158611 194199 158612
rect 194409 158611 194475 158612
rect 195513 158611 195579 158614
rect 196065 158674 196131 158677
rect 196750 158674 196756 158676
rect 196065 158672 196756 158674
rect 196065 158616 196070 158672
rect 196126 158616 196756 158672
rect 196065 158614 196756 158616
rect 196065 158611 196131 158614
rect 196750 158612 196756 158614
rect 196820 158612 196826 158676
rect 196934 158612 196940 158676
rect 197004 158674 197010 158676
rect 197261 158674 197327 158677
rect 197004 158672 197327 158674
rect 197004 158616 197266 158672
rect 197322 158616 197327 158672
rect 197004 158614 197327 158616
rect 197004 158612 197010 158614
rect 197261 158611 197327 158614
rect 198273 158674 198339 158677
rect 198641 158676 198707 158677
rect 198406 158674 198412 158676
rect 198273 158672 198412 158674
rect 198273 158616 198278 158672
rect 198334 158616 198412 158672
rect 198273 158614 198412 158616
rect 198273 158611 198339 158614
rect 198406 158612 198412 158614
rect 198476 158612 198482 158676
rect 198590 158674 198596 158676
rect 198550 158614 198596 158674
rect 198660 158672 198707 158676
rect 198702 158616 198707 158672
rect 198590 158612 198596 158614
rect 198660 158612 198707 158616
rect 198641 158611 198707 158612
rect 199469 158674 199535 158677
rect 199694 158674 199700 158676
rect 199469 158672 199700 158674
rect 199469 158616 199474 158672
rect 199530 158616 199700 158672
rect 199469 158614 199700 158616
rect 199469 158611 199535 158614
rect 199694 158612 199700 158614
rect 199764 158612 199770 158676
rect 200798 158612 200804 158676
rect 200868 158674 200874 158676
rect 201033 158674 201099 158677
rect 202137 158676 202203 158677
rect 202086 158674 202092 158676
rect 200868 158672 201099 158674
rect 200868 158616 201038 158672
rect 201094 158616 201099 158672
rect 200868 158614 201099 158616
rect 202046 158614 202092 158674
rect 202156 158672 202203 158676
rect 202198 158616 202203 158672
rect 200868 158612 200874 158614
rect 201033 158611 201099 158614
rect 202086 158612 202092 158614
rect 202156 158612 202203 158616
rect 202137 158611 202203 158612
rect 203793 158674 203859 158677
rect 204118 158676 204178 158750
rect 205909 158808 270927 158810
rect 205909 158752 205914 158808
rect 205970 158752 270866 158808
rect 270922 158752 270927 158808
rect 205909 158750 270927 158752
rect 205909 158747 205975 158750
rect 270861 158747 270927 158750
rect 203926 158674 203932 158676
rect 203793 158672 203932 158674
rect 203793 158616 203798 158672
rect 203854 158616 203932 158672
rect 203793 158614 203932 158616
rect 203793 158611 203859 158614
rect 203926 158612 203932 158614
rect 203996 158612 204002 158676
rect 204110 158612 204116 158676
rect 204180 158612 204186 158676
rect 204989 158674 205055 158677
rect 205398 158674 205404 158676
rect 204989 158672 205404 158674
rect 204989 158616 204994 158672
rect 205050 158616 205404 158672
rect 204989 158614 205404 158616
rect 204989 158611 205055 158614
rect 205398 158612 205404 158614
rect 205468 158612 205474 158676
rect 206553 158674 206619 158677
rect 206870 158674 206876 158676
rect 206553 158672 206876 158674
rect 206553 158616 206558 158672
rect 206614 158616 206876 158672
rect 206553 158614 206876 158616
rect 206553 158611 206619 158614
rect 206870 158612 206876 158614
rect 206940 158612 206946 158676
rect 192017 158536 192402 158538
rect 192017 158480 192022 158536
rect 192078 158480 192402 158536
rect 192017 158478 192402 158480
rect 192477 158538 192543 158541
rect 192886 158538 192892 158540
rect 192477 158536 192892 158538
rect 192477 158480 192482 158536
rect 192538 158480 192892 158536
rect 192477 158478 192892 158480
rect 192017 158475 192083 158478
rect 192477 158475 192543 158478
rect 192886 158476 192892 158478
rect 192956 158476 192962 158540
rect 193990 158476 193996 158540
rect 194060 158538 194066 158540
rect 194501 158538 194567 158541
rect 194060 158536 194567 158538
rect 194060 158480 194506 158536
rect 194562 158480 194567 158536
rect 194060 158478 194567 158480
rect 194060 158476 194066 158478
rect 194501 158475 194567 158478
rect 195462 158476 195468 158540
rect 195532 158538 195538 158540
rect 195881 158538 195947 158541
rect 195532 158536 195947 158538
rect 195532 158480 195886 158536
rect 195942 158480 195947 158536
rect 195532 158478 195947 158480
rect 195532 158476 195538 158478
rect 195881 158475 195947 158478
rect 199193 158538 199259 158541
rect 199510 158538 199516 158540
rect 199193 158536 199516 158538
rect 199193 158480 199198 158536
rect 199254 158480 199516 158536
rect 199193 158478 199516 158480
rect 199193 158475 199259 158478
rect 199510 158476 199516 158478
rect 199580 158476 199586 158540
rect 200297 158538 200363 158541
rect 201166 158538 201172 158540
rect 200297 158536 201172 158538
rect 200297 158480 200302 158536
rect 200358 158480 201172 158536
rect 200297 158478 201172 158480
rect 200297 158475 200363 158478
rect 201166 158476 201172 158478
rect 201236 158476 201242 158540
rect 201861 158538 201927 158541
rect 202270 158538 202276 158540
rect 201861 158536 202276 158538
rect 201861 158480 201866 158536
rect 201922 158480 202276 158536
rect 201861 158478 202276 158480
rect 201861 158475 201927 158478
rect 202270 158476 202276 158478
rect 202340 158476 202346 158540
rect 203742 158476 203748 158540
rect 203812 158538 203818 158540
rect 204161 158538 204227 158541
rect 203812 158536 204227 158538
rect 203812 158480 204166 158536
rect 204222 158480 204227 158536
rect 203812 158478 204227 158480
rect 203812 158476 203818 158478
rect 204161 158475 204227 158478
rect 206461 158538 206527 158541
rect 208894 158538 208900 158540
rect 206461 158536 208900 158538
rect 206461 158480 206466 158536
rect 206522 158480 208900 158536
rect 206461 158478 208900 158480
rect 206461 158475 206527 158478
rect 208894 158476 208900 158478
rect 208964 158476 208970 158540
rect 168557 158402 168623 158405
rect 168422 158400 168623 158402
rect 168422 158344 168562 158400
rect 168618 158344 168623 158400
rect 168422 158342 168623 158344
rect 161105 158266 161171 158269
rect 166073 158266 166139 158269
rect 161105 158264 166139 158266
rect 161105 158208 161110 158264
rect 161166 158208 166078 158264
rect 166134 158208 166139 158264
rect 161105 158206 166139 158208
rect 161105 158203 161171 158206
rect 166073 158203 166139 158206
rect 159909 158130 159975 158133
rect 166214 158130 166274 158342
rect 168281 158339 168347 158342
rect 168557 158339 168623 158342
rect 168782 158340 168788 158404
rect 168852 158402 168858 158404
rect 169661 158402 169727 158405
rect 168852 158400 169727 158402
rect 168852 158344 169666 158400
rect 169722 158344 169727 158400
rect 168852 158342 169727 158344
rect 168852 158340 168858 158342
rect 169661 158339 169727 158342
rect 174302 158340 174308 158404
rect 174372 158402 174378 158404
rect 175273 158402 175339 158405
rect 174372 158400 175339 158402
rect 174372 158344 175278 158400
rect 175334 158344 175339 158400
rect 174372 158342 175339 158344
rect 174372 158340 174378 158342
rect 175273 158339 175339 158342
rect 190821 158402 190887 158405
rect 191782 158402 191788 158404
rect 190821 158400 191788 158402
rect 190821 158344 190826 158400
rect 190882 158344 191788 158400
rect 190821 158342 191788 158344
rect 190821 158339 190887 158342
rect 191782 158340 191788 158342
rect 191852 158340 191858 158404
rect 193622 158340 193628 158404
rect 193692 158402 193698 158404
rect 194317 158402 194383 158405
rect 193692 158400 194383 158402
rect 193692 158344 194322 158400
rect 194378 158344 194383 158400
rect 193692 158342 194383 158344
rect 193692 158340 193698 158342
rect 194317 158339 194383 158342
rect 194685 158402 194751 158405
rect 195646 158402 195652 158404
rect 194685 158400 195652 158402
rect 194685 158344 194690 158400
rect 194746 158344 195652 158400
rect 194685 158342 195652 158344
rect 194685 158339 194751 158342
rect 195646 158340 195652 158342
rect 195716 158340 195722 158404
rect 198733 158402 198799 158405
rect 199326 158402 199332 158404
rect 198733 158400 199332 158402
rect 198733 158344 198738 158400
rect 198794 158344 199332 158400
rect 198733 158342 199332 158344
rect 198733 158339 198799 158342
rect 199326 158340 199332 158342
rect 199396 158340 199402 158404
rect 200481 158402 200547 158405
rect 201350 158402 201356 158404
rect 200481 158400 201356 158402
rect 200481 158344 200486 158400
rect 200542 158344 201356 158400
rect 200481 158342 201356 158344
rect 200481 158339 200547 158342
rect 201350 158340 201356 158342
rect 201420 158340 201426 158404
rect 203517 158402 203583 158405
rect 204110 158402 204116 158404
rect 203517 158400 204116 158402
rect 203517 158344 203522 158400
rect 203578 158344 204116 158400
rect 203517 158342 204116 158344
rect 203517 158339 203583 158342
rect 204110 158340 204116 158342
rect 204180 158340 204186 158404
rect 205081 158402 205147 158405
rect 209037 158402 209103 158405
rect 205081 158400 209103 158402
rect 205081 158344 205086 158400
rect 205142 158344 209042 158400
rect 209098 158344 209103 158400
rect 205081 158342 209103 158344
rect 205081 158339 205147 158342
rect 209037 158339 209103 158342
rect 166901 158266 166967 158269
rect 172646 158266 172652 158268
rect 166901 158264 172652 158266
rect 166901 158208 166906 158264
rect 166962 158208 172652 158264
rect 166901 158206 172652 158208
rect 166901 158203 166967 158206
rect 172646 158204 172652 158206
rect 172716 158204 172722 158268
rect 175222 158204 175228 158268
rect 175292 158266 175298 158268
rect 175917 158266 175983 158269
rect 175292 158264 175983 158266
rect 175292 158208 175922 158264
rect 175978 158208 175983 158264
rect 175292 158206 175983 158208
rect 175292 158204 175298 158206
rect 175917 158203 175983 158206
rect 191925 158266 191991 158269
rect 192702 158266 192708 158268
rect 191925 158264 192708 158266
rect 191925 158208 191930 158264
rect 191986 158208 192708 158264
rect 191925 158206 192708 158208
rect 191925 158203 191991 158206
rect 192702 158204 192708 158206
rect 192772 158204 192778 158268
rect 193213 158266 193279 158269
rect 194542 158266 194548 158268
rect 193213 158264 194548 158266
rect 193213 158208 193218 158264
rect 193274 158208 194548 158264
rect 193213 158206 194548 158208
rect 193213 158203 193279 158206
rect 194542 158204 194548 158206
rect 194612 158204 194618 158268
rect 199101 158266 199167 158269
rect 200021 158266 200087 158269
rect 199101 158264 200087 158266
rect 199101 158208 199106 158264
rect 199162 158208 200026 158264
rect 200082 158208 200087 158264
rect 199101 158206 200087 158208
rect 199101 158203 199167 158206
rect 200021 158203 200087 158206
rect 202229 158266 202295 158269
rect 202781 158266 202847 158269
rect 202229 158264 202847 158266
rect 202229 158208 202234 158264
rect 202290 158208 202786 158264
rect 202842 158208 202847 158264
rect 202229 158206 202847 158208
rect 202229 158203 202295 158206
rect 202781 158203 202847 158206
rect 204529 158266 204595 158269
rect 209497 158266 209563 158269
rect 204529 158264 209563 158266
rect 204529 158208 204534 158264
rect 204590 158208 209502 158264
rect 209558 158208 209563 158264
rect 204529 158206 209563 158208
rect 204529 158203 204595 158206
rect 209497 158203 209563 158206
rect 172462 158130 172468 158132
rect 159909 158128 166274 158130
rect 159909 158072 159914 158128
rect 159970 158072 166274 158128
rect 159909 158070 166274 158072
rect 166398 158070 172468 158130
rect 159909 158067 159975 158070
rect 158437 157994 158503 157997
rect 166398 157994 166458 158070
rect 172462 158068 172468 158070
rect 172532 158068 172538 158132
rect 192201 158130 192267 158133
rect 193121 158130 193187 158133
rect 192201 158128 193187 158130
rect 192201 158072 192206 158128
rect 192262 158072 193126 158128
rect 193182 158072 193187 158128
rect 192201 158070 193187 158072
rect 192201 158067 192267 158070
rect 193121 158067 193187 158070
rect 196801 158130 196867 158133
rect 199469 158130 199535 158133
rect 196801 158128 199535 158130
rect 196801 158072 196806 158128
rect 196862 158072 199474 158128
rect 199530 158072 199535 158128
rect 196801 158070 199535 158072
rect 196801 158067 196867 158070
rect 199469 158067 199535 158070
rect 201309 158130 201375 158133
rect 202781 158130 202847 158133
rect 201309 158128 202847 158130
rect 201309 158072 201314 158128
rect 201370 158072 202786 158128
rect 202842 158072 202847 158128
rect 201309 158070 202847 158072
rect 201309 158067 201375 158070
rect 202781 158067 202847 158070
rect 203558 158068 203564 158132
rect 203628 158130 203634 158132
rect 203701 158130 203767 158133
rect 203628 158128 203767 158130
rect 203628 158072 203706 158128
rect 203762 158072 203767 158128
rect 203628 158070 203767 158072
rect 203628 158068 203634 158070
rect 203701 158067 203767 158070
rect 206001 158130 206067 158133
rect 206553 158130 206619 158133
rect 206001 158128 206619 158130
rect 206001 158072 206006 158128
rect 206062 158072 206558 158128
rect 206614 158072 206619 158128
rect 206001 158070 206619 158072
rect 206001 158067 206067 158070
rect 206553 158067 206619 158070
rect 207197 158130 207263 158133
rect 208117 158130 208183 158133
rect 227345 158130 227411 158133
rect 207197 158128 227411 158130
rect 207197 158072 207202 158128
rect 207258 158072 208122 158128
rect 208178 158072 227350 158128
rect 227406 158072 227411 158128
rect 207197 158070 227411 158072
rect 207197 158067 207263 158070
rect 208117 158067 208183 158070
rect 227345 158067 227411 158070
rect 167821 157994 167887 157997
rect 158437 157992 166458 157994
rect 158437 157936 158442 157992
rect 158498 157936 166458 157992
rect 158437 157934 166458 157936
rect 166582 157992 167887 157994
rect 166582 157936 167826 157992
rect 167882 157936 167887 157992
rect 166582 157934 167887 157936
rect 158437 157931 158503 157934
rect 158253 157858 158319 157861
rect 166582 157858 166642 157934
rect 167821 157931 167887 157934
rect 178217 157994 178283 157997
rect 179270 157994 179276 157996
rect 178217 157992 179276 157994
rect 178217 157936 178222 157992
rect 178278 157936 179276 157992
rect 178217 157934 179276 157936
rect 178217 157931 178283 157934
rect 179270 157932 179276 157934
rect 179340 157932 179346 157996
rect 180885 157994 180951 157997
rect 181897 157994 181963 157997
rect 180885 157992 181963 157994
rect 180885 157936 180890 157992
rect 180946 157936 181902 157992
rect 181958 157936 181963 157992
rect 180885 157934 181963 157936
rect 180885 157931 180951 157934
rect 181897 157931 181963 157934
rect 192017 157994 192083 157997
rect 196617 157994 196683 157997
rect 192017 157992 196683 157994
rect 192017 157936 192022 157992
rect 192078 157936 196622 157992
rect 196678 157936 196683 157992
rect 192017 157934 196683 157936
rect 192017 157931 192083 157934
rect 196617 157931 196683 157934
rect 199285 157994 199351 157997
rect 203190 157994 203196 157996
rect 199285 157992 203196 157994
rect 199285 157936 199290 157992
rect 199346 157936 203196 157992
rect 199285 157934 203196 157936
rect 199285 157931 199351 157934
rect 203190 157932 203196 157934
rect 203260 157932 203266 157996
rect 208669 157994 208735 157997
rect 245878 157994 245884 157996
rect 208669 157992 245884 157994
rect 208669 157936 208674 157992
rect 208730 157936 245884 157992
rect 208669 157934 245884 157936
rect 208669 157931 208735 157934
rect 245878 157932 245884 157934
rect 245948 157932 245954 157996
rect 158253 157856 166642 157858
rect 158253 157800 158258 157856
rect 158314 157800 166642 157856
rect 158253 157798 166642 157800
rect 166993 157858 167059 157861
rect 168230 157858 168236 157860
rect 166993 157856 168236 157858
rect 166993 157800 166998 157856
rect 167054 157800 168236 157856
rect 166993 157798 168236 157800
rect 158253 157795 158319 157798
rect 166993 157795 167059 157798
rect 168230 157796 168236 157798
rect 168300 157796 168306 157860
rect 168557 157858 168623 157861
rect 174445 157858 174511 157861
rect 168557 157856 174511 157858
rect 168557 157800 168562 157856
rect 168618 157800 174450 157856
rect 174506 157800 174511 157856
rect 168557 157798 174511 157800
rect 168557 157795 168623 157798
rect 174445 157795 174511 157798
rect 176929 157858 176995 157861
rect 177798 157858 177804 157860
rect 176929 157856 177804 157858
rect 176929 157800 176934 157856
rect 176990 157800 177804 157856
rect 176929 157798 177804 157800
rect 176929 157795 176995 157798
rect 177798 157796 177804 157798
rect 177868 157796 177874 157860
rect 178401 157858 178467 157861
rect 179086 157858 179092 157860
rect 178401 157856 179092 157858
rect 178401 157800 178406 157856
rect 178462 157800 179092 157856
rect 178401 157798 179092 157800
rect 178401 157795 178467 157798
rect 179086 157796 179092 157798
rect 179156 157858 179162 157860
rect 179229 157858 179295 157861
rect 179156 157856 179295 157858
rect 179156 157800 179234 157856
rect 179290 157800 179295 157856
rect 179156 157798 179295 157800
rect 179156 157796 179162 157798
rect 179229 157795 179295 157798
rect 202137 157858 202203 157861
rect 238150 157858 238156 157860
rect 202137 157856 238156 157858
rect 202137 157800 202142 157856
rect 202198 157800 238156 157856
rect 202137 157798 238156 157800
rect 202137 157795 202203 157798
rect 238150 157796 238156 157798
rect 238220 157796 238226 157860
rect 157333 157722 157399 157725
rect 158161 157722 158227 157725
rect 166901 157722 166967 157725
rect 157333 157720 166967 157722
rect 157333 157664 157338 157720
rect 157394 157664 158166 157720
rect 158222 157664 166906 157720
rect 166962 157664 166967 157720
rect 157333 157662 166967 157664
rect 157333 157659 157399 157662
rect 158161 157659 158227 157662
rect 166901 157659 166967 157662
rect 168281 157722 168347 157725
rect 174353 157722 174419 157725
rect 168281 157720 174419 157722
rect 168281 157664 168286 157720
rect 168342 157664 174358 157720
rect 174414 157664 174419 157720
rect 168281 157662 174419 157664
rect 168281 157659 168347 157662
rect 174353 157659 174419 157662
rect 177246 157660 177252 157724
rect 177316 157722 177322 157724
rect 177849 157722 177915 157725
rect 178953 157724 179019 157725
rect 177316 157720 177915 157722
rect 177316 157664 177854 157720
rect 177910 157664 177915 157720
rect 177316 157662 177915 157664
rect 177316 157660 177322 157662
rect 177849 157659 177915 157662
rect 178902 157660 178908 157724
rect 178972 157722 179019 157724
rect 179505 157722 179571 157725
rect 180006 157722 180012 157724
rect 178972 157720 179064 157722
rect 179014 157664 179064 157720
rect 178972 157662 179064 157664
rect 179505 157720 180012 157722
rect 179505 157664 179510 157720
rect 179566 157664 180012 157720
rect 179505 157662 180012 157664
rect 178972 157660 179019 157662
rect 178953 157659 179019 157660
rect 179505 157659 179571 157662
rect 180006 157660 180012 157662
rect 180076 157722 180082 157724
rect 180609 157722 180675 157725
rect 180076 157720 180675 157722
rect 180076 157664 180614 157720
rect 180670 157664 180675 157720
rect 180076 157662 180675 157664
rect 180076 157660 180082 157662
rect 180609 157659 180675 157662
rect 181110 157660 181116 157724
rect 181180 157722 181186 157724
rect 181437 157722 181503 157725
rect 210969 157722 211035 157725
rect 181180 157720 181503 157722
rect 181180 157664 181442 157720
rect 181498 157664 181503 157720
rect 181180 157662 181503 157664
rect 181180 157660 181186 157662
rect 181437 157659 181503 157662
rect 195930 157720 211035 157722
rect 195930 157664 210974 157720
rect 211030 157664 211035 157720
rect 195930 157662 211035 157664
rect 160737 157586 160803 157589
rect 163497 157586 163563 157589
rect 195930 157586 195990 157662
rect 210969 157659 211035 157662
rect 160737 157584 168850 157586
rect 160737 157528 160742 157584
rect 160798 157528 163502 157584
rect 163558 157528 168850 157584
rect 160737 157526 168850 157528
rect 160737 157523 160803 157526
rect 163497 157523 163563 157526
rect 155769 157450 155835 157453
rect 163037 157450 163103 157453
rect 164601 157452 164667 157453
rect 155769 157448 163103 157450
rect 155769 157392 155774 157448
rect 155830 157392 163042 157448
rect 163098 157392 163103 157448
rect 155769 157390 163103 157392
rect 155769 157387 155835 157390
rect 163037 157387 163103 157390
rect 164550 157388 164556 157452
rect 164620 157450 164667 157452
rect 164620 157448 164712 157450
rect 164662 157392 164712 157448
rect 164620 157390 164712 157392
rect 164620 157388 164667 157390
rect 164601 157387 164667 157388
rect 157241 157314 157307 157317
rect 164366 157314 164372 157316
rect 157241 157312 164372 157314
rect 157241 157256 157246 157312
rect 157302 157256 164372 157312
rect 157241 157254 164372 157256
rect 157241 157251 157307 157254
rect 164366 157252 164372 157254
rect 164436 157314 164442 157316
rect 164969 157314 165035 157317
rect 164436 157312 165035 157314
rect 164436 157256 164974 157312
rect 165030 157256 165035 157312
rect 164436 157254 165035 157256
rect 168790 157314 168850 157526
rect 169526 157526 195990 157586
rect 202137 157586 202203 157589
rect 202454 157586 202460 157588
rect 202137 157584 202460 157586
rect 202137 157528 202142 157584
rect 202198 157528 202460 157584
rect 202137 157526 202460 157528
rect 169526 157314 169586 157526
rect 202137 157523 202203 157526
rect 202454 157524 202460 157526
rect 202524 157524 202530 157588
rect 206737 157586 206803 157589
rect 206870 157586 206876 157588
rect 206737 157584 206876 157586
rect 206737 157528 206742 157584
rect 206798 157528 206876 157584
rect 206737 157526 206876 157528
rect 206737 157523 206803 157526
rect 206870 157524 206876 157526
rect 206940 157524 206946 157588
rect 176142 157450 176148 157452
rect 171182 157390 176148 157450
rect 168790 157254 169586 157314
rect 171041 157314 171107 157317
rect 171182 157314 171242 157390
rect 176142 157388 176148 157390
rect 176212 157388 176218 157452
rect 177205 157450 177271 157453
rect 177430 157450 177436 157452
rect 177205 157448 177436 157450
rect 177205 157392 177210 157448
rect 177266 157392 177436 157448
rect 177205 157390 177436 157392
rect 177205 157387 177271 157390
rect 177430 157388 177436 157390
rect 177500 157388 177506 157452
rect 177614 157388 177620 157452
rect 177684 157450 177690 157452
rect 177757 157450 177823 157453
rect 177684 157448 177823 157450
rect 177684 157392 177762 157448
rect 177818 157392 177823 157448
rect 177684 157390 177823 157392
rect 177684 157388 177690 157390
rect 177757 157387 177823 157390
rect 178309 157450 178375 157453
rect 179965 157452 180031 157453
rect 179086 157450 179092 157452
rect 178309 157448 179092 157450
rect 178309 157392 178314 157448
rect 178370 157392 179092 157448
rect 178309 157390 179092 157392
rect 178309 157387 178375 157390
rect 179086 157388 179092 157390
rect 179156 157388 179162 157452
rect 179965 157448 180012 157452
rect 180076 157450 180082 157452
rect 180333 157450 180399 157453
rect 180558 157450 180564 157452
rect 179965 157392 179970 157448
rect 179965 157388 180012 157392
rect 180076 157390 180122 157450
rect 180333 157448 180564 157450
rect 180333 157392 180338 157448
rect 180394 157392 180564 157448
rect 180333 157390 180564 157392
rect 180076 157388 180082 157390
rect 179965 157387 180031 157388
rect 180333 157387 180399 157390
rect 180558 157388 180564 157390
rect 180628 157388 180634 157452
rect 181478 157388 181484 157452
rect 181548 157450 181554 157452
rect 181713 157450 181779 157453
rect 181548 157448 181779 157450
rect 181548 157392 181718 157448
rect 181774 157392 181779 157448
rect 181548 157390 181779 157392
rect 181548 157388 181554 157390
rect 181713 157387 181779 157390
rect 183645 157450 183711 157453
rect 185025 157452 185091 157453
rect 184238 157450 184244 157452
rect 183645 157448 184244 157450
rect 183645 157392 183650 157448
rect 183706 157392 184244 157448
rect 183645 157390 184244 157392
rect 183645 157387 183711 157390
rect 184238 157388 184244 157390
rect 184308 157388 184314 157452
rect 184974 157450 184980 157452
rect 184934 157390 184980 157450
rect 185044 157448 185091 157452
rect 185086 157392 185091 157448
rect 184974 157388 184980 157390
rect 185044 157388 185091 157392
rect 185025 157387 185091 157388
rect 200205 157450 200271 157453
rect 200665 157450 200731 157453
rect 200205 157448 200731 157450
rect 200205 157392 200210 157448
rect 200266 157392 200670 157448
rect 200726 157392 200731 157448
rect 200205 157390 200731 157392
rect 200205 157387 200271 157390
rect 200665 157387 200731 157390
rect 205633 157450 205699 157453
rect 206645 157450 206711 157453
rect 205633 157448 206711 157450
rect 205633 157392 205638 157448
rect 205694 157392 206650 157448
rect 206706 157392 206711 157448
rect 205633 157390 206711 157392
rect 205633 157387 205699 157390
rect 206645 157387 206711 157390
rect 171041 157312 171242 157314
rect 171041 157256 171046 157312
rect 171102 157256 171242 157312
rect 171041 157254 171242 157256
rect 172513 157314 172579 157317
rect 173014 157314 173020 157316
rect 172513 157312 173020 157314
rect 172513 157256 172518 157312
rect 172574 157256 173020 157312
rect 172513 157254 173020 157256
rect 164436 157252 164442 157254
rect 164969 157251 165035 157254
rect 171041 157251 171107 157254
rect 172513 157251 172579 157254
rect 173014 157252 173020 157254
rect 173084 157252 173090 157316
rect 191414 157252 191420 157316
rect 191484 157314 191490 157316
rect 191649 157314 191715 157317
rect 191484 157312 191715 157314
rect 191484 157256 191654 157312
rect 191710 157256 191715 157312
rect 191484 157254 191715 157256
rect 191484 157252 191490 157254
rect 191649 157251 191715 157254
rect 198181 157314 198247 157317
rect 290641 157314 290707 157317
rect 291101 157314 291167 157317
rect 198181 157312 291167 157314
rect 198181 157256 198186 157312
rect 198242 157256 290646 157312
rect 290702 157256 291106 157312
rect 291162 157256 291167 157312
rect 198181 157254 291167 157256
rect 198181 157251 198247 157254
rect 290641 157251 290707 157254
rect 291101 157251 291167 157254
rect 162485 157178 162551 157181
rect 162894 157178 162900 157180
rect 162485 157176 162900 157178
rect 162485 157120 162490 157176
rect 162546 157120 162900 157176
rect 162485 157118 162900 157120
rect 162485 157115 162551 157118
rect 162894 157116 162900 157118
rect 162964 157116 162970 157180
rect 202045 157178 202111 157181
rect 274909 157178 274975 157181
rect 202045 157176 274975 157178
rect 202045 157120 202050 157176
rect 202106 157120 274914 157176
rect 274970 157120 274975 157176
rect 202045 157118 274975 157120
rect 202045 157115 202111 157118
rect 274909 157115 274975 157118
rect 156689 157042 156755 157045
rect 157149 157042 157215 157045
rect 166349 157042 166415 157045
rect 156689 157040 166415 157042
rect 156689 156984 156694 157040
rect 156750 156984 157154 157040
rect 157210 156984 166354 157040
rect 166410 156984 166415 157040
rect 156689 156982 166415 156984
rect 156689 156979 156755 156982
rect 157149 156979 157215 156982
rect 166349 156979 166415 156982
rect 199837 157042 199903 157045
rect 270585 157042 270651 157045
rect 199837 157040 270651 157042
rect 199837 156984 199842 157040
rect 199898 156984 270590 157040
rect 270646 156984 270651 157040
rect 199837 156982 270651 156984
rect 199837 156979 199903 156982
rect 270585 156979 270651 156982
rect 155493 156906 155559 156909
rect 167453 156906 167519 156909
rect 155493 156904 167519 156906
rect 155493 156848 155498 156904
rect 155554 156848 167458 156904
rect 167514 156848 167519 156904
rect 155493 156846 167519 156848
rect 155493 156843 155559 156846
rect 167453 156843 167519 156846
rect 175406 156844 175412 156908
rect 175476 156906 175482 156908
rect 216305 156906 216371 156909
rect 175476 156904 216371 156906
rect 175476 156848 216310 156904
rect 216366 156848 216371 156904
rect 175476 156846 216371 156848
rect 175476 156844 175482 156846
rect 216305 156843 216371 156846
rect 156781 156770 156847 156773
rect 167126 156770 167132 156772
rect 156781 156768 167132 156770
rect 156781 156712 156786 156768
rect 156842 156712 167132 156768
rect 156781 156710 167132 156712
rect 156781 156707 156847 156710
rect 167126 156708 167132 156710
rect 167196 156770 167202 156772
rect 167269 156770 167335 156773
rect 167196 156768 167335 156770
rect 167196 156712 167274 156768
rect 167330 156712 167335 156768
rect 167196 156710 167335 156712
rect 167196 156708 167202 156710
rect 167269 156707 167335 156710
rect 200113 156770 200179 156773
rect 239765 156770 239831 156773
rect 200113 156768 239831 156770
rect 200113 156712 200118 156768
rect 200174 156712 239770 156768
rect 239826 156712 239831 156768
rect 200113 156710 239831 156712
rect 200113 156707 200179 156710
rect 239765 156707 239831 156710
rect 193489 156634 193555 156637
rect 208485 156634 208551 156637
rect 193489 156632 208551 156634
rect 193489 156576 193494 156632
rect 193550 156576 208490 156632
rect 208546 156576 208551 156632
rect 193489 156574 208551 156576
rect 193489 156571 193555 156574
rect 208485 156571 208551 156574
rect 291101 156634 291167 156637
rect 431217 156634 431283 156637
rect 291101 156632 431283 156634
rect 291101 156576 291106 156632
rect 291162 156576 431222 156632
rect 431278 156576 431283 156632
rect 291101 156574 431283 156576
rect 291101 156571 291167 156574
rect 431217 156571 431283 156574
rect 171225 155954 171291 155957
rect 175406 155954 175412 155956
rect 171225 155952 175412 155954
rect 171225 155896 171230 155952
rect 171286 155896 175412 155952
rect 171225 155894 175412 155896
rect 171225 155891 171291 155894
rect 175406 155892 175412 155894
rect 175476 155892 175482 155956
rect 200389 155954 200455 155957
rect 211705 155954 211771 155957
rect 200389 155952 211771 155954
rect 200389 155896 200394 155952
rect 200450 155896 211710 155952
rect 211766 155896 211771 155952
rect 200389 155894 211771 155896
rect 200389 155891 200455 155894
rect 211705 155891 211771 155894
rect 203742 155756 203748 155820
rect 203812 155818 203818 155820
rect 268326 155818 268332 155820
rect 203812 155758 268332 155818
rect 203812 155756 203818 155758
rect 268326 155756 268332 155758
rect 268396 155756 268402 155820
rect 179270 155620 179276 155684
rect 179340 155682 179346 155684
rect 219985 155682 220051 155685
rect 179340 155680 220051 155682
rect 179340 155624 219990 155680
rect 220046 155624 220051 155680
rect 179340 155622 220051 155624
rect 179340 155620 179346 155622
rect 219985 155619 220051 155622
rect 205357 155546 205423 155549
rect 236821 155546 236887 155549
rect 205357 155544 236887 155546
rect 205357 155488 205362 155544
rect 205418 155488 236826 155544
rect 236882 155488 236887 155544
rect 205357 155486 236887 155488
rect 205357 155483 205423 155486
rect 236821 155483 236887 155486
rect 201493 155410 201559 155413
rect 233182 155410 233188 155412
rect 201493 155408 233188 155410
rect 201493 155352 201498 155408
rect 201554 155352 233188 155408
rect 201493 155350 233188 155352
rect 201493 155347 201559 155350
rect 233182 155348 233188 155350
rect 233252 155348 233258 155412
rect 206461 155274 206527 155277
rect 206921 155274 206987 155277
rect 220445 155274 220511 155277
rect 206461 155272 220511 155274
rect 206461 155216 206466 155272
rect 206522 155216 206926 155272
rect 206982 155216 220450 155272
rect 220506 155216 220511 155272
rect 206461 155214 220511 155216
rect 206461 155211 206527 155214
rect 206921 155211 206987 155214
rect 220445 155211 220511 155214
rect 195697 155138 195763 155141
rect 200941 155138 201007 155141
rect 195697 155136 201007 155138
rect 195697 155080 195702 155136
rect 195758 155080 200946 155136
rect 201002 155080 201007 155136
rect 195697 155078 201007 155080
rect 195697 155075 195763 155078
rect 200941 155075 201007 155078
rect 203425 155138 203491 155141
rect 204069 155138 204135 155141
rect 270769 155138 270835 155141
rect 203425 155136 270835 155138
rect 203425 155080 203430 155136
rect 203486 155080 204074 155136
rect 204130 155080 270774 155136
rect 270830 155080 270835 155136
rect 203425 155078 270835 155080
rect 203425 155075 203491 155078
rect 204069 155075 204135 155078
rect 270769 155075 270835 155078
rect 197537 154594 197603 154597
rect 204253 154594 204319 154597
rect 197537 154592 204319 154594
rect 197537 154536 197542 154592
rect 197598 154536 204258 154592
rect 204314 154536 204319 154592
rect 197537 154534 204319 154536
rect 197537 154531 197603 154534
rect 204253 154531 204319 154534
rect 205173 154458 205239 154461
rect 276105 154458 276171 154461
rect 205173 154456 276171 154458
rect 205173 154400 205178 154456
rect 205234 154400 276110 154456
rect 276166 154400 276171 154456
rect 205173 154398 276171 154400
rect 205173 154395 205239 154398
rect 276105 154395 276171 154398
rect 205909 154322 205975 154325
rect 273846 154322 273852 154324
rect 205909 154320 273852 154322
rect 205909 154264 205914 154320
rect 205970 154264 273852 154320
rect 205909 154262 273852 154264
rect 205909 154259 205975 154262
rect 273846 154260 273852 154262
rect 273916 154322 273922 154324
rect 273916 154262 277410 154322
rect 273916 154260 273922 154262
rect 203149 154186 203215 154189
rect 262949 154186 263015 154189
rect 203149 154184 263015 154186
rect 203149 154128 203154 154184
rect 203210 154128 262954 154184
rect 263010 154128 263015 154184
rect 203149 154126 263015 154128
rect 203149 154123 203215 154126
rect 262949 154123 263015 154126
rect 131113 154050 131179 154053
rect 157333 154050 157399 154053
rect 131113 154048 157399 154050
rect 131113 153992 131118 154048
rect 131174 153992 157338 154048
rect 157394 153992 157399 154048
rect 131113 153990 157399 153992
rect 131113 153987 131179 153990
rect 157333 153987 157399 153990
rect 199694 153988 199700 154052
rect 199764 154050 199770 154052
rect 240910 154050 240916 154052
rect 199764 153990 240916 154050
rect 199764 153988 199770 153990
rect 240910 153988 240916 153990
rect 240980 153988 240986 154052
rect 71773 153914 71839 153917
rect 155861 153914 155927 153917
rect 71773 153912 155927 153914
rect 71773 153856 71778 153912
rect 71834 153856 155866 153912
rect 155922 153856 155927 153912
rect 71773 153854 155927 153856
rect 71773 153851 71839 153854
rect 155861 153851 155927 153854
rect 198365 153914 198431 153917
rect 236637 153914 236703 153917
rect 198365 153912 236703 153914
rect 198365 153856 198370 153912
rect 198426 153856 236642 153912
rect 236698 153856 236703 153912
rect 198365 153854 236703 153856
rect 198365 153851 198431 153854
rect 236637 153851 236703 153854
rect 6913 153778 6979 153781
rect 155401 153778 155467 153781
rect 6913 153776 155467 153778
rect 6913 153720 6918 153776
rect 6974 153720 155406 153776
rect 155462 153720 155467 153776
rect 6913 153718 155467 153720
rect 277350 153778 277410 154262
rect 557533 153778 557599 153781
rect 277350 153776 557599 153778
rect 277350 153720 557538 153776
rect 557594 153720 557599 153776
rect 277350 153718 557599 153720
rect 6913 153715 6979 153718
rect 155401 153715 155467 153718
rect 557533 153715 557599 153718
rect 186998 153580 187004 153644
rect 187068 153642 187074 153644
rect 208669 153642 208735 153645
rect 187068 153640 208735 153642
rect 187068 153584 208674 153640
rect 208730 153584 208735 153640
rect 187068 153582 208735 153584
rect 187068 153580 187074 153582
rect 208669 153579 208735 153582
rect 196382 153172 196388 153236
rect 196452 153234 196458 153236
rect 197261 153234 197327 153237
rect 196452 153232 197327 153234
rect 196452 153176 197266 153232
rect 197322 153176 197327 153232
rect 196452 153174 197327 153176
rect 196452 153172 196458 153174
rect 197261 153171 197327 153174
rect 154573 153098 154639 153101
rect 158253 153098 158319 153101
rect 154573 153096 158319 153098
rect 154573 153040 154578 153096
rect 154634 153040 158258 153096
rect 158314 153040 158319 153096
rect 154573 153038 158319 153040
rect 154573 153035 154639 153038
rect 158253 153035 158319 153038
rect 196934 153036 196940 153100
rect 197004 153098 197010 153100
rect 276289 153098 276355 153101
rect 197004 153096 276355 153098
rect 197004 153040 276294 153096
rect 276350 153040 276355 153096
rect 197004 153038 276355 153040
rect 197004 153036 197010 153038
rect 276289 153035 276355 153038
rect 195462 152900 195468 152964
rect 195532 152962 195538 152964
rect 273345 152962 273411 152965
rect 195532 152960 273411 152962
rect 195532 152904 273350 152960
rect 273406 152904 273411 152960
rect 195532 152902 273411 152904
rect 195532 152900 195538 152902
rect 273345 152899 273411 152902
rect 204161 152826 204227 152829
rect 262857 152826 262923 152829
rect 204161 152824 262923 152826
rect 204161 152768 204166 152824
rect 204222 152768 262862 152824
rect 262918 152768 262923 152824
rect 204161 152766 262923 152768
rect 204161 152763 204227 152766
rect 262857 152763 262923 152766
rect 194542 152628 194548 152692
rect 194612 152690 194618 152692
rect 253473 152690 253539 152693
rect 194612 152688 253539 152690
rect 194612 152632 253478 152688
rect 253534 152632 253539 152688
rect 194612 152630 253539 152632
rect 194612 152628 194618 152630
rect 253473 152627 253539 152630
rect 579889 152690 579955 152693
rect 583520 152690 584960 152780
rect 579889 152688 584960 152690
rect 579889 152632 579894 152688
rect 579950 152632 584960 152688
rect 579889 152630 584960 152632
rect 579889 152627 579955 152630
rect 198038 152492 198044 152556
rect 198108 152554 198114 152556
rect 198590 152554 198596 152556
rect 198108 152494 198596 152554
rect 198108 152492 198114 152494
rect 198590 152492 198596 152494
rect 198660 152554 198666 152556
rect 239673 152554 239739 152557
rect 198660 152552 239739 152554
rect 198660 152496 239678 152552
rect 239734 152496 239739 152552
rect 583520 152540 584960 152630
rect 198660 152494 239739 152496
rect 198660 152492 198666 152494
rect 239673 152491 239739 152494
rect 51073 152418 51139 152421
rect 156689 152418 156755 152421
rect 51073 152416 156755 152418
rect 51073 152360 51078 152416
rect 51134 152360 156694 152416
rect 156750 152360 156755 152416
rect 51073 152358 156755 152360
rect 51073 152355 51139 152358
rect 156689 152355 156755 152358
rect 193990 152356 193996 152420
rect 194060 152418 194066 152420
rect 217593 152418 217659 152421
rect 194060 152416 217659 152418
rect 194060 152360 217598 152416
rect 217654 152360 217659 152416
rect 194060 152358 217659 152360
rect 194060 152356 194066 152358
rect 217593 152355 217659 152358
rect 195278 152220 195284 152284
rect 195348 152282 195354 152284
rect 213453 152282 213519 152285
rect 195348 152280 213519 152282
rect 195348 152224 213458 152280
rect 213514 152224 213519 152280
rect 195348 152222 213519 152224
rect 195348 152220 195354 152222
rect 213453 152219 213519 152222
rect 193397 151738 193463 151741
rect 284017 151738 284083 151741
rect 193397 151736 284083 151738
rect 193397 151680 193402 151736
rect 193458 151680 284022 151736
rect 284078 151680 284083 151736
rect 193397 151678 284083 151680
rect 193397 151675 193463 151678
rect 284017 151675 284083 151678
rect 201125 151602 201191 151605
rect 284477 151602 284543 151605
rect 201125 151600 284543 151602
rect 201125 151544 201130 151600
rect 201186 151544 284482 151600
rect 284538 151544 284543 151600
rect 201125 151542 284543 151544
rect 201125 151539 201191 151542
rect 284477 151539 284543 151542
rect 197169 151466 197235 151469
rect 257613 151466 257679 151469
rect 197169 151464 257679 151466
rect 197169 151408 197174 151464
rect 197230 151408 257618 151464
rect 257674 151408 257679 151464
rect 197169 151406 257679 151408
rect 197169 151403 197235 151406
rect 257613 151403 257679 151406
rect 179086 151268 179092 151332
rect 179156 151330 179162 151332
rect 238201 151330 238267 151333
rect 179156 151328 238267 151330
rect 179156 151272 238206 151328
rect 238262 151272 238267 151328
rect 179156 151270 238267 151272
rect 179156 151268 179162 151270
rect 238201 151267 238267 151270
rect 192109 151194 192175 151197
rect 234337 151194 234403 151197
rect 192109 151192 234403 151194
rect 192109 151136 192114 151192
rect 192170 151136 234342 151192
rect 234398 151136 234403 151192
rect 192109 151134 234403 151136
rect 192109 151131 192175 151134
rect 234337 151131 234403 151134
rect 284017 151194 284083 151197
rect 376017 151194 376083 151197
rect 284017 151192 376083 151194
rect 284017 151136 284022 151192
rect 284078 151136 376022 151192
rect 376078 151136 376083 151192
rect 284017 151134 376083 151136
rect 284017 151131 284083 151134
rect 376017 151131 376083 151134
rect 284477 151058 284543 151061
rect 498285 151058 498351 151061
rect 284477 151056 498351 151058
rect 284477 151000 284482 151056
rect 284538 151000 498290 151056
rect 498346 151000 498351 151056
rect 284477 150998 498351 151000
rect 284477 150995 284543 150998
rect 498285 150995 498351 150998
rect 151905 150514 151971 150517
rect 159449 150514 159515 150517
rect 151905 150512 159515 150514
rect 151905 150456 151910 150512
rect 151966 150456 159454 150512
rect 159510 150456 159515 150512
rect 151905 150454 159515 150456
rect 151905 150451 151971 150454
rect 159449 150451 159515 150454
rect 203609 150378 203675 150381
rect 298185 150378 298251 150381
rect 299381 150378 299447 150381
rect 203609 150376 299447 150378
rect 203609 150320 203614 150376
rect 203670 150320 298190 150376
rect 298246 150320 299386 150376
rect 299442 150320 299447 150376
rect 203609 150318 299447 150320
rect 203609 150315 203675 150318
rect 298185 150315 298251 150318
rect 299381 150315 299447 150318
rect 196750 150180 196756 150244
rect 196820 150242 196826 150244
rect 256141 150242 256207 150245
rect 196820 150240 256207 150242
rect 196820 150184 256146 150240
rect 256202 150184 256207 150240
rect 196820 150182 256207 150184
rect 196820 150180 196826 150182
rect 256141 150179 256207 150182
rect 177614 150044 177620 150108
rect 177684 150106 177690 150108
rect 222009 150106 222075 150109
rect 177684 150104 222075 150106
rect 177684 150048 222014 150104
rect 222070 150048 222075 150104
rect 177684 150046 222075 150048
rect 177684 150044 177690 150046
rect 222009 150043 222075 150046
rect 127617 149970 127683 149973
rect 155309 149970 155375 149973
rect 127617 149968 155375 149970
rect -960 149834 480 149924
rect 127617 149912 127622 149968
rect 127678 149912 155314 149968
rect 155370 149912 155375 149968
rect 127617 149910 155375 149912
rect 127617 149907 127683 149910
rect 155309 149907 155375 149910
rect 177430 149908 177436 149972
rect 177500 149970 177506 149972
rect 215293 149970 215359 149973
rect 177500 149968 215359 149970
rect 177500 149912 215298 149968
rect 215354 149912 215359 149968
rect 177500 149910 215359 149912
rect 177500 149908 177506 149910
rect 215293 149907 215359 149910
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 100753 149834 100819 149837
rect 154021 149834 154087 149837
rect 100753 149832 154087 149834
rect 100753 149776 100758 149832
rect 100814 149776 154026 149832
rect 154082 149776 154087 149832
rect 100753 149774 154087 149776
rect 100753 149771 100819 149774
rect 154021 149771 154087 149774
rect 177798 149772 177804 149836
rect 177868 149834 177874 149836
rect 214097 149834 214163 149837
rect 177868 149832 214163 149834
rect 177868 149776 214102 149832
rect 214158 149776 214163 149832
rect 177868 149774 214163 149776
rect 177868 149772 177874 149774
rect 214097 149771 214163 149774
rect 71037 149698 71103 149701
rect 156505 149698 156571 149701
rect 71037 149696 156571 149698
rect 71037 149640 71042 149696
rect 71098 149640 156510 149696
rect 156566 149640 156571 149696
rect 71037 149638 156571 149640
rect 71037 149635 71103 149638
rect 156505 149635 156571 149638
rect 299381 149698 299447 149701
rect 529933 149698 529999 149701
rect 299381 149696 529999 149698
rect 299381 149640 299386 149696
rect 299442 149640 529938 149696
rect 529994 149640 529999 149696
rect 299381 149638 529999 149640
rect 299381 149635 299447 149638
rect 529933 149635 529999 149638
rect 204713 149018 204779 149021
rect 282453 149018 282519 149021
rect 204713 149016 282519 149018
rect 204713 148960 204718 149016
rect 204774 148960 282458 149016
rect 282514 148960 282519 149016
rect 204713 148958 282519 148960
rect 204713 148955 204779 148958
rect 282453 148955 282519 148958
rect 201401 148882 201467 148885
rect 274633 148882 274699 148885
rect 201401 148880 277410 148882
rect 201401 148824 201406 148880
rect 201462 148824 274638 148880
rect 274694 148824 277410 148880
rect 201401 148822 277410 148824
rect 201401 148819 201467 148822
rect 274633 148819 274699 148822
rect 198917 148746 198983 148749
rect 269113 148746 269179 148749
rect 198917 148744 269179 148746
rect 198917 148688 198922 148744
rect 198978 148688 269118 148744
rect 269174 148688 269179 148744
rect 198917 148686 269179 148688
rect 198917 148683 198983 148686
rect 269113 148683 269179 148686
rect 116577 148610 116643 148613
rect 158069 148610 158135 148613
rect 116577 148608 158135 148610
rect 116577 148552 116582 148608
rect 116638 148552 158074 148608
rect 158130 148552 158135 148608
rect 116577 148550 158135 148552
rect 116577 148547 116643 148550
rect 158069 148547 158135 148550
rect 202781 148610 202847 148613
rect 269757 148610 269823 148613
rect 202781 148608 269823 148610
rect 202781 148552 202786 148608
rect 202842 148552 269762 148608
rect 269818 148552 269823 148608
rect 202781 148550 269823 148552
rect 202781 148547 202847 148550
rect 269757 148547 269823 148550
rect 103513 148474 103579 148477
rect 156873 148474 156939 148477
rect 103513 148472 156939 148474
rect 103513 148416 103518 148472
rect 103574 148416 156878 148472
rect 156934 148416 156939 148472
rect 103513 148414 156939 148416
rect 103513 148411 103579 148414
rect 156873 148411 156939 148414
rect 170990 148412 170996 148476
rect 171060 148474 171066 148476
rect 230974 148474 230980 148476
rect 171060 148414 230980 148474
rect 171060 148412 171066 148414
rect 230974 148412 230980 148414
rect 231044 148412 231050 148476
rect 277350 148474 277410 148822
rect 500953 148474 501019 148477
rect 277350 148472 501019 148474
rect 277350 148416 500958 148472
rect 501014 148416 501019 148472
rect 277350 148414 501019 148416
rect 500953 148411 501019 148414
rect 31017 148338 31083 148341
rect 151169 148338 151235 148341
rect 31017 148336 151235 148338
rect 31017 148280 31022 148336
rect 31078 148280 151174 148336
rect 151230 148280 151235 148336
rect 31017 148278 151235 148280
rect 31017 148275 31083 148278
rect 151169 148275 151235 148278
rect 282453 148338 282519 148341
rect 543733 148338 543799 148341
rect 282453 148336 543799 148338
rect 282453 148280 282458 148336
rect 282514 148280 543738 148336
rect 543794 148280 543799 148336
rect 282453 148278 543799 148280
rect 282453 148275 282519 148278
rect 543733 148275 543799 148278
rect 153101 147658 153167 147661
rect 168966 147658 168972 147660
rect 142110 147656 168972 147658
rect 142110 147600 153106 147656
rect 153162 147600 168972 147656
rect 142110 147598 168972 147600
rect 89713 147114 89779 147117
rect 142110 147114 142170 147598
rect 153101 147595 153167 147598
rect 168966 147596 168972 147598
rect 169036 147596 169042 147660
rect 206093 147658 206159 147661
rect 295333 147658 295399 147661
rect 206093 147656 295399 147658
rect 206093 147600 206098 147656
rect 206154 147600 295338 147656
rect 295394 147600 295399 147656
rect 206093 147598 295399 147600
rect 206093 147595 206159 147598
rect 295333 147595 295399 147598
rect 234153 147522 234219 147525
rect 173390 147520 234219 147522
rect 173390 147464 234158 147520
rect 234214 147464 234219 147520
rect 173390 147462 234219 147464
rect 172973 147250 173039 147253
rect 173390 147252 173450 147462
rect 234153 147459 234219 147462
rect 203926 147324 203932 147388
rect 203996 147386 204002 147388
rect 264278 147386 264284 147388
rect 203996 147326 264284 147386
rect 203996 147324 204002 147326
rect 264278 147324 264284 147326
rect 264348 147324 264354 147388
rect 173382 147250 173388 147252
rect 172973 147248 173388 147250
rect 172973 147192 172978 147248
rect 173034 147192 173388 147248
rect 172973 147190 173388 147192
rect 172973 147187 173039 147190
rect 173382 147188 173388 147190
rect 173452 147188 173458 147252
rect 174486 147188 174492 147252
rect 174556 147250 174562 147252
rect 232589 147250 232655 147253
rect 174556 147248 232655 147250
rect 174556 147192 232594 147248
rect 232650 147192 232655 147248
rect 174556 147190 232655 147192
rect 174556 147188 174562 147190
rect 232589 147187 232655 147190
rect 89713 147112 142170 147114
rect 89713 147056 89718 147112
rect 89774 147056 142170 147112
rect 89713 147054 142170 147056
rect 89713 147051 89779 147054
rect 173198 147052 173204 147116
rect 173268 147114 173274 147116
rect 227253 147114 227319 147117
rect 173268 147112 227319 147114
rect 173268 147056 227258 147112
rect 227314 147056 227319 147112
rect 173268 147054 227319 147056
rect 173268 147052 173274 147054
rect 227253 147051 227319 147054
rect 16573 146978 16639 146981
rect 162894 146978 162900 146980
rect 16573 146976 162900 146978
rect 16573 146920 16578 146976
rect 16634 146920 162900 146976
rect 16573 146918 162900 146920
rect 16573 146915 16639 146918
rect 162894 146916 162900 146918
rect 162964 146916 162970 146980
rect 187366 146916 187372 146980
rect 187436 146978 187442 146980
rect 211889 146978 211955 146981
rect 187436 146976 211955 146978
rect 187436 146920 211894 146976
rect 211950 146920 211955 146976
rect 187436 146918 211955 146920
rect 187436 146916 187442 146918
rect 211889 146915 211955 146918
rect 295333 146978 295399 146981
rect 296069 146978 296135 146981
rect 561673 146978 561739 146981
rect 295333 146976 561739 146978
rect 295333 146920 295338 146976
rect 295394 146920 296074 146976
rect 296130 146920 561678 146976
rect 561734 146920 561739 146976
rect 295333 146918 561739 146920
rect 295333 146915 295399 146918
rect 296069 146915 296135 146918
rect 561673 146915 561739 146918
rect 154389 146298 154455 146301
rect 168782 146298 168788 146300
rect 142110 146296 168788 146298
rect 142110 146240 154394 146296
rect 154450 146240 168788 146296
rect 142110 146238 168788 146240
rect 93853 145754 93919 145757
rect 142110 145754 142170 146238
rect 154389 146235 154455 146238
rect 168782 146236 168788 146238
rect 168852 146236 168858 146300
rect 173893 146298 173959 146301
rect 175222 146298 175228 146300
rect 173893 146296 175228 146298
rect 173893 146240 173898 146296
rect 173954 146240 175228 146296
rect 173893 146238 175228 146240
rect 173893 146235 173959 146238
rect 175222 146236 175228 146238
rect 175292 146236 175298 146300
rect 184238 146236 184244 146300
rect 184308 146298 184314 146300
rect 212533 146298 212599 146301
rect 184308 146296 212599 146298
rect 184308 146240 212538 146296
rect 212594 146240 212599 146296
rect 184308 146238 212599 146240
rect 184308 146236 184314 146238
rect 212533 146235 212599 146238
rect 154481 146162 154547 146165
rect 168598 146162 168604 146164
rect 93853 145752 142170 145754
rect 93853 145696 93858 145752
rect 93914 145696 142170 145752
rect 93853 145694 142170 145696
rect 151770 146160 168604 146162
rect 151770 146104 154486 146160
rect 154542 146104 168604 146160
rect 151770 146102 168604 146104
rect 93853 145691 93919 145694
rect 88977 145618 89043 145621
rect 151770 145618 151830 146102
rect 154481 146099 154547 146102
rect 168598 146100 168604 146102
rect 168668 146100 168674 146164
rect 201166 146100 201172 146164
rect 201236 146162 201242 146164
rect 260046 146162 260052 146164
rect 201236 146102 260052 146162
rect 201236 146100 201242 146102
rect 260046 146100 260052 146102
rect 260116 146100 260122 146164
rect 180006 145964 180012 146028
rect 180076 146026 180082 146028
rect 218053 146026 218119 146029
rect 180076 146024 218119 146026
rect 180076 145968 218058 146024
rect 218114 145968 218119 146024
rect 180076 145966 218119 145968
rect 180076 145964 180082 145966
rect 218053 145963 218119 145966
rect 176510 145828 176516 145892
rect 176580 145890 176586 145892
rect 214189 145890 214255 145893
rect 176580 145888 214255 145890
rect 176580 145832 214194 145888
rect 214250 145832 214255 145888
rect 176580 145830 214255 145832
rect 176580 145828 176586 145830
rect 214189 145827 214255 145830
rect 205398 145692 205404 145756
rect 205468 145754 205474 145756
rect 267774 145754 267780 145756
rect 205468 145694 267780 145754
rect 205468 145692 205474 145694
rect 267774 145692 267780 145694
rect 267844 145692 267850 145756
rect 88977 145616 151830 145618
rect 88977 145560 88982 145616
rect 89038 145560 151830 145616
rect 88977 145558 151830 145560
rect 218053 145618 218119 145621
rect 218789 145618 218855 145621
rect 226333 145618 226399 145621
rect 218053 145616 226399 145618
rect 218053 145560 218058 145616
rect 218114 145560 218794 145616
rect 218850 145560 226338 145616
rect 226394 145560 226399 145616
rect 218053 145558 226399 145560
rect 88977 145555 89043 145558
rect 218053 145555 218119 145558
rect 218789 145555 218855 145558
rect 226333 145555 226399 145558
rect 202965 144802 203031 144805
rect 203885 144802 203951 144805
rect 202965 144800 203994 144802
rect 202965 144744 202970 144800
rect 203026 144744 203890 144800
rect 203946 144744 203994 144800
rect 202965 144742 203994 144744
rect 202965 144739 203031 144742
rect 203885 144739 203994 144742
rect 204110 144740 204116 144804
rect 204180 144802 204186 144804
rect 278865 144802 278931 144805
rect 204180 144800 278931 144802
rect 204180 144744 278870 144800
rect 278926 144744 278931 144800
rect 204180 144742 278931 144744
rect 204180 144740 204186 144742
rect 278865 144739 278931 144742
rect 203934 144666 203994 144739
rect 262438 144666 262444 144668
rect 203934 144606 262444 144666
rect 262438 144604 262444 144606
rect 262508 144604 262514 144668
rect 228633 144530 228699 144533
rect 171090 144528 228699 144530
rect 171090 144472 228638 144528
rect 228694 144472 228699 144528
rect 171090 144470 228699 144472
rect 107653 144258 107719 144261
rect 169661 144258 169727 144261
rect 171090 144258 171150 144470
rect 228633 144467 228699 144470
rect 191782 144332 191788 144396
rect 191852 144394 191858 144396
rect 217409 144394 217475 144397
rect 191852 144392 217475 144394
rect 191852 144336 217414 144392
rect 217470 144336 217475 144392
rect 191852 144334 217475 144336
rect 191852 144332 191858 144334
rect 217409 144331 217475 144334
rect 107653 144256 171150 144258
rect 107653 144200 107658 144256
rect 107714 144200 169666 144256
rect 169722 144200 171150 144256
rect 107653 144198 171150 144200
rect 107653 144195 107719 144198
rect 169661 144195 169727 144198
rect 191230 144196 191236 144260
rect 191300 144258 191306 144260
rect 215937 144258 216003 144261
rect 191300 144256 216003 144258
rect 191300 144200 215942 144256
rect 215998 144200 216003 144256
rect 191300 144198 216003 144200
rect 191300 144196 191306 144198
rect 215937 144195 216003 144198
rect 33133 144122 33199 144125
rect 164366 144122 164372 144124
rect 33133 144120 164372 144122
rect 33133 144064 33138 144120
rect 33194 144064 164372 144120
rect 33133 144062 164372 144064
rect 33133 144059 33199 144062
rect 164366 144060 164372 144062
rect 164436 144060 164442 144124
rect 178902 144060 178908 144124
rect 178972 144122 178978 144124
rect 212533 144122 212599 144125
rect 178972 144120 212599 144122
rect 178972 144064 212538 144120
rect 212594 144064 212599 144120
rect 178972 144062 212599 144064
rect 178972 144060 178978 144062
rect 212533 144059 212599 144062
rect 174302 143380 174308 143444
rect 174372 143442 174378 143444
rect 174629 143442 174695 143445
rect 174372 143440 174695 143442
rect 174372 143384 174634 143440
rect 174690 143384 174695 143440
rect 174372 143382 174695 143384
rect 174372 143380 174378 143382
rect 174629 143379 174695 143382
rect 200205 143442 200271 143445
rect 201309 143442 201375 143445
rect 200205 143440 201375 143442
rect 200205 143384 200210 143440
rect 200266 143384 201314 143440
rect 201370 143384 201375 143440
rect 200205 143382 201375 143384
rect 200205 143379 200271 143382
rect 201309 143379 201375 143382
rect 202086 143380 202092 143444
rect 202156 143442 202162 143444
rect 202689 143442 202755 143445
rect 202156 143440 202755 143442
rect 202156 143384 202694 143440
rect 202750 143384 202755 143440
rect 202156 143382 202755 143384
rect 202156 143380 202162 143382
rect 202689 143379 202755 143382
rect 200798 143244 200804 143308
rect 200868 143306 200874 143308
rect 261702 143306 261708 143308
rect 200868 143246 261708 143306
rect 200868 143244 200874 143246
rect 261702 143244 261708 143246
rect 261772 143244 261778 143308
rect 173014 143108 173020 143172
rect 173084 143170 173090 143172
rect 232681 143170 232747 143173
rect 173084 143168 232747 143170
rect 173084 143112 232686 143168
rect 232742 143112 232747 143168
rect 173084 143110 232747 143112
rect 173084 143108 173090 143110
rect 232681 143107 232747 143110
rect 201309 143034 201375 143037
rect 259678 143034 259684 143036
rect 201309 143032 259684 143034
rect 201309 142976 201314 143032
rect 201370 142976 259684 143032
rect 201309 142974 259684 142976
rect 201309 142971 201375 142974
rect 259678 142972 259684 142974
rect 259748 142972 259754 143036
rect 202270 142836 202276 142900
rect 202340 142898 202346 142900
rect 261518 142898 261524 142900
rect 202340 142838 261524 142898
rect 202340 142836 202346 142838
rect 261518 142836 261524 142838
rect 261588 142836 261594 142900
rect 263593 142898 263659 142901
rect 264094 142898 264100 142900
rect 263593 142896 264100 142898
rect 263593 142840 263598 142896
rect 263654 142840 264100 142896
rect 263593 142838 264100 142840
rect 263593 142835 263659 142838
rect 264094 142836 264100 142838
rect 264164 142836 264170 142900
rect 171726 142700 171732 142764
rect 171796 142762 171802 142764
rect 172278 142762 172284 142764
rect 171796 142702 172284 142762
rect 171796 142700 171802 142702
rect 172278 142700 172284 142702
rect 172348 142762 172354 142764
rect 221457 142762 221523 142765
rect 172348 142760 221523 142762
rect 172348 142704 221462 142760
rect 221518 142704 221523 142760
rect 172348 142702 221523 142704
rect 172348 142700 172354 142702
rect 221457 142699 221523 142702
rect 189942 142564 189948 142628
rect 190012 142626 190018 142628
rect 221641 142626 221707 142629
rect 190012 142624 221707 142626
rect 190012 142568 221646 142624
rect 221702 142568 221707 142624
rect 190012 142566 221707 142568
rect 190012 142564 190018 142566
rect 221641 142563 221707 142566
rect 201350 142292 201356 142356
rect 201420 142354 201426 142356
rect 272057 142354 272123 142357
rect 201420 142352 272123 142354
rect 201420 142296 272062 142352
rect 272118 142296 272123 142352
rect 201420 142294 272123 142296
rect 201420 142292 201426 142294
rect 272057 142291 272123 142294
rect 260833 142218 260899 142221
rect 261334 142218 261340 142220
rect 260833 142216 261340 142218
rect 260833 142160 260838 142216
rect 260894 142160 261340 142216
rect 260833 142158 261340 142160
rect 260833 142155 260899 142158
rect 261334 142156 261340 142158
rect 261404 142156 261410 142220
rect 172421 142082 172487 142085
rect 232630 142082 232636 142084
rect 172421 142080 232636 142082
rect 172421 142024 172426 142080
rect 172482 142024 232636 142080
rect 172421 142022 232636 142024
rect 172421 142019 172487 142022
rect 232630 142020 232636 142022
rect 232700 142020 232706 142084
rect 188838 141884 188844 141948
rect 188908 141946 188914 141948
rect 249374 141946 249380 141948
rect 188908 141886 249380 141946
rect 188908 141884 188914 141886
rect 249374 141884 249380 141886
rect 249444 141884 249450 141948
rect 187550 141748 187556 141812
rect 187620 141810 187626 141812
rect 238017 141810 238083 141813
rect 187620 141808 238083 141810
rect 187620 141752 238022 141808
rect 238078 141752 238083 141808
rect 187620 141750 238083 141752
rect 187620 141748 187626 141750
rect 238017 141747 238083 141750
rect 187182 141612 187188 141676
rect 187252 141674 187258 141676
rect 232773 141674 232839 141677
rect 187252 141672 232839 141674
rect 187252 141616 232778 141672
rect 232834 141616 232839 141672
rect 187252 141614 232839 141616
rect 187252 141612 187258 141614
rect 232773 141611 232839 141614
rect 147673 141538 147739 141541
rect 174486 141538 174492 141540
rect 147673 141536 174492 141538
rect 147673 141480 147678 141536
rect 147734 141480 174492 141536
rect 147673 141478 174492 141480
rect 147673 141475 147739 141478
rect 174486 141476 174492 141478
rect 174556 141476 174562 141540
rect 191414 141476 191420 141540
rect 191484 141538 191490 141540
rect 235349 141538 235415 141541
rect 191484 141536 235415 141538
rect 191484 141480 235354 141536
rect 235410 141480 235415 141536
rect 191484 141478 235415 141480
rect 191484 141476 191490 141478
rect 235349 141475 235415 141478
rect 110413 141402 110479 141405
rect 170254 141402 170260 141404
rect 110413 141400 170260 141402
rect 110413 141344 110418 141400
rect 110474 141344 170260 141400
rect 110413 141342 170260 141344
rect 110413 141339 110479 141342
rect 170254 141340 170260 141342
rect 170324 141340 170330 141404
rect 188654 141340 188660 141404
rect 188724 141402 188730 141404
rect 224309 141402 224375 141405
rect 188724 141400 224375 141402
rect 188724 141344 224314 141400
rect 224370 141344 224375 141400
rect 188724 141342 224375 141344
rect 188724 141340 188730 141342
rect 224309 141339 224375 141342
rect 190310 141204 190316 141268
rect 190380 141266 190386 141268
rect 223113 141266 223179 141269
rect 190380 141264 223179 141266
rect 190380 141208 223118 141264
rect 223174 141208 223179 141264
rect 190380 141206 223179 141208
rect 190380 141204 190386 141206
rect 223113 141203 223179 141206
rect 191046 140796 191052 140860
rect 191116 140858 191122 140860
rect 191649 140858 191715 140861
rect 191116 140856 191715 140858
rect 191116 140800 191654 140856
rect 191710 140800 191715 140856
rect 191116 140798 191715 140800
rect 191116 140796 191122 140798
rect 191649 140795 191715 140798
rect 150525 140722 150591 140725
rect 151721 140722 151787 140725
rect 168414 140722 168420 140724
rect 150525 140720 168420 140722
rect 150525 140664 150530 140720
rect 150586 140664 151726 140720
rect 151782 140664 168420 140720
rect 150525 140662 168420 140664
rect 150525 140659 150591 140662
rect 151721 140659 151787 140662
rect 168414 140660 168420 140662
rect 168484 140660 168490 140724
rect 181478 140660 181484 140724
rect 181548 140722 181554 140724
rect 242198 140722 242204 140724
rect 181548 140662 242204 140722
rect 181548 140660 181554 140662
rect 242198 140660 242204 140662
rect 242268 140660 242274 140724
rect 177246 140524 177252 140588
rect 177316 140586 177322 140588
rect 237966 140586 237972 140588
rect 177316 140526 237972 140586
rect 177316 140524 177322 140526
rect 237966 140524 237972 140526
rect 238036 140524 238042 140588
rect 189758 140388 189764 140452
rect 189828 140450 189834 140452
rect 189993 140450 190059 140453
rect 246430 140450 246436 140452
rect 189828 140448 190059 140450
rect 189828 140392 189998 140448
rect 190054 140392 190059 140448
rect 189828 140390 190059 140392
rect 189828 140388 189834 140390
rect 189993 140387 190059 140390
rect 195286 140390 246436 140450
rect 187509 140314 187575 140317
rect 195286 140314 195346 140390
rect 246430 140388 246436 140390
rect 246500 140388 246506 140452
rect 187509 140312 195346 140314
rect 187509 140256 187514 140312
rect 187570 140256 195346 140312
rect 187509 140254 195346 140256
rect 195421 140314 195487 140317
rect 240726 140314 240732 140316
rect 195421 140312 240732 140314
rect 195421 140256 195426 140312
rect 195482 140256 240732 140312
rect 195421 140254 240732 140256
rect 187509 140251 187575 140254
rect 195421 140251 195487 140254
rect 240726 140252 240732 140254
rect 240796 140252 240802 140316
rect 121453 140178 121519 140181
rect 172421 140178 172487 140181
rect 121453 140176 172487 140178
rect 121453 140120 121458 140176
rect 121514 140120 172426 140176
rect 172482 140120 172487 140176
rect 121453 140118 172487 140120
rect 121453 140115 121519 140118
rect 172421 140115 172487 140118
rect 187601 140178 187667 140181
rect 242014 140178 242020 140180
rect 187601 140176 242020 140178
rect 187601 140120 187606 140176
rect 187662 140120 242020 140176
rect 187601 140118 242020 140120
rect 187601 140115 187667 140118
rect 242014 140116 242020 140118
rect 242084 140116 242090 140180
rect 80053 140042 80119 140045
rect 150525 140042 150591 140045
rect 80053 140040 150591 140042
rect 80053 139984 80058 140040
rect 80114 139984 150530 140040
rect 150586 139984 150591 140040
rect 80053 139982 150591 139984
rect 80053 139979 80119 139982
rect 150525 139979 150591 139982
rect 188286 139980 188292 140044
rect 188356 140042 188362 140044
rect 229921 140042 229987 140045
rect 188356 140040 229987 140042
rect 188356 139984 229926 140040
rect 229982 139984 229987 140040
rect 188356 139982 229987 139984
rect 188356 139980 188362 139982
rect 229921 139979 229987 139982
rect 178718 139844 178724 139908
rect 178788 139906 178794 139908
rect 216673 139906 216739 139909
rect 178788 139904 216739 139906
rect 178788 139848 216678 139904
rect 216734 139848 216739 139904
rect 178788 139846 216739 139848
rect 178788 139844 178794 139846
rect 216673 139843 216739 139846
rect 184974 139708 184980 139772
rect 185044 139770 185050 139772
rect 195421 139770 195487 139773
rect 185044 139768 195487 139770
rect 185044 139712 195426 139768
rect 195482 139712 195487 139768
rect 185044 139710 195487 139712
rect 185044 139708 185050 139710
rect 195421 139707 195487 139710
rect 198406 139708 198412 139772
rect 198476 139770 198482 139772
rect 198641 139770 198707 139773
rect 198476 139768 198707 139770
rect 198476 139712 198646 139768
rect 198702 139712 198707 139768
rect 198476 139710 198707 139712
rect 198476 139708 198482 139710
rect 198641 139707 198707 139710
rect 186313 139634 186379 139637
rect 187509 139634 187575 139637
rect 186313 139632 187575 139634
rect 186313 139576 186318 139632
rect 186374 139576 187514 139632
rect 187570 139576 187575 139632
rect 186313 139574 187575 139576
rect 186313 139571 186379 139574
rect 187509 139571 187575 139574
rect 186681 139498 186747 139501
rect 187601 139498 187667 139501
rect 186681 139496 187667 139498
rect 186681 139440 186686 139496
rect 186742 139440 187606 139496
rect 187662 139440 187667 139496
rect 186681 139438 187667 139440
rect 186681 139435 186747 139438
rect 187601 139435 187667 139438
rect 168649 139362 168715 139365
rect 169017 139362 169083 139365
rect 234654 139362 234660 139364
rect 168649 139360 234660 139362
rect 168649 139304 168654 139360
rect 168710 139304 169022 139360
rect 169078 139304 234660 139360
rect 168649 139302 234660 139304
rect 168649 139299 168715 139302
rect 169017 139299 169083 139302
rect 234654 139300 234660 139302
rect 234724 139300 234730 139364
rect 580257 139362 580323 139365
rect 583520 139362 584960 139452
rect 580257 139360 584960 139362
rect 580257 139304 580262 139360
rect 580318 139304 584960 139360
rect 580257 139302 584960 139304
rect 580257 139299 580323 139302
rect 195646 139164 195652 139228
rect 195716 139226 195722 139228
rect 258717 139226 258783 139229
rect 195716 139224 258783 139226
rect 195716 139168 258722 139224
rect 258778 139168 258783 139224
rect 583520 139212 584960 139302
rect 195716 139166 258783 139168
rect 195716 139164 195722 139166
rect 258717 139163 258783 139166
rect 168833 139090 168899 139093
rect 169201 139090 169267 139093
rect 230422 139090 230428 139092
rect 168833 139088 230428 139090
rect 168833 139032 168838 139088
rect 168894 139032 169206 139088
rect 169262 139032 230428 139088
rect 168833 139030 230428 139032
rect 168833 139027 168899 139030
rect 169201 139027 169267 139030
rect 230422 139028 230428 139030
rect 230492 139028 230498 139092
rect 167126 138892 167132 138956
rect 167196 138954 167202 138956
rect 168230 138954 168236 138956
rect 167196 138894 168236 138954
rect 167196 138892 167202 138894
rect 168230 138892 168236 138894
rect 168300 138954 168306 138956
rect 226425 138954 226491 138957
rect 168300 138952 226491 138954
rect 168300 138896 226430 138952
rect 226486 138896 226491 138952
rect 168300 138894 226491 138896
rect 168300 138892 168306 138894
rect 226425 138891 226491 138894
rect 62113 138682 62179 138685
rect 166942 138682 166948 138684
rect 62113 138680 166948 138682
rect 62113 138624 62118 138680
rect 62174 138624 166948 138680
rect 62113 138622 166948 138624
rect 62113 138619 62179 138622
rect 166942 138620 166948 138622
rect 167012 138620 167018 138684
rect 177798 138620 177804 138684
rect 177868 138682 177874 138684
rect 186313 138682 186379 138685
rect 177868 138680 186379 138682
rect 177868 138624 186318 138680
rect 186374 138624 186379 138680
rect 177868 138622 186379 138624
rect 177868 138620 177874 138622
rect 186313 138619 186379 138622
rect 166165 138002 166231 138005
rect 227161 138002 227227 138005
rect 166165 138000 227227 138002
rect 166165 137944 166170 138000
rect 166226 137944 227166 138000
rect 227222 137944 227227 138000
rect 166165 137942 227227 137944
rect 166165 137939 166231 137942
rect 227161 137939 227227 137942
rect 194174 137804 194180 137868
rect 194244 137866 194250 137868
rect 254577 137866 254643 137869
rect 194244 137864 254643 137866
rect 194244 137808 254582 137864
rect 254638 137808 254643 137864
rect 194244 137806 254643 137808
rect 194244 137804 194250 137806
rect 254577 137803 254643 137806
rect 193070 137668 193076 137732
rect 193140 137730 193146 137732
rect 253289 137730 253355 137733
rect 193140 137728 253355 137730
rect 193140 137672 253294 137728
rect 253350 137672 253355 137728
rect 193140 137670 253355 137672
rect 193140 137668 193146 137670
rect 253289 137667 253355 137670
rect 166165 137596 166231 137597
rect 166165 137594 166212 137596
rect 166120 137592 166212 137594
rect 166120 137536 166170 137592
rect 166120 137534 166212 137536
rect 166165 137532 166212 137534
rect 166276 137532 166282 137596
rect 192702 137532 192708 137596
rect 192772 137594 192778 137596
rect 251766 137594 251772 137596
rect 192772 137534 251772 137594
rect 192772 137532 192778 137534
rect 251766 137532 251772 137534
rect 251836 137532 251842 137596
rect 166165 137531 166231 137532
rect 192518 137396 192524 137460
rect 192588 137458 192594 137460
rect 250294 137458 250300 137460
rect 192588 137398 250300 137458
rect 192588 137396 192594 137398
rect 250294 137396 250300 137398
rect 250364 137396 250370 137460
rect 59353 137322 59419 137325
rect 167126 137322 167132 137324
rect 59353 137320 167132 137322
rect 59353 137264 59358 137320
rect 59414 137264 167132 137320
rect 59353 137262 167132 137264
rect 59353 137259 59419 137262
rect 167126 137260 167132 137262
rect 167196 137260 167202 137324
rect 194358 137260 194364 137324
rect 194428 137322 194434 137324
rect 239489 137322 239555 137325
rect 194428 137320 239555 137322
rect 194428 137264 239494 137320
rect 239550 137264 239555 137320
rect 194428 137262 239555 137264
rect 194428 137260 194434 137262
rect 239489 137259 239555 137262
rect 192886 137124 192892 137188
rect 192956 137186 192962 137188
rect 236494 137186 236500 137188
rect 192956 137126 236500 137186
rect 192956 137124 192962 137126
rect 236494 137124 236500 137126
rect 236564 137124 236570 137188
rect -960 136778 480 136868
rect 3049 136778 3115 136781
rect -960 136776 3115 136778
rect -960 136720 3054 136776
rect 3110 136720 3115 136776
rect -960 136718 3115 136720
rect -960 136628 480 136718
rect 3049 136715 3115 136718
rect 177430 136580 177436 136644
rect 177500 136642 177506 136644
rect 180149 136642 180215 136645
rect 177500 136640 180215 136642
rect 177500 136584 180154 136640
rect 180210 136584 180215 136640
rect 177500 136582 180215 136584
rect 177500 136580 177506 136582
rect 180149 136579 180215 136582
rect 271822 136580 271828 136644
rect 271892 136642 271898 136644
rect 272241 136642 272307 136645
rect 271892 136640 272307 136642
rect 271892 136584 272246 136640
rect 272302 136584 272307 136640
rect 271892 136582 272307 136584
rect 271892 136580 271898 136582
rect 272241 136579 272307 136582
rect 143625 135962 143691 135965
rect 173382 135962 173388 135964
rect 143625 135960 173388 135962
rect 143625 135904 143630 135960
rect 143686 135904 173388 135960
rect 143625 135902 173388 135904
rect 143625 135899 143691 135902
rect 173382 135900 173388 135902
rect 173452 135900 173458 135964
rect 180190 135900 180196 135964
rect 180260 135962 180266 135964
rect 223573 135962 223639 135965
rect 180260 135960 223639 135962
rect 180260 135904 223578 135960
rect 223634 135904 223639 135960
rect 180260 135902 223639 135904
rect 180260 135900 180266 135902
rect 223573 135899 223639 135902
rect 126973 134466 127039 134469
rect 171726 134466 171732 134468
rect 126973 134464 171732 134466
rect 126973 134408 126978 134464
rect 127034 134408 171732 134464
rect 126973 134406 171732 134408
rect 126973 134403 127039 134406
rect 171726 134404 171732 134406
rect 171796 134404 171802 134468
rect 52453 131746 52519 131749
rect 166206 131746 166212 131748
rect 52453 131744 166212 131746
rect 52453 131688 52458 131744
rect 52514 131688 166212 131744
rect 52453 131686 166212 131688
rect 52453 131683 52519 131686
rect 166206 131684 166212 131686
rect 166276 131684 166282 131748
rect 199326 131684 199332 131748
rect 199396 131746 199402 131748
rect 468477 131746 468543 131749
rect 199396 131744 468543 131746
rect 199396 131688 468482 131744
rect 468538 131688 468543 131744
rect 199396 131686 468543 131688
rect 199396 131684 199402 131686
rect 468477 131683 468543 131686
rect 171777 131202 171843 131205
rect 175774 131202 175780 131204
rect 171777 131200 175780 131202
rect 171777 131144 171782 131200
rect 171838 131144 175780 131200
rect 171777 131142 175780 131144
rect 171777 131139 171843 131142
rect 175774 131140 175780 131142
rect 175844 131140 175850 131204
rect 32397 130386 32463 130389
rect 164366 130386 164372 130388
rect 32397 130384 164372 130386
rect 32397 130328 32402 130384
rect 32458 130328 164372 130384
rect 32397 130326 164372 130328
rect 32397 130323 32463 130326
rect 164366 130324 164372 130326
rect 164436 130324 164442 130388
rect 180374 130324 180380 130388
rect 180444 130386 180450 130388
rect 226425 130386 226491 130389
rect 180444 130384 226491 130386
rect 180444 130328 226430 130384
rect 226486 130328 226491 130384
rect 180444 130326 226491 130328
rect 180444 130324 180450 130326
rect 226425 130323 226491 130326
rect 182950 127604 182956 127668
rect 183020 127666 183026 127668
rect 255313 127666 255379 127669
rect 183020 127664 255379 127666
rect 183020 127608 255318 127664
rect 255374 127608 255379 127664
rect 183020 127606 255379 127608
rect 183020 127604 183026 127606
rect 255313 127603 255379 127606
rect 181110 126924 181116 126988
rect 181180 126986 181186 126988
rect 233877 126986 233943 126989
rect 181180 126984 233943 126986
rect 181180 126928 233882 126984
rect 233938 126928 233943 126984
rect 181180 126926 233943 126928
rect 181180 126924 181186 126926
rect 233877 126923 233943 126926
rect 136633 126306 136699 126309
rect 173198 126306 173204 126308
rect 136633 126304 173204 126306
rect 136633 126248 136638 126304
rect 136694 126248 173204 126304
rect 136633 126246 173204 126248
rect 136633 126243 136699 126246
rect 173198 126244 173204 126246
rect 173268 126244 173274 126308
rect 233877 126306 233943 126309
rect 244273 126306 244339 126309
rect 233877 126304 244339 126306
rect 233877 126248 233882 126304
rect 233938 126248 244278 126304
rect 244334 126248 244339 126304
rect 233877 126246 244339 126248
rect 233877 126243 233943 126246
rect 244273 126243 244339 126246
rect 580533 126034 580599 126037
rect 583520 126034 584960 126124
rect 580533 126032 584960 126034
rect 580533 125976 580538 126032
rect 580594 125976 584960 126032
rect 580533 125974 584960 125976
rect 580533 125971 580599 125974
rect 583520 125884 584960 125974
rect 199510 125428 199516 125492
rect 199580 125490 199586 125492
rect 292573 125490 292639 125493
rect 293217 125490 293283 125493
rect 199580 125488 293283 125490
rect 199580 125432 292578 125488
rect 292634 125432 293222 125488
rect 293278 125432 293283 125488
rect 199580 125430 293283 125432
rect 199580 125428 199586 125430
rect 292573 125427 292639 125430
rect 293217 125427 293283 125430
rect 182582 124748 182588 124812
rect 182652 124810 182658 124812
rect 258717 124810 258783 124813
rect 182652 124808 258783 124810
rect 182652 124752 258722 124808
rect 258778 124752 258783 124808
rect 182652 124750 258783 124752
rect 182652 124748 182658 124750
rect 258717 124747 258783 124750
rect 292573 124810 292639 124813
rect 472617 124810 472683 124813
rect 292573 124808 472683 124810
rect 292573 124752 292578 124808
rect 292634 124752 472622 124808
rect 472678 124752 472683 124808
rect 292573 124750 472683 124752
rect 292573 124747 292639 124750
rect 472617 124747 472683 124750
rect 180558 124068 180564 124132
rect 180628 124130 180634 124132
rect 229001 124130 229067 124133
rect 180628 124128 229067 124130
rect 180628 124072 229006 124128
rect 229062 124072 229067 124128
rect 180628 124070 229067 124072
rect 180628 124068 180634 124070
rect 229001 124067 229067 124070
rect -960 123572 480 123812
rect 229001 122906 229067 122909
rect 230473 122906 230539 122909
rect 229001 122904 230539 122906
rect 229001 122848 229006 122904
rect 229062 122848 230478 122904
rect 230534 122848 230539 122904
rect 229001 122846 230539 122848
rect 229001 122843 229067 122846
rect 230473 122843 230539 122846
rect 182766 122164 182772 122228
rect 182836 122226 182842 122228
rect 265617 122226 265683 122229
rect 182836 122224 265683 122226
rect 182836 122168 265622 122224
rect 265678 122168 265683 122224
rect 182836 122166 265683 122168
rect 182836 122164 182842 122166
rect 265617 122163 265683 122166
rect 193990 122028 193996 122092
rect 194060 122090 194066 122092
rect 412633 122090 412699 122093
rect 194060 122088 412699 122090
rect 194060 122032 412638 122088
rect 412694 122032 412699 122088
rect 194060 122030 412699 122032
rect 194060 122028 194066 122030
rect 412633 122027 412699 122030
rect 177614 120804 177620 120868
rect 177684 120866 177690 120868
rect 196617 120866 196683 120869
rect 177684 120864 196683 120866
rect 177684 120808 196622 120864
rect 196678 120808 196683 120864
rect 177684 120806 196683 120808
rect 177684 120804 177690 120806
rect 196617 120803 196683 120806
rect 195278 120668 195284 120732
rect 195348 120730 195354 120732
rect 426433 120730 426499 120733
rect 195348 120728 426499 120730
rect 195348 120672 426438 120728
rect 426494 120672 426499 120728
rect 195348 120670 426499 120672
rect 195348 120668 195354 120670
rect 426433 120667 426499 120670
rect 187182 119444 187188 119508
rect 187252 119506 187258 119508
rect 318793 119506 318859 119509
rect 187252 119504 318859 119506
rect 187252 119448 318798 119504
rect 318854 119448 318859 119504
rect 187252 119446 318859 119448
rect 187252 119444 187258 119446
rect 318793 119443 318859 119446
rect 203742 119308 203748 119372
rect 203812 119370 203818 119372
rect 536833 119370 536899 119373
rect 203812 119368 536899 119370
rect 203812 119312 536838 119368
rect 536894 119312 536899 119368
rect 203812 119310 536899 119312
rect 203812 119308 203818 119310
rect 536833 119307 536899 119310
rect 196934 117948 196940 118012
rect 197004 118010 197010 118012
rect 447777 118010 447843 118013
rect 197004 118008 447843 118010
rect 197004 117952 447782 118008
rect 447838 117952 447843 118008
rect 197004 117950 447843 117952
rect 197004 117948 197010 117950
rect 447777 117947 447843 117950
rect 189758 115228 189764 115292
rect 189828 115290 189834 115292
rect 343633 115290 343699 115293
rect 189828 115288 343699 115290
rect 189828 115232 343638 115288
rect 343694 115232 343699 115288
rect 189828 115230 343699 115232
rect 189828 115228 189834 115230
rect 343633 115227 343699 115230
rect 198038 115092 198044 115156
rect 198108 115154 198114 115156
rect 465073 115154 465139 115157
rect 198108 115152 465139 115154
rect 198108 115096 465078 115152
rect 465134 115096 465139 115152
rect 198108 115094 465139 115096
rect 198108 115092 198114 115094
rect 465073 115091 465139 115094
rect 188286 113868 188292 113932
rect 188356 113930 188362 113932
rect 315297 113930 315363 113933
rect 188356 113928 315363 113930
rect 188356 113872 315302 113928
rect 315358 113872 315363 113928
rect 188356 113870 315363 113872
rect 188356 113868 188362 113870
rect 315297 113867 315363 113870
rect 44817 113794 44883 113797
rect 165838 113794 165844 113796
rect 44817 113792 165844 113794
rect 44817 113736 44822 113792
rect 44878 113736 165844 113792
rect 44817 113734 165844 113736
rect 44817 113731 44883 113734
rect 165838 113732 165844 113734
rect 165908 113732 165914 113796
rect 199694 113732 199700 113796
rect 199764 113794 199770 113796
rect 476113 113794 476179 113797
rect 199764 113792 476179 113794
rect 199764 113736 476118 113792
rect 476174 113736 476179 113792
rect 199764 113734 476179 113736
rect 199764 113732 199770 113734
rect 476113 113731 476179 113734
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 44173 112434 44239 112437
rect 166022 112434 166028 112436
rect 44173 112432 166028 112434
rect 44173 112376 44178 112432
rect 44234 112376 166028 112432
rect 44173 112374 166028 112376
rect 44173 112371 44239 112374
rect 166022 112372 166028 112374
rect 166092 112372 166098 112436
rect 181478 112372 181484 112436
rect 181548 112434 181554 112436
rect 247677 112434 247743 112437
rect 181548 112432 247743 112434
rect 181548 112376 247682 112432
rect 247738 112376 247743 112432
rect 181548 112374 247743 112376
rect 181548 112372 181554 112374
rect 247677 112371 247743 112374
rect 331806 111828 331812 111892
rect 331876 111890 331882 111892
rect 583526 111890 583586 112646
rect 331876 111830 583586 111890
rect 331876 111828 331882 111830
rect 129733 111074 129799 111077
rect 173014 111074 173020 111076
rect 129733 111072 173020 111074
rect 129733 111016 129738 111072
rect 129794 111016 173020 111072
rect 129733 111014 173020 111016
rect 129733 111011 129799 111014
rect 173014 111012 173020 111014
rect 173084 111012 173090 111076
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 200982 109652 200988 109716
rect 201052 109714 201058 109716
rect 485773 109714 485839 109717
rect 201052 109712 485839 109714
rect 201052 109656 485778 109712
rect 485834 109656 485839 109712
rect 201052 109654 485839 109656
rect 201052 109652 201058 109654
rect 485773 109651 485839 109654
rect 200798 106796 200804 106860
rect 200868 106858 200874 106860
rect 496813 106858 496879 106861
rect 200868 106856 496879 106858
rect 200868 106800 496818 106856
rect 496874 106800 496879 106856
rect 200868 106798 496879 106800
rect 200868 106796 200874 106798
rect 496813 106795 496879 106798
rect 187366 105436 187372 105500
rect 187436 105498 187442 105500
rect 311157 105498 311223 105501
rect 187436 105496 311223 105498
rect 187436 105440 311162 105496
rect 311218 105440 311223 105496
rect 187436 105438 311223 105440
rect 187436 105436 187442 105438
rect 311157 105435 311223 105438
rect 202270 104076 202276 104140
rect 202340 104138 202346 104140
rect 506565 104138 506631 104141
rect 202340 104136 506631 104138
rect 202340 104080 506570 104136
rect 506626 104080 506631 104136
rect 202340 104078 506631 104080
rect 202340 104076 202346 104078
rect 506565 104075 506631 104078
rect 188470 102716 188476 102780
rect 188540 102778 188546 102780
rect 332685 102778 332751 102781
rect 188540 102776 332751 102778
rect 188540 102720 332690 102776
rect 332746 102720 332751 102776
rect 188540 102718 332751 102720
rect 188540 102716 188546 102718
rect 332685 102715 332751 102718
rect 202454 101356 202460 101420
rect 202524 101418 202530 101420
rect 514845 101418 514911 101421
rect 202524 101416 514911 101418
rect 202524 101360 514850 101416
rect 514906 101360 514911 101416
rect 202524 101358 514911 101360
rect 202524 101356 202530 101358
rect 514845 101355 514911 101358
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 181294 98772 181300 98836
rect 181364 98834 181370 98836
rect 251265 98834 251331 98837
rect 181364 98832 251331 98834
rect 181364 98776 251270 98832
rect 251326 98776 251331 98832
rect 181364 98774 251331 98776
rect 181364 98772 181370 98774
rect 251265 98771 251331 98774
rect 198222 98636 198228 98700
rect 198292 98698 198298 98700
rect 454033 98698 454099 98701
rect 198292 98696 454099 98698
rect 198292 98640 454038 98696
rect 454094 98640 454099 98696
rect 198292 98638 454099 98640
rect 198292 98636 198298 98638
rect 454033 98635 454099 98638
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 203926 95780 203932 95844
rect 203996 95842 204002 95844
rect 531405 95842 531471 95845
rect 203996 95840 531471 95842
rect 203996 95784 531410 95840
rect 531466 95784 531471 95840
rect 203996 95782 531471 95784
rect 203996 95780 204002 95782
rect 531405 95779 531471 95782
rect 179086 91700 179092 91764
rect 179156 91762 179162 91764
rect 204253 91762 204319 91765
rect 179156 91760 204319 91762
rect 179156 91704 204258 91760
rect 204314 91704 204319 91760
rect 179156 91702 204319 91704
rect 179156 91700 179162 91702
rect 204253 91699 204319 91702
rect 205214 90340 205220 90404
rect 205284 90402 205290 90404
rect 548517 90402 548583 90405
rect 205284 90400 548583 90402
rect 205284 90344 548522 90400
rect 548578 90344 548583 90400
rect 205284 90342 548583 90344
rect 205284 90340 205290 90342
rect 548517 90339 548583 90342
rect 580257 86186 580323 86189
rect 583520 86186 584960 86276
rect 580257 86184 584960 86186
rect 580257 86128 580262 86184
rect 580318 86128 584960 86184
rect 580257 86126 584960 86128
rect 580257 86123 580323 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 205766 84764 205772 84828
rect 205836 84826 205842 84828
rect 564433 84826 564499 84829
rect 205836 84824 564499 84826
rect 205836 84768 564438 84824
rect 564494 84768 564499 84824
rect 205836 84766 564499 84768
rect 205836 84764 205842 84766
rect 564433 84763 564499 84766
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 280654 71844 280660 71908
rect 280724 71906 280730 71908
rect 583526 71906 583586 72798
rect 280724 71846 583586 71906
rect 280724 71844 280730 71846
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 202638 71028 202644 71092
rect 202708 71090 202714 71092
rect 517513 71090 517579 71093
rect 202708 71088 517579 71090
rect 202708 71032 517518 71088
rect 517574 71032 517579 71088
rect 202708 71030 517579 71032
rect 202708 71028 202714 71030
rect 517513 71027 517579 71030
rect 204110 69532 204116 69596
rect 204180 69594 204186 69596
rect 528553 69594 528619 69597
rect 204180 69592 528619 69594
rect 204180 69536 528558 69592
rect 528614 69536 528619 69592
rect 204180 69534 528619 69536
rect 204180 69532 204186 69534
rect 528553 69531 528619 69534
rect 187550 68172 187556 68236
rect 187620 68234 187626 68236
rect 322933 68234 322999 68237
rect 187620 68232 322999 68234
rect 187620 68176 322938 68232
rect 322994 68176 322999 68232
rect 187620 68174 322999 68176
rect 187620 68172 187626 68174
rect 322933 68171 322999 68174
rect 188654 66812 188660 66876
rect 188724 66874 188730 66876
rect 336733 66874 336799 66877
rect 188724 66872 336799 66874
rect 188724 66816 336738 66872
rect 336794 66816 336799 66872
rect 188724 66814 336799 66816
rect 188724 66812 188730 66814
rect 336733 66811 336799 66814
rect 188838 65452 188844 65516
rect 188908 65514 188914 65516
rect 340965 65514 341031 65517
rect 188908 65512 341031 65514
rect 188908 65456 340970 65512
rect 341026 65456 341031 65512
rect 188908 65454 341031 65456
rect 188908 65452 188914 65454
rect 340965 65451 341031 65454
rect 190126 64092 190132 64156
rect 190196 64154 190202 64156
rect 350533 64154 350599 64157
rect 190196 64152 350599 64154
rect 190196 64096 350538 64152
rect 350594 64096 350599 64152
rect 190196 64094 350599 64096
rect 190196 64092 190202 64094
rect 350533 64091 350599 64094
rect 189942 62732 189948 62796
rect 190012 62794 190018 62796
rect 354673 62794 354739 62797
rect 190012 62792 354739 62794
rect 190012 62736 354678 62792
rect 354734 62736 354739 62792
rect 190012 62734 354739 62736
rect 190012 62732 190018 62734
rect 354673 62731 354739 62734
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 335854 59332 335860 59396
rect 335924 59394 335930 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 335924 59334 567210 59394
rect 335924 59332 335930 59334
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 194174 54436 194180 54500
rect 194244 54498 194250 54500
rect 407205 54498 407271 54501
rect 194244 54496 407271 54498
rect 194244 54440 407210 54496
rect 407266 54440 407271 54496
rect 194244 54438 407271 54440
rect 194244 54436 194250 54438
rect 407205 54435 407271 54438
rect 194358 51716 194364 51780
rect 194428 51778 194434 51780
rect 411253 51778 411319 51781
rect 194428 51776 411319 51778
rect 194428 51720 411258 51776
rect 411314 51720 411319 51776
rect 194428 51718 411319 51720
rect 194428 51716 194434 51718
rect 411253 51715 411319 51718
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 197854 46140 197860 46204
rect 197924 46202 197930 46204
rect 456885 46202 456951 46205
rect 197924 46200 456951 46202
rect 197924 46144 456890 46200
rect 456946 46144 456951 46200
rect 583520 46188 584960 46278
rect 197924 46142 456951 46144
rect 197924 46140 197930 46142
rect 456885 46139 456951 46142
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 198406 44780 198412 44844
rect 198476 44842 198482 44844
rect 460933 44842 460999 44845
rect 198476 44840 460999 44842
rect 198476 44784 460938 44840
rect 460994 44784 460999 44840
rect 198476 44782 460999 44784
rect 198476 44780 198482 44782
rect 460933 44779 460999 44782
rect 199878 42060 199884 42124
rect 199948 42122 199954 42124
rect 474733 42122 474799 42125
rect 199948 42120 474799 42122
rect 199948 42064 474738 42120
rect 474794 42064 474799 42120
rect 199948 42062 474799 42064
rect 199948 42060 199954 42062
rect 474733 42059 474799 42062
rect 190310 40564 190316 40628
rect 190380 40626 190386 40628
rect 357525 40626 357591 40629
rect 190380 40624 357591 40626
rect 190380 40568 357530 40624
rect 357586 40568 357591 40624
rect 190380 40566 357591 40568
rect 190380 40564 190386 40566
rect 357525 40563 357591 40566
rect 201166 37844 201172 37908
rect 201236 37906 201242 37908
rect 487153 37906 487219 37909
rect 201236 37904 487219 37906
rect 201236 37848 487158 37904
rect 487214 37848 487219 37904
rect 201236 37846 487219 37848
rect 201236 37844 201242 37846
rect 487153 37843 487219 37846
rect 205398 35124 205404 35188
rect 205468 35186 205474 35188
rect 547965 35186 548031 35189
rect 205468 35184 548031 35186
rect 205468 35128 547970 35184
rect 548026 35128 548031 35184
rect 205468 35126 548031 35128
rect 205468 35124 205474 35126
rect 547965 35123 548031 35126
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 195462 30908 195468 30972
rect 195532 30970 195538 30972
rect 430573 30970 430639 30973
rect 195532 30968 430639 30970
rect 195532 30912 430578 30968
rect 430634 30912 430639 30968
rect 195532 30910 430639 30912
rect 195532 30908 195538 30910
rect 430573 30907 430639 30910
rect 177246 24108 177252 24172
rect 177316 24170 177322 24172
rect 197997 24170 198063 24173
rect 177316 24168 198063 24170
rect 177316 24112 198002 24168
rect 198058 24112 198063 24168
rect 177316 24110 198063 24112
rect 177316 24108 177322 24110
rect 197997 24107 198063 24110
rect 580073 19818 580139 19821
rect 583520 19818 584960 19908
rect 580073 19816 584960 19818
rect 580073 19760 580078 19816
rect 580134 19760 584960 19816
rect 580073 19758 584960 19760
rect 580073 19755 580139 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 201350 18532 201356 18596
rect 201420 18594 201426 18596
rect 490005 18594 490071 18597
rect 201420 18592 490071 18594
rect 201420 18536 490010 18592
rect 490066 18536 490071 18592
rect 201420 18534 490071 18536
rect 201420 18532 201426 18534
rect 490005 18531 490071 18534
rect 197118 11596 197124 11660
rect 197188 11658 197194 11660
rect 440325 11658 440391 11661
rect 197188 11656 440391 11658
rect 197188 11600 440330 11656
rect 440386 11600 440391 11656
rect 197188 11598 440391 11600
rect 197188 11596 197194 11598
rect 440325 11595 440391 11598
rect 192702 9420 192708 9484
rect 192772 9482 192778 9484
rect 379973 9482 380039 9485
rect 192772 9480 380039 9482
rect 192772 9424 379978 9480
rect 380034 9424 380039 9480
rect 192772 9422 380039 9424
rect 192772 9420 192778 9422
rect 379973 9419 380039 9422
rect 192886 9284 192892 9348
rect 192956 9346 192962 9348
rect 387149 9346 387215 9349
rect 192956 9344 387215 9346
rect 192956 9288 387154 9344
rect 387210 9288 387215 9344
rect 192956 9286 387215 9288
rect 192956 9284 192962 9286
rect 387149 9283 387215 9286
rect 192518 9148 192524 9212
rect 192588 9210 192594 9212
rect 394233 9210 394299 9213
rect 192588 9208 394299 9210
rect 192588 9152 394238 9208
rect 394294 9152 394299 9208
rect 192588 9150 394299 9152
rect 192588 9148 192594 9150
rect 394233 9147 394299 9150
rect 195646 9012 195652 9076
rect 195716 9074 195722 9076
rect 415485 9074 415551 9077
rect 195716 9072 415551 9074
rect 195716 9016 415490 9072
rect 415546 9016 415551 9072
rect 195716 9014 415551 9016
rect 195716 9012 195722 9014
rect 415485 9011 415551 9014
rect 195094 8876 195100 8940
rect 195164 8938 195170 8940
rect 422569 8938 422635 8941
rect 195164 8936 422635 8938
rect 195164 8880 422574 8936
rect 422630 8880 422635 8936
rect 195164 8878 422635 8880
rect 195164 8876 195170 8878
rect 422569 8875 422635 8878
rect 205950 7516 205956 7580
rect 206020 7578 206026 7580
rect 571517 7578 571583 7581
rect 206020 7576 571583 7578
rect 206020 7520 571522 7576
rect 571578 7520 571583 7576
rect 206020 7518 571583 7520
rect 206020 7516 206026 7518
rect 571517 7515 571583 7518
rect 184606 6836 184612 6900
rect 184676 6898 184682 6900
rect 284293 6898 284359 6901
rect 184676 6896 284359 6898
rect 184676 6840 284298 6896
rect 284354 6840 284359 6896
rect 184676 6838 284359 6840
rect 184676 6836 184682 6838
rect 284293 6835 284359 6838
rect 184974 6700 184980 6764
rect 185044 6762 185050 6764
rect 291377 6762 291443 6765
rect 185044 6760 291443 6762
rect 185044 6704 291382 6760
rect 291438 6704 291443 6760
rect 185044 6702 291443 6704
rect 185044 6700 185050 6702
rect 291377 6699 291443 6702
rect -960 6490 480 6580
rect 185158 6564 185164 6628
rect 185228 6626 185234 6628
rect 294873 6626 294939 6629
rect 185228 6624 294939 6626
rect 185228 6568 294878 6624
rect 294934 6568 294939 6624
rect 185228 6566 294939 6568
rect 185228 6564 185234 6566
rect 294873 6563 294939 6566
rect 580349 6626 580415 6629
rect 583520 6626 584960 6716
rect 580349 6624 584960 6626
rect 580349 6568 580354 6624
rect 580410 6568 584960 6624
rect 580349 6566 584960 6568
rect 580349 6563 580415 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 191598 6428 191604 6492
rect 191668 6490 191674 6492
rect 365805 6490 365871 6493
rect 191668 6488 365871 6490
rect 191668 6432 365810 6488
rect 365866 6432 365871 6488
rect 583520 6476 584960 6566
rect 191668 6430 365871 6432
rect 191668 6428 191674 6430
rect 365805 6427 365871 6430
rect 191414 6292 191420 6356
rect 191484 6354 191490 6356
rect 376477 6354 376543 6357
rect 191484 6352 376543 6354
rect 191484 6296 376482 6352
rect 376538 6296 376543 6352
rect 191484 6294 376543 6296
rect 191484 6292 191490 6294
rect 376477 6291 376543 6294
rect 193070 6156 193076 6220
rect 193140 6218 193146 6220
rect 390645 6218 390711 6221
rect 193140 6216 390711 6218
rect 193140 6160 390650 6216
rect 390706 6160 390711 6216
rect 193140 6158 390711 6160
rect 193140 6156 193146 6158
rect 390645 6155 390711 6158
rect 184422 6020 184428 6084
rect 184492 6082 184498 6084
rect 280705 6082 280771 6085
rect 184492 6080 280771 6082
rect 184492 6024 280710 6080
rect 280766 6024 280771 6080
rect 184492 6022 280771 6024
rect 184492 6020 184498 6022
rect 280705 6019 280771 6022
rect 179270 3572 179276 3636
rect 179340 3634 179346 3636
rect 203885 3634 203951 3637
rect 179340 3632 203951 3634
rect 179340 3576 203890 3632
rect 203946 3576 203951 3632
rect 179340 3574 203951 3576
rect 179340 3572 179346 3574
rect 203885 3571 203951 3574
rect 184238 3436 184244 3500
rect 184308 3498 184314 3500
rect 273621 3498 273687 3501
rect 184308 3496 273687 3498
rect 184308 3440 273626 3496
rect 273682 3440 273687 3496
rect 184308 3438 273687 3440
rect 184308 3436 184314 3438
rect 273621 3435 273687 3438
rect 184054 3300 184060 3364
rect 184124 3362 184130 3364
rect 277117 3362 277183 3365
rect 184124 3360 277183 3362
rect 184124 3304 277122 3360
rect 277178 3304 277183 3360
rect 184124 3302 277183 3304
rect 184124 3300 184130 3302
rect 277117 3299 277183 3302
<< via3 >>
rect 374132 452508 374196 452572
rect 278636 451828 278700 451892
rect 343956 451556 344020 451620
rect 355180 451284 355244 451348
rect 362908 451284 362972 451348
rect 368244 451284 368308 451348
rect 376892 451284 376956 451348
rect 360332 449984 360396 449988
rect 360332 449928 360382 449984
rect 360382 449928 360396 449984
rect 360332 449924 360396 449928
rect 363276 449924 363340 449988
rect 364380 449924 364444 449988
rect 360516 449788 360580 449852
rect 374132 449516 374196 449580
rect 343772 449440 343836 449444
rect 343772 449384 343822 449440
rect 343822 449384 343836 449440
rect 343772 449380 343836 449384
rect 345796 449440 345860 449444
rect 345796 449384 345800 449440
rect 345800 449384 345856 449440
rect 345856 449384 345860 449440
rect 345796 449380 345860 449384
rect 347452 449380 347516 449444
rect 370452 449380 370516 449444
rect 373212 449440 373276 449444
rect 373212 449384 373226 449440
rect 373226 449384 373276 449440
rect 373212 449380 373276 449384
rect 374316 449440 374380 449444
rect 374316 449384 374330 449440
rect 374330 449384 374380 449440
rect 374316 449380 374380 449384
rect 384988 449380 385052 449444
rect 347636 449304 347700 449308
rect 347636 449248 347640 449304
rect 347640 449248 347696 449304
rect 347696 449248 347700 449304
rect 347636 449244 347700 449248
rect 371188 449304 371252 449308
rect 371188 449248 371192 449304
rect 371192 449248 371248 449304
rect 371248 449248 371252 449304
rect 371188 449244 371252 449248
rect 382228 449304 382292 449308
rect 382228 449248 382232 449304
rect 382232 449248 382288 449304
rect 382288 449248 382292 449304
rect 382228 449244 382292 449248
rect 383700 449304 383764 449308
rect 383700 449248 383704 449304
rect 383704 449248 383760 449304
rect 383760 449248 383764 449304
rect 383700 449244 383764 449248
rect 347636 448564 347700 448628
rect 347452 447884 347516 447948
rect 345796 447748 345860 447812
rect 360148 447476 360212 447540
rect 360516 447476 360580 447540
rect 343956 443532 344020 443596
rect 307708 404288 307772 404292
rect 307708 404232 307722 404288
rect 307722 404232 307772 404288
rect 307708 404228 307772 404232
rect 343956 402188 344020 402252
rect 343036 402052 343100 402116
rect 360148 401916 360212 401980
rect 360516 401916 360580 401980
rect 347636 401644 347700 401708
rect 371188 401508 371252 401572
rect 355180 401236 355244 401300
rect 362908 401100 362972 401164
rect 360332 400964 360396 401028
rect 374316 400828 374380 400892
rect 352420 400692 352484 400756
rect 355364 400556 355428 400620
rect 343772 400420 343836 400484
rect 345796 400284 345860 400348
rect 354076 400284 354140 400348
rect 355548 400148 355612 400212
rect 357388 400148 357452 400212
rect 370452 400148 370516 400212
rect 354444 400012 354508 400076
rect 354628 400012 354692 400076
rect 343036 399936 343100 399940
rect 343036 399880 343040 399936
rect 343040 399880 343096 399936
rect 343096 399880 343100 399936
rect 343036 399876 343100 399880
rect 343772 399936 343836 399940
rect 343772 399880 343776 399936
rect 343776 399880 343832 399936
rect 343832 399880 343836 399936
rect 343772 399876 343836 399880
rect 344692 399936 344756 399940
rect 344692 399880 344696 399936
rect 344696 399880 344752 399936
rect 344752 399880 344756 399936
rect 344692 399876 344756 399880
rect 345060 399936 345124 399940
rect 345060 399880 345064 399936
rect 345064 399880 345120 399936
rect 345120 399880 345124 399936
rect 345060 399876 345124 399880
rect 345428 399876 345492 399940
rect 345796 399876 345860 399940
rect 347268 399936 347332 399940
rect 347268 399880 347272 399936
rect 347272 399880 347328 399936
rect 347328 399880 347332 399936
rect 342300 399740 342364 399804
rect 343220 399800 343284 399804
rect 343220 399744 343224 399800
rect 343224 399744 343280 399800
rect 343280 399744 343284 399800
rect 343220 399740 343284 399744
rect 345244 399740 345308 399804
rect 347268 399876 347332 399880
rect 347636 399876 347700 399940
rect 348004 399936 348068 399940
rect 348004 399880 348008 399936
rect 348008 399880 348064 399936
rect 348064 399880 348068 399936
rect 348004 399876 348068 399880
rect 348372 399936 348436 399940
rect 348372 399880 348376 399936
rect 348376 399880 348432 399936
rect 348432 399880 348436 399936
rect 348372 399876 348436 399880
rect 348556 399876 348620 399940
rect 350396 399936 350460 399940
rect 350396 399880 350400 399936
rect 350400 399880 350456 399936
rect 350456 399880 350460 399936
rect 350396 399876 350460 399880
rect 350580 399876 350644 399940
rect 346348 399740 346412 399804
rect 350028 399800 350092 399804
rect 350028 399744 350032 399800
rect 350032 399744 350088 399800
rect 350088 399744 350092 399800
rect 350028 399740 350092 399744
rect 351684 399740 351748 399804
rect 352236 399876 352300 399940
rect 353708 399876 353772 399940
rect 354628 399876 354692 399940
rect 355180 400012 355244 400076
rect 364380 400012 364444 400076
rect 355548 399876 355612 399940
rect 374132 400012 374196 400076
rect 366588 399876 366652 399940
rect 366772 399936 366836 399940
rect 366772 399880 366776 399936
rect 366776 399880 366832 399936
rect 366832 399880 366836 399936
rect 366772 399876 366836 399880
rect 368060 399936 368124 399940
rect 368060 399880 368064 399936
rect 368064 399880 368120 399936
rect 368120 399880 368124 399936
rect 368060 399876 368124 399880
rect 368428 399876 368492 399940
rect 369716 399936 369780 399940
rect 369716 399880 369720 399936
rect 369720 399880 369776 399936
rect 369776 399880 369780 399936
rect 369716 399876 369780 399880
rect 371004 399936 371068 399940
rect 371004 399880 371008 399936
rect 371008 399880 371064 399936
rect 371064 399880 371068 399936
rect 371004 399876 371068 399880
rect 371188 399876 371252 399940
rect 352420 399800 352484 399804
rect 352420 399744 352470 399800
rect 352470 399744 352484 399800
rect 352420 399740 352484 399744
rect 353156 399740 353220 399804
rect 354076 399740 354140 399804
rect 360516 399740 360580 399804
rect 360884 399740 360948 399804
rect 362540 399800 362604 399804
rect 362540 399744 362544 399800
rect 362544 399744 362600 399800
rect 362600 399744 362604 399800
rect 355180 399604 355244 399668
rect 355364 399664 355428 399668
rect 355364 399608 355414 399664
rect 355414 399608 355428 399664
rect 355364 399604 355428 399608
rect 355548 399604 355612 399668
rect 358676 399604 358740 399668
rect 360700 399604 360764 399668
rect 362540 399740 362604 399744
rect 363092 399740 363156 399804
rect 364196 399740 364260 399804
rect 371740 399936 371804 399940
rect 371740 399880 371744 399936
rect 371744 399880 371800 399936
rect 371800 399880 371804 399936
rect 371740 399876 371804 399880
rect 366588 399740 366652 399804
rect 367508 399740 367572 399804
rect 369900 399740 369964 399804
rect 366220 399604 366284 399668
rect 368244 399604 368308 399668
rect 343956 399332 344020 399396
rect 357388 399392 357452 399396
rect 357388 399336 357402 399392
rect 357402 399336 357452 399392
rect 357388 399332 357452 399336
rect 370452 399468 370516 399532
rect 371556 399740 371620 399804
rect 372844 399740 372908 399804
rect 374316 399876 374380 399940
rect 372292 399604 372356 399668
rect 374868 399800 374932 399804
rect 374868 399744 374872 399800
rect 374872 399744 374928 399800
rect 374928 399744 374932 399800
rect 374868 399740 374932 399744
rect 377628 399936 377692 399940
rect 377628 399880 377632 399936
rect 377632 399880 377688 399936
rect 377688 399880 377692 399936
rect 377628 399876 377692 399880
rect 378364 400148 378428 400212
rect 379284 400012 379348 400076
rect 379100 399876 379164 399940
rect 378180 399740 378244 399804
rect 381676 400012 381740 400076
rect 382412 399876 382476 399940
rect 378548 399528 378612 399532
rect 378548 399472 378598 399528
rect 378598 399472 378612 399528
rect 378548 399468 378612 399472
rect 379836 399740 379900 399804
rect 382228 399332 382292 399396
rect 289124 398924 289188 398988
rect 349108 399196 349172 399260
rect 353340 399196 353404 399260
rect 310284 398788 310348 398852
rect 358124 399196 358188 399260
rect 373212 399196 373276 399260
rect 373948 399196 374012 399260
rect 368428 399060 368492 399124
rect 371740 399060 371804 399124
rect 371740 398924 371804 398988
rect 365116 398652 365180 398716
rect 371004 398652 371068 398716
rect 350764 398516 350828 398580
rect 352420 398244 352484 398308
rect 343220 398108 343284 398172
rect 348004 398108 348068 398172
rect 357572 398108 357636 398172
rect 355180 397972 355244 398036
rect 368980 397972 369044 398036
rect 357388 397836 357452 397900
rect 375972 397836 376036 397900
rect 360332 397700 360396 397764
rect 377260 397700 377324 397764
rect 372292 397624 372356 397628
rect 372292 397568 372306 397624
rect 372306 397568 372356 397624
rect 372292 397564 372356 397568
rect 380940 397564 381004 397628
rect 382228 397564 382292 397628
rect 350396 397428 350460 397492
rect 353156 397428 353220 397492
rect 356468 397488 356532 397492
rect 356468 397432 356518 397488
rect 356518 397432 356532 397488
rect 356468 397428 356532 397432
rect 358124 397428 358188 397492
rect 359412 397428 359476 397492
rect 372844 397428 372908 397492
rect 382044 397428 382108 397492
rect 364380 397292 364444 397356
rect 367876 397352 367940 397356
rect 367876 397296 367926 397352
rect 367926 397296 367940 397352
rect 367876 397292 367940 397296
rect 369164 397292 369228 397356
rect 375420 397292 375484 397356
rect 382412 397352 382476 397356
rect 382412 397296 382462 397352
rect 382462 397296 382476 397352
rect 382412 397292 382476 397296
rect 382780 397292 382844 397356
rect 283420 397156 283484 397220
rect 358124 397156 358188 397220
rect 372292 397216 372356 397220
rect 372292 397160 372342 397216
rect 372342 397160 372356 397216
rect 372292 397156 372356 397160
rect 355548 397020 355612 397084
rect 357020 397020 357084 397084
rect 374316 397020 374380 397084
rect 358860 396944 358924 396948
rect 358860 396888 358910 396944
rect 358910 396888 358924 396944
rect 358860 396884 358924 396888
rect 362908 396884 362972 396948
rect 356652 396748 356716 396812
rect 378180 396748 378244 396812
rect 355180 396476 355244 396540
rect 357388 396612 357452 396676
rect 358308 396612 358372 396676
rect 378180 396612 378244 396676
rect 379836 396612 379900 396676
rect 363460 396476 363524 396540
rect 377628 396476 377692 396540
rect 354260 396204 354324 396268
rect 354812 395932 354876 395996
rect 342300 395524 342364 395588
rect 368612 395524 368676 395588
rect 373764 395388 373828 395452
rect 374132 395388 374196 395452
rect 354628 395252 354692 395316
rect 356836 395252 356900 395316
rect 379652 395252 379716 395316
rect 368428 395176 368492 395180
rect 368428 395120 368442 395176
rect 368442 395120 368492 395176
rect 368428 395116 368492 395120
rect 379100 395116 379164 395180
rect 345428 394708 345492 394772
rect 297220 394572 297284 394636
rect 372292 394572 372356 394636
rect 297956 394436 298020 394500
rect 357572 394436 357636 394500
rect 296484 394300 296548 394364
rect 321324 394164 321388 394228
rect 372660 393892 372724 393956
rect 350028 393484 350092 393548
rect 357940 393484 358004 393548
rect 378364 393484 378428 393548
rect 344692 393348 344756 393412
rect 347820 393348 347884 393412
rect 349292 393408 349356 393412
rect 349292 393352 349342 393408
rect 349342 393352 349356 393408
rect 349292 393348 349356 393352
rect 362540 393348 362604 393412
rect 369716 393348 369780 393412
rect 299244 393212 299308 393276
rect 360884 393212 360948 393276
rect 364932 393212 364996 393276
rect 367876 393212 367940 393276
rect 306236 393076 306300 393140
rect 364196 393076 364260 393140
rect 366772 393076 366836 393140
rect 367692 393076 367756 393140
rect 304764 392940 304828 393004
rect 366220 392940 366284 393004
rect 300716 392804 300780 392868
rect 368060 392804 368124 392868
rect 304580 392668 304644 392732
rect 293172 392532 293236 392596
rect 352236 392532 352300 392596
rect 358676 392532 358740 392596
rect 303476 392396 303540 392460
rect 282868 392048 282932 392052
rect 282868 391992 282918 392048
rect 282918 391992 282932 392048
rect 282868 391988 282932 391992
rect 341012 391988 341076 392052
rect 311756 391716 311820 391780
rect 371188 391716 371252 391780
rect 295012 391580 295076 391644
rect 353708 391580 353772 391644
rect 295196 391036 295260 391100
rect 314148 390900 314212 390964
rect 294644 390492 294708 390556
rect 317276 390356 317340 390420
rect 345060 389812 345124 389876
rect 316724 389676 316788 389740
rect 378548 389268 378612 389332
rect 373948 389192 374012 389196
rect 373948 389136 373962 389192
rect 373962 389136 374012 389192
rect 373948 389132 374012 389136
rect 291700 388996 291764 389060
rect 288020 388860 288084 388924
rect 287468 388724 287532 388788
rect 348372 388724 348436 388788
rect 289492 388588 289556 388652
rect 348556 388588 348620 388652
rect 344876 388452 344940 388516
rect 383700 388452 383764 388516
rect 345244 388316 345308 388380
rect 384988 388316 385052 388380
rect 286732 388180 286796 388244
rect 307524 387636 307588 387700
rect 366588 387636 366652 387700
rect 287836 387500 287900 387564
rect 297588 387364 297652 387428
rect 281396 387092 281460 387156
rect 357020 387092 357084 387156
rect 347268 386956 347332 387020
rect 302004 385868 302068 385932
rect 376892 385732 376956 385796
rect 360332 385596 360396 385660
rect 298876 384372 298940 384436
rect 363276 384236 363340 384300
rect 373948 383828 374012 383892
rect 373948 383420 374012 383484
rect 366404 382060 366468 382124
rect 364380 381924 364444 381988
rect 371740 381788 371804 381852
rect 286364 381652 286428 381716
rect 368612 381652 368676 381716
rect 292988 381516 293052 381580
rect 291884 379340 291948 379404
rect 290964 379204 291028 379268
rect 291332 379068 291396 379132
rect 292252 378932 292316 378996
rect 290780 378796 290844 378860
rect 288756 378660 288820 378724
rect 289308 378524 289372 378588
rect 354812 377980 354876 378044
rect 353340 377844 353404 377908
rect 308996 377436 309060 377500
rect 314700 377300 314764 377364
rect 285076 376756 285140 376820
rect 296300 375940 296364 376004
rect 279372 375396 279436 375460
rect 292804 374716 292868 374780
rect 297404 374580 297468 374644
rect 373948 374096 374012 374100
rect 373948 374040 373962 374096
rect 373962 374040 374012 374096
rect 373948 374036 374012 374040
rect 373948 373764 374012 373828
rect 220676 373356 220740 373420
rect 280476 372948 280540 373012
rect 279924 372676 279988 372740
rect 280660 372268 280724 372332
rect 277900 372132 277964 372196
rect 276612 371996 276676 372060
rect 314332 371860 314396 371924
rect 372660 371860 372724 371924
rect 279556 371452 279620 371516
rect 307708 371452 307772 371516
rect 282684 371316 282748 371380
rect 323164 371316 323228 371380
rect 316908 370500 316972 370564
rect 285260 369820 285324 369884
rect 312492 370092 312556 370156
rect 315620 369820 315684 369884
rect 319668 369820 319732 369884
rect 331812 369956 331876 370020
rect 335860 369820 335924 369884
rect 282132 369684 282196 369748
rect 319300 369548 319364 369612
rect 281580 369412 281644 369476
rect 282684 369412 282748 369476
rect 286548 369412 286612 369476
rect 287284 369472 287348 369476
rect 287284 369416 287288 369472
rect 287288 369416 287344 369472
rect 287344 369416 287348 369472
rect 287284 369412 287348 369416
rect 304948 369412 305012 369476
rect 306972 369412 307036 369476
rect 311020 369412 311084 369476
rect 313780 369412 313844 369476
rect 318012 369412 318076 369476
rect 319852 369472 319916 369476
rect 319852 369416 319902 369472
rect 319902 369416 319916 369472
rect 319852 369412 319916 369416
rect 320772 369412 320836 369476
rect 322060 369412 322124 369476
rect 278636 369276 278700 369340
rect 288940 369276 289004 369340
rect 315436 369004 315500 369068
rect 278636 368596 278700 368660
rect 285260 368732 285324 368796
rect 288940 368596 289004 368660
rect 287284 368460 287348 368524
rect 307708 367644 307772 367708
rect 321140 367644 321204 367708
rect 379652 367644 379716 367708
rect 280476 366284 280540 366348
rect 323164 366284 323228 366348
rect 373948 364440 374012 364444
rect 373948 364384 373962 364440
rect 373962 364384 374012 364440
rect 373948 364380 374012 364384
rect 373948 364108 374012 364172
rect 281580 361796 281644 361860
rect 280660 360980 280724 361044
rect 282132 360844 282196 360908
rect 279924 359348 279988 359412
rect 280660 359348 280724 359412
rect 373948 354784 374012 354788
rect 373948 354728 373962 354784
rect 373962 354728 374012 354784
rect 373948 354724 374012 354728
rect 373948 354452 374012 354516
rect 325372 345612 325436 345676
rect 381676 345612 381740 345676
rect 373948 345128 374012 345132
rect 373948 345072 373962 345128
rect 373962 345072 374012 345128
rect 373948 345068 374012 345072
rect 373948 344992 374012 344996
rect 373948 344936 373962 344992
rect 373962 344936 374012 344992
rect 373948 344932 374012 344936
rect 324268 342892 324332 342956
rect 382780 342892 382844 342956
rect 373948 340776 374012 340780
rect 373948 340720 373962 340776
rect 373962 340720 374012 340776
rect 373948 340716 374012 340720
rect 379284 337316 379348 337380
rect 373948 331256 374012 331260
rect 373948 331200 373962 331256
rect 373962 331200 374012 331256
rect 373948 331196 374012 331200
rect 276612 330380 276676 330444
rect 382044 329836 382108 329900
rect 368428 329292 368492 329356
rect 326844 328476 326908 328540
rect 338252 329020 338316 329084
rect 375236 328476 375300 328540
rect 375236 327660 375300 327724
rect 378180 326572 378244 326636
rect 374132 326436 374196 326500
rect 327580 326300 327644 326364
rect 373948 325892 374012 325956
rect 323348 325756 323412 325820
rect 371372 325348 371436 325412
rect 374132 325212 374196 325276
rect 330340 325076 330404 325140
rect 323532 324940 323596 325004
rect 382228 324940 382292 325004
rect 327764 324396 327828 324460
rect 330340 324396 330404 324460
rect 373764 324396 373828 324460
rect 277900 323580 277964 323644
rect 323716 322900 323780 322964
rect 279556 322220 279620 322284
rect 288940 321948 289004 322012
rect 293356 321948 293420 322012
rect 321692 321948 321756 322012
rect 325188 321948 325252 322012
rect 282684 321812 282748 321876
rect 284340 321812 284404 321876
rect 288572 321812 288636 321876
rect 298324 321812 298388 321876
rect 324084 321812 324148 321876
rect 330708 321812 330772 321876
rect 301268 321676 301332 321740
rect 321508 321676 321572 321740
rect 282684 321540 282748 321604
rect 284524 321540 284588 321604
rect 286364 321540 286428 321604
rect 290596 321540 290660 321604
rect 299060 321540 299124 321604
rect 326660 321540 326724 321604
rect 330524 321540 330588 321604
rect 288940 321268 289004 321332
rect 291148 321404 291212 321468
rect 292620 321268 292684 321332
rect 293356 321268 293420 321332
rect 314516 321268 314580 321332
rect 320220 321404 320284 321468
rect 283236 320996 283300 321060
rect 288572 320996 288636 321060
rect 288388 320860 288452 320924
rect 282684 320784 282748 320788
rect 282684 320728 282688 320784
rect 282688 320728 282744 320784
rect 282744 320728 282748 320784
rect 282684 320724 282748 320728
rect 283972 320784 284036 320788
rect 283972 320728 283976 320784
rect 283976 320728 284032 320784
rect 284032 320728 284036 320784
rect 283972 320724 284036 320728
rect 285076 320724 285140 320788
rect 287468 320724 287532 320788
rect 288204 320724 288268 320788
rect 288572 320724 288636 320788
rect 289308 320784 289372 320788
rect 289308 320728 289312 320784
rect 289312 320728 289368 320784
rect 289368 320728 289372 320784
rect 289308 320724 289372 320728
rect 284708 320648 284772 320652
rect 284708 320592 284712 320648
rect 284712 320592 284768 320648
rect 284768 320592 284772 320648
rect 284708 320588 284772 320592
rect 284892 320588 284956 320652
rect 287468 320588 287532 320652
rect 290964 321132 291028 321196
rect 294276 321132 294340 321196
rect 295012 321132 295076 321196
rect 350764 321268 350828 321332
rect 298324 320996 298388 321060
rect 291884 320724 291948 320788
rect 292620 320724 292684 320788
rect 297220 320724 297284 320788
rect 292436 320588 292500 320652
rect 293172 320588 293236 320652
rect 295564 320588 295628 320652
rect 299244 320724 299308 320788
rect 298324 320588 298388 320652
rect 298508 320648 298572 320652
rect 298508 320592 298512 320648
rect 298512 320592 298568 320648
rect 298568 320592 298572 320648
rect 298508 320588 298572 320592
rect 299244 320648 299308 320652
rect 299244 320592 299248 320648
rect 299248 320592 299304 320648
rect 299304 320592 299308 320648
rect 299244 320588 299308 320592
rect 301268 320784 301332 320788
rect 301268 320728 301272 320784
rect 301272 320728 301328 320784
rect 301328 320728 301332 320784
rect 301268 320724 301332 320728
rect 304764 320784 304828 320788
rect 304764 320728 304768 320784
rect 304768 320728 304824 320784
rect 304824 320728 304828 320784
rect 304764 320724 304828 320728
rect 306420 320724 306484 320788
rect 306972 320724 307036 320788
rect 310652 320724 310716 320788
rect 311756 320724 311820 320788
rect 314516 320724 314580 320788
rect 315436 320724 315500 320788
rect 321508 320860 321572 320924
rect 325556 320860 325620 320924
rect 321692 320784 321756 320788
rect 321692 320728 321696 320784
rect 321696 320728 321752 320784
rect 321752 320728 321756 320784
rect 321692 320724 321756 320728
rect 322060 320724 322124 320788
rect 324084 320784 324148 320788
rect 324084 320728 324088 320784
rect 324088 320728 324144 320784
rect 324144 320728 324148 320784
rect 324084 320724 324148 320728
rect 325188 320784 325252 320788
rect 325188 320728 325192 320784
rect 325192 320728 325248 320784
rect 325248 320728 325252 320784
rect 325188 320724 325252 320728
rect 326660 320724 326724 320788
rect 327396 320784 327460 320788
rect 327396 320728 327400 320784
rect 327400 320728 327456 320784
rect 327456 320728 327460 320784
rect 327396 320724 327460 320728
rect 304028 320588 304092 320652
rect 305868 320588 305932 320652
rect 313596 320588 313660 320652
rect 320220 320588 320284 320652
rect 324820 320588 324884 320652
rect 300348 320452 300412 320516
rect 301636 320452 301700 320516
rect 305684 320452 305748 320516
rect 327580 320588 327644 320652
rect 312308 320452 312372 320516
rect 313964 320452 314028 320516
rect 318932 320452 318996 320516
rect 319852 320452 319916 320516
rect 323164 320452 323228 320516
rect 324636 320452 324700 320516
rect 326844 320452 326908 320516
rect 327764 320512 327828 320516
rect 327764 320456 327778 320512
rect 327778 320456 327828 320512
rect 327764 320452 327828 320456
rect 283788 320044 283852 320108
rect 284524 320044 284588 320108
rect 283604 319908 283668 319972
rect 284340 319908 284404 319972
rect 286548 320180 286612 320244
rect 287284 320240 287348 320244
rect 287284 320184 287288 320240
rect 287288 320184 287344 320240
rect 287344 320184 287348 320240
rect 287284 320180 287348 320184
rect 288388 320180 288452 320244
rect 308260 320316 308324 320380
rect 309180 320316 309244 320380
rect 310284 320316 310348 320380
rect 311204 320316 311268 320380
rect 285628 320104 285692 320108
rect 285628 320048 285632 320104
rect 285632 320048 285688 320104
rect 285688 320048 285692 320104
rect 285628 320044 285692 320048
rect 286732 320044 286796 320108
rect 286916 320104 286980 320108
rect 286916 320048 286920 320104
rect 286920 320048 286976 320104
rect 286976 320048 286980 320104
rect 286916 320044 286980 320048
rect 287652 320044 287716 320108
rect 285076 319636 285140 319700
rect 287468 319696 287532 319700
rect 287468 319640 287482 319696
rect 287482 319640 287532 319696
rect 287468 319636 287532 319640
rect 288020 319696 288084 319700
rect 288020 319640 288034 319696
rect 288034 319640 288084 319696
rect 288020 319636 288084 319640
rect 288940 320044 289004 320108
rect 289492 320044 289556 320108
rect 288572 319908 288636 319972
rect 288756 319636 288820 319700
rect 291148 320180 291212 320244
rect 292252 320180 292316 320244
rect 292988 320180 293052 320244
rect 293356 320180 293420 320244
rect 291332 320044 291396 320108
rect 292068 320044 292132 320108
rect 292620 320044 292684 320108
rect 294828 320180 294892 320244
rect 295012 320240 295076 320244
rect 295012 320184 295016 320240
rect 295016 320184 295072 320240
rect 295072 320184 295076 320240
rect 295012 320180 295076 320184
rect 295748 320180 295812 320244
rect 296300 320180 296364 320244
rect 298692 320240 298756 320244
rect 298692 320184 298696 320240
rect 298696 320184 298752 320240
rect 298752 320184 298756 320240
rect 294276 320044 294340 320108
rect 294460 320044 294524 320108
rect 295196 320044 295260 320108
rect 295380 320044 295444 320108
rect 296484 320044 296548 320108
rect 290780 319908 290844 319972
rect 290780 319772 290844 319836
rect 292988 319908 293052 319972
rect 298692 320180 298756 320184
rect 299428 320180 299492 320244
rect 300164 320240 300228 320244
rect 300164 320184 300168 320240
rect 300168 320184 300224 320240
rect 300224 320184 300228 320240
rect 300164 320180 300228 320184
rect 302740 320240 302804 320244
rect 302740 320184 302744 320240
rect 302744 320184 302800 320240
rect 302800 320184 302804 320240
rect 296852 320044 296916 320108
rect 297588 320104 297652 320108
rect 297588 320048 297592 320104
rect 297592 320048 297648 320104
rect 297648 320048 297652 320104
rect 297588 320044 297652 320048
rect 297772 320104 297836 320108
rect 297772 320048 297776 320104
rect 297776 320048 297832 320104
rect 297832 320048 297836 320104
rect 297772 320044 297836 320048
rect 298140 320044 298204 320108
rect 298876 320044 298940 320108
rect 299060 320104 299124 320108
rect 299060 320048 299064 320104
rect 299064 320048 299120 320104
rect 299120 320048 299124 320104
rect 299060 320044 299124 320048
rect 299796 320044 299860 320108
rect 300532 320044 300596 320108
rect 300900 320104 300964 320108
rect 300900 320048 300904 320104
rect 300904 320048 300960 320104
rect 300960 320048 300964 320104
rect 300900 320044 300964 320048
rect 302004 320044 302068 320108
rect 298876 319908 298940 319972
rect 302740 320180 302804 320184
rect 304764 320180 304828 320244
rect 305500 320180 305564 320244
rect 306788 320180 306852 320244
rect 308444 320240 308508 320244
rect 308444 320184 308448 320240
rect 308448 320184 308504 320240
rect 308504 320184 308508 320240
rect 308444 320180 308508 320184
rect 308628 320240 308692 320244
rect 308628 320184 308632 320240
rect 308632 320184 308688 320240
rect 308688 320184 308692 320240
rect 308628 320180 308692 320184
rect 309364 320180 309428 320244
rect 312676 320180 312740 320244
rect 313780 320180 313844 320244
rect 315620 320180 315684 320244
rect 316356 320180 316420 320244
rect 319668 320180 319732 320244
rect 319852 320240 319916 320244
rect 319852 320184 319856 320240
rect 319856 320184 319912 320240
rect 319912 320184 319916 320240
rect 319852 320180 319916 320184
rect 320588 320240 320652 320244
rect 320588 320184 320592 320240
rect 320592 320184 320648 320240
rect 320648 320184 320652 320240
rect 320588 320180 320652 320184
rect 322980 320316 323044 320380
rect 323532 320376 323596 320380
rect 323532 320320 323536 320376
rect 323536 320320 323592 320376
rect 323592 320320 323596 320376
rect 323532 320316 323596 320320
rect 324268 320316 324332 320380
rect 325188 320316 325252 320380
rect 302556 320044 302620 320108
rect 303292 320044 303356 320108
rect 303660 320104 303724 320108
rect 303660 320048 303664 320104
rect 303664 320048 303720 320104
rect 303720 320048 303724 320104
rect 303660 320044 303724 320048
rect 305132 320044 305196 320108
rect 306236 320044 306300 320108
rect 306972 320104 307036 320108
rect 306972 320048 306976 320104
rect 306976 320048 307032 320104
rect 307032 320048 307036 320104
rect 306972 320044 307036 320048
rect 307340 320104 307404 320108
rect 307340 320048 307344 320104
rect 307344 320048 307400 320104
rect 307400 320048 307404 320104
rect 307340 320044 307404 320048
rect 308076 320104 308140 320108
rect 308076 320048 308080 320104
rect 308080 320048 308136 320104
rect 308136 320048 308140 320104
rect 308076 320044 308140 320048
rect 308996 320044 309060 320108
rect 309548 320044 309612 320108
rect 310100 320044 310164 320108
rect 310836 320044 310900 320108
rect 312124 320104 312188 320108
rect 312124 320048 312128 320104
rect 312128 320048 312184 320104
rect 312184 320048 312188 320104
rect 312124 320044 312188 320048
rect 312492 320044 312556 320108
rect 314148 320044 314212 320108
rect 314700 320044 314764 320108
rect 316908 320044 316972 320108
rect 317644 320044 317708 320108
rect 319300 320044 319364 320108
rect 319484 320104 319548 320108
rect 319484 320048 319488 320104
rect 319488 320048 319544 320104
rect 319544 320048 319548 320104
rect 319484 320044 319548 320048
rect 320036 320104 320100 320108
rect 320036 320048 320040 320104
rect 320040 320048 320096 320104
rect 320096 320048 320100 320104
rect 320036 320044 320100 320048
rect 320956 320044 321020 320108
rect 321324 320104 321388 320108
rect 321324 320048 321328 320104
rect 321328 320048 321384 320104
rect 321384 320048 321388 320104
rect 321324 320044 321388 320048
rect 322796 320104 322860 320108
rect 322796 320048 322800 320104
rect 322800 320048 322856 320104
rect 322856 320048 322860 320104
rect 322796 320044 322860 320048
rect 323532 320044 323596 320108
rect 324452 320104 324516 320108
rect 324452 320048 324456 320104
rect 324456 320048 324512 320104
rect 324512 320048 324516 320104
rect 324452 320044 324516 320048
rect 325372 320044 325436 320108
rect 306052 319908 306116 319972
rect 325004 319908 325068 319972
rect 325372 319908 325436 319972
rect 295196 319772 295260 319836
rect 327212 320044 327276 320108
rect 326660 319908 326724 319972
rect 327580 319968 327644 319972
rect 327580 319912 327594 319968
rect 327594 319912 327644 319968
rect 327580 319908 327644 319912
rect 283788 319364 283852 319428
rect 294828 319364 294892 319428
rect 295564 319364 295628 319428
rect 297956 319364 298020 319428
rect 300164 319364 300228 319428
rect 300532 319424 300596 319428
rect 300532 319368 300546 319424
rect 300546 319368 300596 319424
rect 300532 319364 300596 319368
rect 301636 319364 301700 319428
rect 305500 319500 305564 319564
rect 305868 319500 305932 319564
rect 306052 319560 306116 319564
rect 306052 319504 306102 319560
rect 306102 319504 306116 319560
rect 306052 319500 306116 319504
rect 306788 319560 306852 319564
rect 306788 319504 306802 319560
rect 306802 319504 306852 319560
rect 306788 319500 306852 319504
rect 307892 319560 307956 319564
rect 307892 319504 307942 319560
rect 307942 319504 307956 319560
rect 307892 319500 307956 319504
rect 308444 319500 308508 319564
rect 309364 319500 309428 319564
rect 309548 319500 309612 319564
rect 313964 319560 314028 319564
rect 313964 319504 314014 319560
rect 314014 319504 314028 319560
rect 313964 319500 314028 319504
rect 317276 319500 317340 319564
rect 320588 319560 320652 319564
rect 320588 319504 320638 319560
rect 320638 319504 320652 319560
rect 320588 319500 320652 319504
rect 323532 319560 323596 319564
rect 323532 319504 323546 319560
rect 323546 319504 323596 319560
rect 323532 319500 323596 319504
rect 323716 319560 323780 319564
rect 323716 319504 323766 319560
rect 323766 319504 323780 319560
rect 323716 319500 323780 319504
rect 325372 319560 325436 319564
rect 325372 319504 325386 319560
rect 325386 319504 325436 319560
rect 325372 319500 325436 319504
rect 326660 319560 326724 319564
rect 326660 319504 326674 319560
rect 326674 319504 326724 319560
rect 326660 319500 326724 319504
rect 327212 319500 327276 319564
rect 327396 319560 327460 319564
rect 327396 319504 327446 319560
rect 327446 319504 327460 319560
rect 327396 319500 327460 319504
rect 307340 319424 307404 319428
rect 307340 319368 307354 319424
rect 307354 319368 307404 319424
rect 307340 319364 307404 319368
rect 308628 319364 308692 319428
rect 309732 319424 309796 319428
rect 309732 319368 309746 319424
rect 309746 319368 309796 319424
rect 309732 319364 309796 319368
rect 311204 319364 311268 319428
rect 312308 319424 312372 319428
rect 312308 319368 312322 319424
rect 312322 319368 312372 319424
rect 312308 319364 312372 319368
rect 313596 319364 313660 319428
rect 283420 319228 283484 319292
rect 283972 319228 284036 319292
rect 285628 319228 285692 319292
rect 286916 319228 286980 319292
rect 288388 319228 288452 319292
rect 288572 319228 288636 319292
rect 292620 319288 292684 319292
rect 292620 319232 292670 319288
rect 292670 319232 292684 319288
rect 283236 318956 283300 319020
rect 283604 318956 283668 319020
rect 284708 319016 284772 319020
rect 284708 318960 284758 319016
rect 284758 318960 284772 319016
rect 284708 318956 284772 318960
rect 284892 318956 284956 319020
rect 287284 319016 287348 319020
rect 287284 318960 287298 319016
rect 287298 318960 287348 319016
rect 287284 318956 287348 318960
rect 288940 318956 289004 319020
rect 290596 318820 290660 318884
rect 291148 319092 291212 319156
rect 292252 319092 292316 319156
rect 292620 319228 292684 319232
rect 292988 319288 293052 319292
rect 292988 319232 293002 319288
rect 293002 319232 293052 319288
rect 292988 319228 293052 319232
rect 295012 319228 295076 319292
rect 295380 319228 295444 319292
rect 295748 319016 295812 319020
rect 295748 318960 295762 319016
rect 295762 318960 295812 319016
rect 295748 318956 295812 318960
rect 297404 319016 297468 319020
rect 297404 318960 297418 319016
rect 297418 318960 297468 319016
rect 297404 318956 297468 318960
rect 297772 319016 297836 319020
rect 297772 318960 297786 319016
rect 297786 318960 297836 319016
rect 297772 318956 297836 318960
rect 298692 319016 298756 319020
rect 298692 318960 298742 319016
rect 298742 318960 298756 319016
rect 298692 318956 298756 318960
rect 300348 318956 300412 319020
rect 304764 318956 304828 319020
rect 305684 318956 305748 319020
rect 308260 319016 308324 319020
rect 308260 318960 308274 319016
rect 308274 318960 308324 319016
rect 308260 318956 308324 318960
rect 312124 319016 312188 319020
rect 312124 318960 312138 319016
rect 312138 318960 312188 319016
rect 312124 318956 312188 318960
rect 319484 318956 319548 319020
rect 319852 318956 319916 319020
rect 324452 318956 324516 319020
rect 325004 318956 325068 319020
rect 295196 318820 295260 318884
rect 298508 318820 298572 318884
rect 299796 318820 299860 318884
rect 307892 318820 307956 318884
rect 320036 318820 320100 318884
rect 324636 318820 324700 318884
rect 324820 318820 324884 318884
rect 325188 318820 325252 318884
rect 328500 318820 328564 318884
rect 283420 318684 283484 318748
rect 287836 318684 287900 318748
rect 294644 318744 294708 318748
rect 294644 318688 294658 318744
rect 294658 318688 294708 318744
rect 236500 318412 236564 318476
rect 292804 318548 292868 318612
rect 294644 318684 294708 318688
rect 296668 318684 296732 318748
rect 297956 318684 298020 318748
rect 300716 318684 300780 318748
rect 307524 318684 307588 318748
rect 308076 318684 308140 318748
rect 314332 318684 314396 318748
rect 325556 318744 325620 318748
rect 325556 318688 325570 318744
rect 325570 318688 325620 318744
rect 325556 318684 325620 318688
rect 237972 318276 238036 318340
rect 285812 318276 285876 318340
rect 292068 318276 292132 318340
rect 296852 318412 296916 318476
rect 300716 318412 300780 318476
rect 306972 318412 307036 318476
rect 323348 318548 323412 318612
rect 321324 318276 321388 318340
rect 285628 318004 285692 318068
rect 286548 318004 286612 318068
rect 289124 318004 289188 318068
rect 290596 318064 290660 318068
rect 290596 318008 290610 318064
rect 290610 318008 290660 318064
rect 290596 318004 290660 318008
rect 292436 318004 292500 318068
rect 302740 318004 302804 318068
rect 304764 318004 304828 318068
rect 284524 317868 284588 317932
rect 287100 317868 287164 317932
rect 288388 317868 288452 317932
rect 306604 317868 306668 317932
rect 315068 318004 315132 318068
rect 316540 318004 316604 318068
rect 317460 318004 317524 318068
rect 326660 318004 326724 318068
rect 318748 317928 318812 317932
rect 318748 317872 318798 317928
rect 318798 317872 318812 317928
rect 318748 317868 318812 317872
rect 320772 317868 320836 317932
rect 322796 317928 322860 317932
rect 322796 317872 322846 317928
rect 322846 317872 322860 317928
rect 322796 317868 322860 317872
rect 324452 317868 324516 317932
rect 367692 318140 367756 318204
rect 369900 318004 369964 318068
rect 327580 317868 327644 317932
rect 328684 317868 328748 317932
rect 300532 317792 300596 317796
rect 300532 317736 300582 317792
rect 300582 317736 300596 317792
rect 300532 317732 300596 317736
rect 301268 317732 301332 317796
rect 303292 317792 303356 317796
rect 303292 317736 303342 317792
rect 303342 317736 303356 317792
rect 303292 317732 303356 317736
rect 305316 317732 305380 317796
rect 307708 317732 307772 317796
rect 309732 317732 309796 317796
rect 310284 317732 310348 317796
rect 312860 317792 312924 317796
rect 312860 317736 312910 317792
rect 312910 317736 312924 317792
rect 312860 317732 312924 317736
rect 316172 317732 316236 317796
rect 318196 317732 318260 317796
rect 325556 317732 325620 317796
rect 327028 317732 327092 317796
rect 322796 317596 322860 317660
rect 283052 317460 283116 317524
rect 284340 317460 284404 317524
rect 290780 317460 290844 317524
rect 291700 317460 291764 317524
rect 299612 317460 299676 317524
rect 301084 317460 301148 317524
rect 302004 317460 302068 317524
rect 302740 317460 302804 317524
rect 303476 317460 303540 317524
rect 305500 317460 305564 317524
rect 306788 317520 306852 317524
rect 306788 317464 306838 317520
rect 306838 317464 306852 317520
rect 306788 317460 306852 317464
rect 308260 317460 308324 317524
rect 309732 317520 309796 317524
rect 309732 317464 309782 317520
rect 309782 317464 309796 317520
rect 309732 317460 309796 317464
rect 309916 317520 309980 317524
rect 309916 317464 309966 317520
rect 309966 317464 309980 317520
rect 309916 317460 309980 317464
rect 313044 317460 313108 317524
rect 313412 317460 313476 317524
rect 314516 317520 314580 317524
rect 314516 317464 314530 317520
rect 314530 317464 314580 317520
rect 314516 317460 314580 317464
rect 318380 317460 318444 317524
rect 320588 317460 320652 317524
rect 322612 317520 322676 317524
rect 322612 317464 322662 317520
rect 322662 317464 322676 317520
rect 223252 317052 223316 317116
rect 223436 316916 223500 316980
rect 287652 317324 287716 317388
rect 292436 317324 292500 317388
rect 322612 317460 322676 317464
rect 326844 317520 326908 317524
rect 326844 317464 326858 317520
rect 326858 317464 326908 317520
rect 326844 317460 326908 317464
rect 303660 317188 303724 317252
rect 281396 316916 281460 316980
rect 326660 316916 326724 316980
rect 325556 316780 325620 316844
rect 340828 316644 340892 316708
rect 299428 316508 299492 316572
rect 299244 316372 299308 316436
rect 298876 316236 298940 316300
rect 222700 315964 222764 316028
rect 298508 315964 298572 316028
rect 296484 315828 296548 315892
rect 296300 315692 296364 315756
rect 310100 315752 310164 315756
rect 310100 315696 310114 315752
rect 310114 315696 310164 315752
rect 310100 315692 310164 315696
rect 236684 315556 236748 315620
rect 297036 315556 297100 315620
rect 365116 315556 365180 315620
rect 237052 315420 237116 315484
rect 297404 315420 297468 315484
rect 352420 315420 352484 315484
rect 224724 315148 224788 315212
rect 301084 315148 301148 315212
rect 244780 314604 244844 314668
rect 288204 314604 288268 314668
rect 306788 314604 306852 314668
rect 312492 314664 312556 314668
rect 312492 314608 312506 314664
rect 312506 314608 312556 314664
rect 312492 314604 312556 314608
rect 312860 314604 312924 314668
rect 232268 314468 232332 314532
rect 301268 314468 301332 314532
rect 312676 314468 312740 314532
rect 232820 314332 232884 314396
rect 245516 314196 245580 314260
rect 304580 314196 304644 314260
rect 242572 314060 242636 314124
rect 302556 314060 302620 314124
rect 241284 313924 241348 313988
rect 356836 313924 356900 313988
rect 242756 313788 242820 313852
rect 234108 313108 234172 313172
rect 293356 313108 293420 313172
rect 309732 313168 309796 313172
rect 309732 313112 309782 313168
rect 309782 313112 309796 313168
rect 309732 313108 309796 313112
rect 320772 313108 320836 313172
rect 323164 313108 323228 313172
rect 249564 312972 249628 313036
rect 309180 312972 309244 313036
rect 251036 312836 251100 312900
rect 234476 312700 234540 312764
rect 294644 312700 294708 312764
rect 316172 312700 316236 312764
rect 233556 312564 233620 312628
rect 294276 312564 294340 312628
rect 315068 312564 315132 312628
rect 233740 312428 233804 312492
rect 294460 312428 294524 312492
rect 250852 312292 250916 312356
rect 232636 311748 232700 311812
rect 259316 311476 259380 311540
rect 231532 311340 231596 311404
rect 231716 311204 231780 311268
rect 231164 311068 231228 311132
rect 291700 311068 291764 311132
rect 313780 311068 313844 311132
rect 322612 311068 322676 311132
rect 291884 310932 291948 310996
rect 227484 310388 227548 310452
rect 297588 310388 297652 310452
rect 326844 310388 326908 310452
rect 239996 310252 240060 310316
rect 299612 310252 299676 310316
rect 226196 310116 226260 310180
rect 241100 309980 241164 310044
rect 300532 309980 300596 310044
rect 375972 309980 376036 310044
rect 231348 309844 231412 309908
rect 291332 309844 291396 309908
rect 230244 309708 230308 309772
rect 290780 309708 290844 309772
rect 228956 309572 229020 309636
rect 328684 309436 328748 309500
rect 284340 309028 284404 309092
rect 358308 308756 358372 308820
rect 319668 308620 319732 308684
rect 270356 308484 270420 308548
rect 356468 308348 356532 308412
rect 281396 307668 281460 307732
rect 302740 307668 302804 307732
rect 362724 307668 362788 307732
rect 282868 307532 282932 307596
rect 322796 307532 322860 307596
rect 380940 307532 381004 307596
rect 369164 307396 369228 307460
rect 359412 307260 359476 307324
rect 271092 307124 271156 307188
rect 313412 306988 313476 307052
rect 345060 306988 345124 307052
rect 327580 306444 327644 306508
rect 364932 306308 364996 306372
rect 363460 306172 363524 306236
rect 358124 306036 358188 306100
rect 223988 305764 224052 305828
rect 357940 305900 358004 305964
rect 356652 305764 356716 305828
rect 246988 304948 247052 305012
rect 320588 304948 320652 305012
rect 301452 304812 301516 304876
rect 360700 304812 360764 304876
rect 377260 304540 377324 304604
rect 246804 304132 246868 304196
rect 305500 304132 305564 304196
rect 317460 303512 317524 303516
rect 317460 303456 317510 303512
rect 317510 303456 317524 303512
rect 317460 303452 317524 303456
rect 367324 303316 367388 303380
rect 304764 302908 304828 302972
rect 239444 302772 239508 302836
rect 358860 302092 358924 302156
rect 313044 301956 313108 302020
rect 235212 301548 235276 301612
rect 299612 301548 299676 301612
rect 300716 301608 300780 301612
rect 300716 301552 300766 301608
rect 300766 301552 300780 301608
rect 300716 301548 300780 301552
rect 240916 301412 240980 301476
rect 300900 301412 300964 301476
rect 317460 300732 317524 300796
rect 318380 300732 318444 300796
rect 271276 300188 271340 300252
rect 330708 300188 330772 300252
rect 269620 300052 269684 300116
rect 237788 299372 237852 299436
rect 309732 299372 309796 299436
rect 313780 299372 313844 299436
rect 314516 299372 314580 299436
rect 375420 299372 375484 299436
rect 292436 299236 292500 299300
rect 350580 299236 350644 299300
rect 349292 299100 349356 299164
rect 370452 298964 370516 299028
rect 318196 298828 318260 298892
rect 349108 298692 349172 298756
rect 223804 298012 223868 298076
rect 308260 298012 308324 298076
rect 303292 297876 303356 297940
rect 363092 297876 363156 297940
rect 303476 297740 303540 297804
rect 362908 297740 362972 297804
rect 307708 297604 307772 297668
rect 310284 297604 310348 297668
rect 362540 297604 362604 297668
rect 239260 297468 239324 297532
rect 368980 297468 369044 297532
rect 238340 297332 238404 297396
rect 298324 297332 298388 297396
rect 346348 296924 346412 296988
rect 227300 296516 227364 296580
rect 285628 296516 285692 296580
rect 225828 296380 225892 296444
rect 285812 296380 285876 296444
rect 227116 296244 227180 296308
rect 228772 296108 228836 296172
rect 226932 295972 226996 296036
rect 229692 295156 229756 295220
rect 288756 295156 288820 295220
rect 354444 295156 354508 295220
rect 223068 295020 223132 295084
rect 352052 295020 352116 295084
rect 227852 294884 227916 294948
rect 229876 294748 229940 294812
rect 317644 294748 317708 294812
rect 223620 294612 223684 294676
rect 347820 294612 347884 294676
rect 230060 294476 230124 294540
rect 228220 294340 228284 294404
rect 232452 294204 232516 294268
rect 291148 294340 291212 294404
rect 245148 293524 245212 293588
rect 304028 293524 304092 293588
rect 238156 293388 238220 293452
rect 298140 293388 298204 293452
rect 236868 293252 236932 293316
rect 239076 293116 239140 293180
rect 246620 291756 246684 291820
rect 306604 291756 306668 291820
rect 220124 291484 220188 291548
rect 219940 291348 220004 291412
rect 221228 291212 221292 291276
rect 279372 290668 279436 290732
rect 220676 290320 220740 290324
rect 220676 290264 220726 290320
rect 220726 290264 220740 290320
rect 220676 290260 220740 290264
rect 245700 290260 245764 290324
rect 245700 289852 245764 289916
rect 225460 289580 225524 289644
rect 246436 289640 246500 289644
rect 246436 289584 246450 289640
rect 246450 289584 246500 289640
rect 246436 289580 246500 289584
rect 247172 289580 247236 289644
rect 246252 289444 246316 289508
rect 247540 289444 247604 289508
rect 251772 289444 251836 289508
rect 252692 289444 252756 289508
rect 240732 289308 240796 289372
rect 244044 289308 244108 289372
rect 244964 289036 245028 289100
rect 246436 288628 246500 288692
rect 240732 288492 240796 288556
rect 250668 287676 250732 287740
rect 257108 286316 257172 286380
rect 316540 286316 316604 286380
rect 221228 282100 221292 282164
rect 220124 272444 220188 272508
rect 265020 271084 265084 271148
rect 256924 267140 256988 267204
rect 316356 267140 316420 267204
rect 255820 267004 255884 267068
rect 256372 265508 256436 265572
rect 314884 265508 314948 265572
rect 260604 264284 260668 264348
rect 318932 264284 318996 264348
rect 267596 264148 267660 264212
rect 259132 260068 259196 260132
rect 262812 258708 262876 258772
rect 287100 257484 287164 257548
rect 256188 257348 256252 257412
rect 260972 253132 261036 253196
rect 264468 250412 264532 250476
rect 327028 249188 327092 249252
rect 262260 249052 262324 249116
rect 290596 247828 290660 247892
rect 262444 246196 262508 246260
rect 289308 245380 289372 245444
rect 305132 245244 305196 245308
rect 316172 245108 316236 245172
rect 264836 244972 264900 245036
rect 266124 244836 266188 244900
rect 260788 243748 260852 243812
rect 322980 243748 323044 243812
rect 320956 243612 321020 243676
rect 265020 243476 265084 243540
rect 324452 243476 324516 243540
rect 267412 243068 267476 243132
rect 265940 242796 266004 242860
rect 263732 242660 263796 242724
rect 259868 242388 259932 242452
rect 257292 242252 257356 242316
rect 316908 242252 316972 242316
rect 219940 242116 220004 242180
rect 260236 242116 260300 242180
rect 264652 241980 264716 242044
rect 273852 241980 273916 242044
rect 222884 241708 222948 241772
rect 226012 241708 226076 241772
rect 237972 241708 238036 241772
rect 265756 241708 265820 241772
rect 273852 241708 273916 241772
rect 228220 241572 228284 241636
rect 231900 241572 231964 241636
rect 233004 241436 233068 241500
rect 232084 241300 232148 241364
rect 232636 241300 232700 241364
rect 234844 241572 234908 241636
rect 256556 241572 256620 241636
rect 271828 241572 271892 241636
rect 288388 241436 288452 241500
rect 226748 241164 226812 241228
rect 225276 241028 225340 241092
rect 232636 240892 232700 240956
rect 233372 240892 233436 240956
rect 292620 240892 292684 240956
rect 242020 240756 242084 240820
rect 233924 240620 233988 240684
rect 234292 240620 234356 240684
rect 328500 240756 328564 240820
rect 265388 240620 265452 240684
rect 235028 240484 235092 240548
rect 222700 240348 222764 240412
rect 223436 240348 223500 240412
rect 232636 240348 232700 240412
rect 238892 240348 238956 240412
rect 225276 240212 225340 240276
rect 228036 240212 228100 240276
rect 235212 240212 235276 240276
rect 236316 240212 236380 240276
rect 236868 240212 236932 240276
rect 224724 239804 224788 239868
rect 225276 239864 225340 239868
rect 225276 239808 225280 239864
rect 225280 239808 225336 239864
rect 225336 239808 225340 239864
rect 225276 239804 225340 239808
rect 225460 239864 225524 239868
rect 225460 239808 225464 239864
rect 225464 239808 225520 239864
rect 225520 239808 225524 239864
rect 225460 239804 225524 239808
rect 226380 240076 226444 240140
rect 269620 240348 269684 240412
rect 225828 239940 225892 240004
rect 227852 239940 227916 240004
rect 230428 239940 230492 240004
rect 233740 239940 233804 240004
rect 226564 239804 226628 239868
rect 227116 239864 227180 239868
rect 227116 239808 227120 239864
rect 227120 239808 227176 239864
rect 227176 239808 227180 239864
rect 227116 239804 227180 239808
rect 227852 239804 227916 239868
rect 228036 239864 228100 239868
rect 228036 239808 228050 239864
rect 228050 239808 228100 239864
rect 228036 239804 228100 239808
rect 229140 239804 229204 239868
rect 229876 239804 229940 239868
rect 230612 239864 230676 239868
rect 230612 239808 230616 239864
rect 230616 239808 230672 239864
rect 230672 239808 230676 239864
rect 230612 239804 230676 239808
rect 231716 239804 231780 239868
rect 232452 239804 232516 239868
rect 232820 239804 232884 239868
rect 233372 239804 233436 239868
rect 234108 239804 234172 239868
rect 234660 239804 234724 239868
rect 236316 239804 236380 239868
rect 237604 239864 237668 239868
rect 237604 239808 237608 239864
rect 237608 239808 237664 239864
rect 237664 239808 237668 239864
rect 237604 239804 237668 239808
rect 237788 239804 237852 239868
rect 239260 239842 239264 239868
rect 239264 239842 239320 239868
rect 239320 239842 239324 239868
rect 239260 239804 239324 239842
rect 239628 239842 239632 239868
rect 239632 239842 239688 239868
rect 239688 239842 239692 239868
rect 239628 239804 239692 239842
rect 223252 239668 223316 239732
rect 223436 239728 223500 239732
rect 223436 239672 223450 239728
rect 223450 239672 223500 239728
rect 223436 239668 223500 239672
rect 223804 239668 223868 239732
rect 224172 239668 224236 239732
rect 228772 239728 228836 239732
rect 228772 239672 228786 239728
rect 228786 239672 228836 239728
rect 228772 239668 228836 239672
rect 230612 239668 230676 239732
rect 231164 239728 231228 239732
rect 231164 239672 231178 239728
rect 231178 239672 231228 239728
rect 231164 239668 231228 239672
rect 231348 239728 231412 239732
rect 231348 239672 231398 239728
rect 231398 239672 231412 239728
rect 231348 239668 231412 239672
rect 232084 239668 232148 239732
rect 232268 239668 232332 239732
rect 234292 239668 234356 239732
rect 234476 239668 234540 239732
rect 235028 239668 235092 239732
rect 236684 239668 236748 239732
rect 238340 239728 238404 239732
rect 238340 239672 238390 239728
rect 238390 239672 238404 239728
rect 238340 239668 238404 239672
rect 238892 239668 238956 239732
rect 239812 239706 239816 239732
rect 239816 239706 239872 239732
rect 239872 239706 239876 239732
rect 239812 239668 239876 239706
rect 240548 239804 240612 239868
rect 241100 239804 241164 239868
rect 240548 239668 240612 239732
rect 240916 239668 240980 239732
rect 241100 239668 241164 239732
rect 242020 239804 242084 239868
rect 242572 239804 242636 239868
rect 241652 239668 241716 239732
rect 243492 239668 243556 239732
rect 244044 239728 244108 239732
rect 244044 239672 244058 239728
rect 244058 239672 244108 239728
rect 244044 239668 244108 239672
rect 245516 239804 245580 239868
rect 246068 239804 246132 239868
rect 246436 239804 246500 239868
rect 245884 239668 245948 239732
rect 246804 239668 246868 239732
rect 247356 239804 247420 239868
rect 247540 239804 247604 239868
rect 257108 239940 257172 240004
rect 248828 239804 248892 239868
rect 249932 239804 249996 239868
rect 250116 239804 250180 239868
rect 251956 239842 251960 239868
rect 251960 239842 252016 239868
rect 252016 239842 252020 239868
rect 251956 239804 252020 239842
rect 252692 239804 252756 239868
rect 253428 239804 253492 239868
rect 254716 239842 254720 239868
rect 254720 239842 254776 239868
rect 254776 239842 254780 239868
rect 254716 239804 254780 239842
rect 256004 239804 256068 239868
rect 258396 239940 258460 240004
rect 259316 239940 259380 240004
rect 261524 239940 261588 240004
rect 258764 239864 258828 239868
rect 258764 239808 258768 239864
rect 258768 239808 258824 239864
rect 258824 239808 258828 239864
rect 258764 239804 258828 239808
rect 259132 239804 259196 239868
rect 259684 239804 259748 239868
rect 260236 239804 260300 239868
rect 262812 239940 262876 240004
rect 271092 240076 271156 240140
rect 266308 239940 266372 240004
rect 262628 239864 262692 239868
rect 262628 239808 262632 239864
rect 262632 239808 262688 239864
rect 262688 239808 262692 239864
rect 262628 239804 262692 239808
rect 264652 239804 264716 239868
rect 265388 239864 265452 239868
rect 265388 239808 265392 239864
rect 265392 239808 265448 239864
rect 265448 239808 265452 239864
rect 265388 239804 265452 239808
rect 265756 239864 265820 239868
rect 265756 239808 265760 239864
rect 265760 239808 265816 239864
rect 265816 239808 265820 239864
rect 265756 239804 265820 239808
rect 266124 239804 266188 239868
rect 267596 239864 267660 239868
rect 267596 239808 267646 239864
rect 267646 239808 267660 239864
rect 267596 239804 267660 239808
rect 223068 239456 223132 239460
rect 223068 239400 223118 239456
rect 223118 239400 223132 239456
rect 223068 239396 223132 239400
rect 223620 239396 223684 239460
rect 226196 239396 226260 239460
rect 226564 239396 226628 239460
rect 226748 239456 226812 239460
rect 226748 239400 226798 239456
rect 226798 239400 226812 239456
rect 226748 239396 226812 239400
rect 227484 239396 227548 239460
rect 228220 239396 228284 239460
rect 229692 239456 229756 239460
rect 229692 239400 229706 239456
rect 229706 239400 229756 239456
rect 229692 239396 229756 239400
rect 231532 239396 231596 239460
rect 231900 239456 231964 239460
rect 231900 239400 231950 239456
rect 231950 239400 231964 239456
rect 231900 239396 231964 239400
rect 232084 239396 232148 239460
rect 232636 239396 232700 239460
rect 233004 239396 233068 239460
rect 233924 239396 233988 239460
rect 235396 239396 235460 239460
rect 237052 239456 237116 239460
rect 237052 239400 237102 239456
rect 237102 239400 237116 239456
rect 237052 239396 237116 239400
rect 238156 239396 238220 239460
rect 239076 239396 239140 239460
rect 239996 239396 240060 239460
rect 241284 239456 241348 239460
rect 241284 239400 241334 239456
rect 241334 239400 241348 239456
rect 241284 239396 241348 239400
rect 242756 239396 242820 239460
rect 244780 239396 244844 239460
rect 246252 239532 246316 239596
rect 247172 239532 247236 239596
rect 247908 239532 247972 239596
rect 248828 239532 248892 239596
rect 249564 239532 249628 239596
rect 250668 239592 250732 239596
rect 250668 239536 250682 239592
rect 250682 239536 250732 239592
rect 250668 239532 250732 239536
rect 251036 239532 251100 239596
rect 251772 239532 251836 239596
rect 255820 239668 255884 239732
rect 256556 239668 256620 239732
rect 256924 239668 256988 239732
rect 259500 239668 259564 239732
rect 259868 239668 259932 239732
rect 260788 239728 260852 239732
rect 260788 239672 260838 239728
rect 260838 239672 260852 239728
rect 260788 239668 260852 239672
rect 260972 239668 261036 239732
rect 262260 239728 262324 239732
rect 262260 239672 262274 239728
rect 262274 239672 262324 239728
rect 262260 239668 262324 239672
rect 266308 239668 266372 239732
rect 271828 239668 271892 239732
rect 249380 239396 249444 239460
rect 250116 239396 250180 239460
rect 250852 239396 250916 239460
rect 256188 239396 256252 239460
rect 257292 239396 257356 239460
rect 260604 239396 260668 239460
rect 261340 239396 261404 239460
rect 263180 239396 263244 239460
rect 227300 239320 227364 239324
rect 227300 239264 227350 239320
rect 227350 239264 227364 239320
rect 227300 239260 227364 239264
rect 233556 239260 233620 239324
rect 234660 239260 234724 239324
rect 237236 239260 237300 239324
rect 247172 239260 247236 239324
rect 229876 239124 229940 239188
rect 230060 239184 230124 239188
rect 230060 239128 230110 239184
rect 230110 239128 230124 239184
rect 230060 239124 230124 239128
rect 232452 239124 232516 239188
rect 233188 239124 233252 239188
rect 225460 238988 225524 239052
rect 226380 238988 226444 239052
rect 227116 238988 227180 239052
rect 228036 238988 228100 239052
rect 237236 238988 237300 239052
rect 244964 239124 245028 239188
rect 246068 239124 246132 239188
rect 249196 239184 249260 239188
rect 266124 239320 266188 239324
rect 266124 239264 266138 239320
rect 266138 239264 266188 239320
rect 266124 239260 266188 239264
rect 267412 239260 267476 239324
rect 249196 239128 249210 239184
rect 249210 239128 249260 239184
rect 249196 239124 249260 239128
rect 247540 238852 247604 238916
rect 256372 238988 256436 239052
rect 260972 238852 261036 238916
rect 262444 238852 262508 238916
rect 264100 238988 264164 239052
rect 264468 239048 264532 239052
rect 264468 238992 264482 239048
rect 264482 238992 264532 239048
rect 264468 238988 264532 238992
rect 265020 239048 265084 239052
rect 265020 238992 265034 239048
rect 265034 238992 265084 239048
rect 265020 238988 265084 238992
rect 222700 238716 222764 238780
rect 223988 238776 224052 238780
rect 223988 238720 224002 238776
rect 224002 238720 224052 238776
rect 223988 238716 224052 238720
rect 236500 238716 236564 238780
rect 237236 238776 237300 238780
rect 237236 238720 237250 238776
rect 237250 238720 237300 238776
rect 237236 238716 237300 238720
rect 239260 238716 239324 238780
rect 240732 238716 240796 238780
rect 265204 238716 265268 238780
rect 188292 238444 188356 238508
rect 226932 238580 226996 238644
rect 228956 238580 229020 238644
rect 230244 238580 230308 238644
rect 230612 238640 230676 238644
rect 230612 238584 230662 238640
rect 230662 238584 230676 238640
rect 230612 238580 230676 238584
rect 234660 238580 234724 238644
rect 245148 238580 245212 238644
rect 245516 238580 245580 238644
rect 247172 238580 247236 238644
rect 248276 238580 248340 238644
rect 250300 238580 250364 238644
rect 252692 238580 252756 238644
rect 255636 238580 255700 238644
rect 264836 238580 264900 238644
rect 223804 238444 223868 238508
rect 226012 238444 226076 238508
rect 230980 238368 231044 238372
rect 230980 238312 231030 238368
rect 231030 238312 231044 238368
rect 230980 238308 231044 238312
rect 264284 238444 264348 238508
rect 266308 238444 266372 238508
rect 186820 238172 186884 238236
rect 175780 238036 175844 238100
rect 259132 238172 259196 238236
rect 263732 238172 263796 238236
rect 175964 237900 176028 237964
rect 241652 237960 241716 237964
rect 241652 237904 241666 237960
rect 241666 237904 241716 237960
rect 241652 237900 241716 237904
rect 249564 237900 249628 237964
rect 262628 237900 262692 237964
rect 310652 238036 310716 238100
rect 177252 237628 177316 237692
rect 231164 237764 231228 237828
rect 237604 237764 237668 237828
rect 242020 237764 242084 237828
rect 246252 237764 246316 237828
rect 259684 237824 259748 237828
rect 259684 237768 259734 237824
rect 259734 237768 259748 237824
rect 259684 237764 259748 237768
rect 260604 237764 260668 237828
rect 267780 237764 267844 237828
rect 247908 237628 247972 237692
rect 252324 237628 252388 237692
rect 255452 237628 255516 237692
rect 265940 237628 266004 237692
rect 231348 237356 231412 237420
rect 251036 237356 251100 237420
rect 252692 237356 252756 237420
rect 258764 237356 258828 237420
rect 260420 237416 260484 237420
rect 260420 237360 260434 237416
rect 260434 237360 260484 237416
rect 260420 237356 260484 237360
rect 268332 237220 268396 237284
rect 244412 236948 244476 237012
rect 252140 236948 252204 237012
rect 247356 236872 247420 236876
rect 247356 236816 247406 236872
rect 247406 236816 247420 236872
rect 247356 236812 247420 236816
rect 258396 236812 258460 236876
rect 262076 236812 262140 236876
rect 165844 236676 165908 236740
rect 238156 236676 238220 236740
rect 262628 236676 262692 236740
rect 270356 236676 270420 236740
rect 173756 236540 173820 236604
rect 236500 236540 236564 236604
rect 251772 236540 251836 236604
rect 255268 236540 255332 236604
rect 227484 236268 227548 236332
rect 234844 236268 234908 236332
rect 256004 236268 256068 236332
rect 224356 235996 224420 236060
rect 235580 235996 235644 236060
rect 242756 235996 242820 236060
rect 247172 236056 247236 236060
rect 247172 236000 247222 236056
rect 247222 236000 247236 236056
rect 247172 235996 247236 236000
rect 247724 236056 247788 236060
rect 247724 236000 247774 236056
rect 247774 236000 247788 236056
rect 247724 235996 247788 236000
rect 250668 236056 250732 236060
rect 250668 236000 250718 236056
rect 250718 236000 250732 236056
rect 250668 235996 250732 236000
rect 242572 235724 242636 235788
rect 236316 235588 236380 235652
rect 243860 235588 243924 235652
rect 162900 235452 162964 235516
rect 244044 235452 244108 235516
rect 176516 235316 176580 235380
rect 239996 235316 240060 235380
rect 240916 235316 240980 235380
rect 231900 235044 231964 235108
rect 239628 235104 239692 235108
rect 239628 235048 239678 235104
rect 239678 235048 239692 235104
rect 239628 235044 239692 235048
rect 243492 235104 243556 235108
rect 243492 235048 243506 235104
rect 243506 235048 243556 235104
rect 243492 235044 243556 235048
rect 241100 234772 241164 234836
rect 234476 234636 234540 234700
rect 180380 234364 180444 234428
rect 184428 234228 184492 234292
rect 181484 233956 181548 234020
rect 180564 233820 180628 233884
rect 240364 233820 240428 233884
rect 182588 233684 182652 233748
rect 173572 233548 173636 233612
rect 232820 233548 232884 233612
rect 258580 233548 258644 233612
rect 173020 233412 173084 233476
rect 232268 233412 232332 233476
rect 257108 233412 257172 233476
rect 165476 233140 165540 233204
rect 229140 233140 229204 233204
rect 252692 233004 252756 233068
rect 191604 232868 191668 232932
rect 174308 232732 174372 232796
rect 237236 232732 237300 232796
rect 175044 232596 175108 232660
rect 251956 232596 252020 232660
rect 163820 232460 163884 232524
rect 193076 232460 193140 232524
rect 164740 232324 164804 232388
rect 194364 231916 194428 231980
rect 172284 231780 172348 231844
rect 230796 231840 230860 231844
rect 230796 231784 230846 231840
rect 230846 231784 230860 231840
rect 230796 231780 230860 231784
rect 237972 231840 238036 231844
rect 237972 231784 237986 231840
rect 237986 231784 238036 231840
rect 237972 231780 238036 231784
rect 174676 231644 174740 231708
rect 234292 231644 234356 231708
rect 166396 231508 166460 231572
rect 168236 231372 168300 231436
rect 166580 231236 166644 231300
rect 317460 231644 317524 231708
rect 165660 231100 165724 231164
rect 250668 231100 250732 231164
rect 327580 231236 327644 231300
rect 176148 230964 176212 231028
rect 255268 230284 255332 230348
rect 184612 230148 184676 230212
rect 271276 230148 271340 230212
rect 181300 230012 181364 230076
rect 249012 230012 249076 230076
rect 168788 229876 168852 229940
rect 168052 229740 168116 229804
rect 338252 228924 338316 228988
rect 330340 228788 330404 228852
rect 181116 228516 181180 228580
rect 240548 228516 240612 228580
rect 249748 228516 249812 228580
rect 251036 228516 251100 228580
rect 309180 228516 309244 228580
rect 225460 228380 225524 228444
rect 235580 228244 235644 228308
rect 259132 227564 259196 227628
rect 330524 227428 330588 227492
rect 248276 227292 248340 227356
rect 249748 227020 249812 227084
rect 183140 226884 183204 226948
rect 259132 226400 259196 226404
rect 259132 226344 259146 226400
rect 259146 226344 259196 226400
rect 259132 226340 259196 226344
rect 306420 226068 306484 226132
rect 254900 225932 254964 225996
rect 261708 225932 261772 225996
rect 260420 225796 260484 225860
rect 197124 225660 197188 225724
rect 255636 225660 255700 225724
rect 188844 225524 188908 225588
rect 234476 224844 234540 224908
rect 167684 224300 167748 224364
rect 313964 224708 314028 224772
rect 169340 224164 169404 224228
rect 260604 223484 260668 223548
rect 252140 223348 252204 223412
rect 252508 223348 252572 223412
rect 263364 223212 263428 223276
rect 321508 223076 321572 223140
rect 235396 222940 235460 223004
rect 234844 222804 234908 222868
rect 252508 222804 252572 222868
rect 252508 222668 252572 222732
rect 249012 222532 249076 222596
rect 249748 222532 249812 222596
rect 253428 222184 253492 222188
rect 253428 222128 253478 222184
rect 253478 222128 253492 222184
rect 253428 222124 253492 222128
rect 258396 221988 258460 222052
rect 259132 221988 259196 222052
rect 249380 221852 249444 221916
rect 252508 221716 252572 221780
rect 257108 221716 257172 221780
rect 249748 221580 249812 221644
rect 173204 221444 173268 221508
rect 259132 221036 259196 221100
rect 249196 220900 249260 220964
rect 178540 220764 178604 220828
rect 224356 220628 224420 220692
rect 249564 220764 249628 220828
rect 309732 220628 309796 220692
rect 246988 220492 247052 220556
rect 247724 220492 247788 220556
rect 307708 220492 307772 220556
rect 310836 220356 310900 220420
rect 169156 220220 169220 220284
rect 246988 220220 247052 220284
rect 314700 220220 314764 220284
rect 163636 220084 163700 220148
rect 255452 220084 255516 220148
rect 313780 220084 313844 220148
rect 291700 219948 291764 220012
rect 242204 219268 242268 219332
rect 301452 219268 301516 219332
rect 243860 219132 243924 219196
rect 302924 219132 302988 219196
rect 182956 218996 183020 219060
rect 244044 218996 244108 219060
rect 302740 218996 302804 219060
rect 165108 218860 165172 218924
rect 237972 218860 238036 218924
rect 296852 218860 296916 218924
rect 167868 218724 167932 218788
rect 299612 218724 299676 218788
rect 164924 218588 164988 218652
rect 239996 218588 240060 218652
rect 244044 218240 244108 218244
rect 244044 218184 244058 218240
rect 244058 218184 244108 218240
rect 244044 218180 244108 218184
rect 239996 218104 240060 218108
rect 239996 218048 240010 218104
rect 240010 218048 240060 218104
rect 239996 218044 240060 218048
rect 243860 218104 243924 218108
rect 243860 218048 243874 218104
rect 243874 218048 243924 218104
rect 243860 218044 243924 218048
rect 170996 217772 171060 217836
rect 168972 217636 169036 217700
rect 171732 217500 171796 217564
rect 170628 217364 170692 217428
rect 171916 217228 171980 217292
rect 172100 217092 172164 217156
rect 170812 216956 170876 217020
rect 318932 216548 318996 216612
rect 230980 216412 231044 216476
rect 259316 216276 259380 216340
rect 259316 215324 259380 215388
rect 196940 214916 197004 214980
rect 255820 214916 255884 214980
rect 195652 214780 195716 214844
rect 195836 214644 195900 214708
rect 170444 214508 170508 214572
rect 179092 213828 179156 213892
rect 178908 213692 178972 213756
rect 185164 213556 185228 213620
rect 244412 213556 244476 213620
rect 180196 213420 180260 213484
rect 239444 213420 239508 213484
rect 182772 213284 182836 213348
rect 174492 213148 174556 213212
rect 180012 213012 180076 213076
rect 203196 212060 203260 212124
rect 180932 211924 180996 211988
rect 178724 211788 178788 211852
rect 198412 210428 198476 210492
rect 190316 210292 190380 210356
rect 198044 210020 198108 210084
rect 199332 209748 199396 209812
rect 163452 209476 163516 209540
rect 184060 209476 184124 209540
rect 189580 209536 189644 209540
rect 189580 209480 189594 209536
rect 189594 209480 189644 209536
rect 189580 209476 189644 209480
rect 193812 209476 193876 209540
rect 195468 209476 195532 209540
rect 197860 209476 197924 209540
rect 199148 209536 199212 209540
rect 199148 209480 199198 209536
rect 199198 209480 199212 209536
rect 199148 209476 199212 209480
rect 199884 209536 199948 209540
rect 199884 209480 199898 209536
rect 199898 209480 199948 209536
rect 199884 209476 199948 209480
rect 189580 208932 189644 208996
rect 201356 207572 201420 207636
rect 203196 206212 203260 206276
rect 208900 204852 208964 204916
rect 207796 182820 207860 182884
rect 205772 179964 205836 180028
rect 205956 175884 206020 175948
rect 266308 175884 266372 175948
rect 207980 171668 208044 171732
rect 204852 170308 204916 170372
rect 204668 167588 204732 167652
rect 206140 166228 206204 166292
rect 205404 165004 205468 165068
rect 204116 164868 204180 164932
rect 203564 163508 203628 163572
rect 205220 163372 205284 163436
rect 203380 162284 203444 162348
rect 203196 162148 203260 162212
rect 206876 162012 206940 162076
rect 202644 161876 202708 161940
rect 169524 160652 169588 160716
rect 186820 160652 186884 160716
rect 164004 160380 164068 160444
rect 162716 160244 162780 160308
rect 171364 160244 171428 160308
rect 172284 160244 172348 160308
rect 162716 159836 162780 159900
rect 163452 159836 163516 159900
rect 163820 159836 163884 159900
rect 164004 159896 164068 159900
rect 165660 159972 165724 160036
rect 164004 159840 164054 159896
rect 164054 159840 164068 159896
rect 164004 159836 164068 159840
rect 164740 159836 164804 159900
rect 165844 159836 165908 159900
rect 166580 159896 166644 159900
rect 166580 159840 166594 159896
rect 166594 159840 166644 159896
rect 166580 159836 166644 159840
rect 167868 159836 167932 159900
rect 168052 159836 168116 159900
rect 169340 159972 169404 160036
rect 169156 159836 169220 159900
rect 169524 159896 169588 159900
rect 169524 159840 169574 159896
rect 169574 159840 169588 159896
rect 169524 159836 169588 159840
rect 162900 159760 162964 159764
rect 162900 159704 162914 159760
rect 162914 159704 162964 159760
rect 162900 159700 162964 159704
rect 163636 159700 163700 159764
rect 164556 159700 164620 159764
rect 165476 159700 165540 159764
rect 166396 159700 166460 159764
rect 168236 159700 168300 159764
rect 168972 159700 169036 159764
rect 168788 159564 168852 159628
rect 170260 159896 170324 159900
rect 170260 159840 170310 159896
rect 170310 159840 170324 159896
rect 170260 159836 170324 159840
rect 170812 159836 170876 159900
rect 175964 160108 176028 160172
rect 203564 161196 203628 161260
rect 198780 161060 198844 161124
rect 198044 160924 198108 160988
rect 171180 159836 171244 159900
rect 171548 159896 171612 159900
rect 171548 159840 171562 159896
rect 171562 159840 171612 159896
rect 171548 159836 171612 159840
rect 171732 159836 171796 159900
rect 172652 159896 172716 159900
rect 172652 159840 172666 159896
rect 172666 159840 172716 159896
rect 172652 159836 172716 159840
rect 173020 159836 173084 159900
rect 173204 159836 173268 159900
rect 173756 159896 173820 159900
rect 173756 159840 173770 159896
rect 173770 159840 173820 159896
rect 173756 159836 173820 159840
rect 174308 159896 174372 159900
rect 174308 159840 174322 159896
rect 174322 159840 174372 159896
rect 174308 159836 174372 159840
rect 174676 159836 174740 159900
rect 198780 160108 198844 160172
rect 175228 159836 175292 159900
rect 176516 159836 176580 159900
rect 178908 159836 178972 159900
rect 180380 159836 180444 159900
rect 180564 159896 180628 159900
rect 180564 159840 180614 159896
rect 180614 159840 180628 159896
rect 180564 159836 180628 159840
rect 181484 159836 181548 159900
rect 182588 159896 182652 159900
rect 182588 159840 182602 159896
rect 182602 159840 182652 159896
rect 182588 159836 182652 159840
rect 183140 159836 183204 159900
rect 184060 159836 184124 159900
rect 184612 159836 184676 159900
rect 185164 159836 185228 159900
rect 188476 159836 188540 159900
rect 188844 159836 188908 159900
rect 190316 159836 190380 159900
rect 193076 159836 193140 159900
rect 193628 159896 193692 159900
rect 193628 159840 193642 159896
rect 193642 159840 193692 159896
rect 193628 159836 193692 159840
rect 194364 159836 194428 159900
rect 195284 159896 195348 159900
rect 195284 159840 195298 159896
rect 195298 159840 195348 159896
rect 195284 159836 195348 159840
rect 195836 159896 195900 159900
rect 195836 159840 195850 159896
rect 195850 159840 195900 159896
rect 195836 159836 195900 159840
rect 197124 159836 197188 159900
rect 197860 159836 197924 159900
rect 198228 159836 198292 159900
rect 199148 159896 199212 159900
rect 199148 159840 199162 159896
rect 199162 159840 199212 159896
rect 199148 159836 199212 159840
rect 199884 159836 199948 159900
rect 200988 159836 201052 159900
rect 201356 159836 201420 159900
rect 170076 159700 170140 159764
rect 170628 159760 170692 159764
rect 170628 159704 170678 159760
rect 170678 159704 170692 159760
rect 170628 159700 170692 159704
rect 171364 159700 171428 159764
rect 171916 159700 171980 159764
rect 173572 159700 173636 159764
rect 174492 159700 174556 159764
rect 176332 159760 176396 159764
rect 176332 159704 176382 159760
rect 176382 159704 176396 159760
rect 176332 159700 176396 159704
rect 178540 159700 178604 159764
rect 180932 159700 180996 159764
rect 182772 159700 182836 159764
rect 184428 159700 184492 159764
rect 191604 159700 191668 159764
rect 195652 159700 195716 159764
rect 196388 159760 196452 159764
rect 196388 159704 196402 159760
rect 196402 159704 196452 159760
rect 196388 159700 196452 159704
rect 196940 159700 197004 159764
rect 198412 159700 198476 159764
rect 199332 159700 199396 159764
rect 203564 160244 203628 160308
rect 204116 159896 204180 159900
rect 204116 159840 204130 159896
rect 204130 159840 204180 159896
rect 204116 159836 204180 159840
rect 204668 159836 204732 159900
rect 205220 159896 205284 159900
rect 205220 159840 205234 159896
rect 205234 159840 205284 159896
rect 205220 159836 205284 159840
rect 205404 159896 205468 159900
rect 205404 159840 205454 159896
rect 205454 159840 205468 159896
rect 205404 159836 205468 159840
rect 205772 159836 205836 159900
rect 207980 159836 208044 159900
rect 202460 159760 202524 159764
rect 202460 159704 202474 159760
rect 202474 159704 202524 159760
rect 202460 159700 202524 159704
rect 202644 159760 202708 159764
rect 202644 159704 202694 159760
rect 202694 159704 202708 159760
rect 202644 159700 202708 159704
rect 204852 159700 204916 159764
rect 205956 159700 206020 159764
rect 207796 159700 207860 159764
rect 170444 159564 170508 159628
rect 172100 159564 172164 159628
rect 175044 159564 175108 159628
rect 181116 159564 181180 159628
rect 198044 159564 198108 159628
rect 175780 159428 175844 159492
rect 170996 159352 171060 159356
rect 177252 159428 177316 159492
rect 227668 159428 227732 159492
rect 170996 159296 171010 159352
rect 171010 159296 171060 159352
rect 170996 159292 171060 159296
rect 172468 159156 172532 159220
rect 203380 159156 203444 159220
rect 206140 159156 206204 159220
rect 192524 159020 192588 159084
rect 170076 158884 170140 158948
rect 171548 158944 171612 158948
rect 171548 158888 171562 158944
rect 171562 158888 171612 158944
rect 171548 158884 171612 158888
rect 199148 158884 199212 158948
rect 163452 158612 163516 158676
rect 164188 158672 164252 158676
rect 164188 158616 164238 158672
rect 164238 158616 164252 158672
rect 164188 158612 164252 158616
rect 164740 158672 164804 158676
rect 164740 158616 164790 158672
rect 164790 158616 164804 158672
rect 164740 158612 164804 158616
rect 165292 158612 165356 158676
rect 165660 158672 165724 158676
rect 165660 158616 165710 158672
rect 165710 158616 165724 158672
rect 165660 158612 165724 158616
rect 166028 158672 166092 158676
rect 166028 158616 166078 158672
rect 166078 158616 166092 158672
rect 166028 158612 166092 158616
rect 167684 158612 167748 158676
rect 188292 158748 188356 158812
rect 168420 158612 168484 158676
rect 168972 158612 169036 158676
rect 170260 158612 170324 158676
rect 171732 158612 171796 158676
rect 172284 158672 172348 158676
rect 172284 158616 172334 158672
rect 172334 158616 172348 158672
rect 172284 158612 172348 158616
rect 173204 158612 173268 158676
rect 175044 158612 175108 158676
rect 175412 158612 175476 158676
rect 176332 158612 176396 158676
rect 178724 158612 178788 158676
rect 180196 158612 180260 158676
rect 181300 158612 181364 158676
rect 182956 158612 183020 158676
rect 187004 158612 187068 158676
rect 187188 158672 187252 158676
rect 187188 158616 187238 158672
rect 187238 158616 187252 158672
rect 187188 158612 187252 158616
rect 187556 158672 187620 158676
rect 187556 158616 187570 158672
rect 187570 158616 187620 158672
rect 187556 158612 187620 158616
rect 188292 158612 188356 158676
rect 188660 158672 188724 158676
rect 188660 158616 188674 158672
rect 188674 158616 188724 158672
rect 188660 158612 188724 158616
rect 188844 158672 188908 158676
rect 188844 158616 188894 158672
rect 188894 158616 188908 158672
rect 188844 158612 188908 158616
rect 189580 158612 189644 158676
rect 189948 158672 190012 158676
rect 189948 158616 189998 158672
rect 189998 158616 190012 158672
rect 189948 158612 190012 158616
rect 190316 158672 190380 158676
rect 190316 158616 190330 158672
rect 190330 158616 190380 158672
rect 190316 158612 190380 158616
rect 191236 158612 191300 158676
rect 165108 158340 165172 158404
rect 168604 158476 168668 158540
rect 171916 158476 171980 158540
rect 172100 158536 172164 158540
rect 172100 158480 172150 158536
rect 172150 158480 172164 158536
rect 172100 158476 172164 158480
rect 174676 158476 174740 158540
rect 175228 158476 175292 158540
rect 176516 158476 176580 158540
rect 187372 158476 187436 158540
rect 191052 158476 191116 158540
rect 193076 158612 193140 158676
rect 194180 158672 194244 158676
rect 194180 158616 194194 158672
rect 194194 158616 194244 158672
rect 194180 158612 194244 158616
rect 194364 158672 194428 158676
rect 194364 158616 194414 158672
rect 194414 158616 194428 158672
rect 194364 158612 194428 158616
rect 195284 158612 195348 158676
rect 196756 158612 196820 158676
rect 196940 158612 197004 158676
rect 198412 158612 198476 158676
rect 198596 158672 198660 158676
rect 198596 158616 198646 158672
rect 198646 158616 198660 158672
rect 198596 158612 198660 158616
rect 199700 158612 199764 158676
rect 200804 158612 200868 158676
rect 202092 158672 202156 158676
rect 202092 158616 202142 158672
rect 202142 158616 202156 158672
rect 202092 158612 202156 158616
rect 203932 158612 203996 158676
rect 204116 158612 204180 158676
rect 205404 158612 205468 158676
rect 206876 158612 206940 158676
rect 192892 158476 192956 158540
rect 193996 158476 194060 158540
rect 195468 158476 195532 158540
rect 199516 158476 199580 158540
rect 201172 158476 201236 158540
rect 202276 158476 202340 158540
rect 203748 158476 203812 158540
rect 208900 158476 208964 158540
rect 168788 158340 168852 158404
rect 174308 158340 174372 158404
rect 191788 158340 191852 158404
rect 193628 158340 193692 158404
rect 195652 158340 195716 158404
rect 199332 158340 199396 158404
rect 201356 158340 201420 158404
rect 204116 158340 204180 158404
rect 172652 158204 172716 158268
rect 175228 158204 175292 158268
rect 192708 158204 192772 158268
rect 194548 158204 194612 158268
rect 172468 158068 172532 158132
rect 203564 158068 203628 158132
rect 179276 157932 179340 157996
rect 203196 157932 203260 157996
rect 245884 157932 245948 157996
rect 168236 157796 168300 157860
rect 177804 157796 177868 157860
rect 179092 157796 179156 157860
rect 238156 157796 238220 157860
rect 177252 157660 177316 157724
rect 178908 157720 178972 157724
rect 178908 157664 178958 157720
rect 178958 157664 178972 157720
rect 178908 157660 178972 157664
rect 180012 157660 180076 157724
rect 181116 157660 181180 157724
rect 164556 157448 164620 157452
rect 164556 157392 164606 157448
rect 164606 157392 164620 157448
rect 164556 157388 164620 157392
rect 164372 157252 164436 157316
rect 202460 157524 202524 157588
rect 206876 157524 206940 157588
rect 176148 157388 176212 157452
rect 177436 157388 177500 157452
rect 177620 157388 177684 157452
rect 179092 157388 179156 157452
rect 180012 157448 180076 157452
rect 180012 157392 180026 157448
rect 180026 157392 180076 157448
rect 180012 157388 180076 157392
rect 180564 157388 180628 157452
rect 181484 157388 181548 157452
rect 184244 157388 184308 157452
rect 184980 157448 185044 157452
rect 184980 157392 185030 157448
rect 185030 157392 185044 157448
rect 184980 157388 185044 157392
rect 173020 157252 173084 157316
rect 191420 157252 191484 157316
rect 162900 157116 162964 157180
rect 175412 156844 175476 156908
rect 167132 156708 167196 156772
rect 175412 155892 175476 155956
rect 203748 155756 203812 155820
rect 268332 155756 268396 155820
rect 179276 155620 179340 155684
rect 233188 155348 233252 155412
rect 273852 154260 273916 154324
rect 199700 153988 199764 154052
rect 240916 153988 240980 154052
rect 187004 153580 187068 153644
rect 196388 153172 196452 153236
rect 196940 153036 197004 153100
rect 195468 152900 195532 152964
rect 194548 152628 194612 152692
rect 198044 152492 198108 152556
rect 198596 152492 198660 152556
rect 193996 152356 194060 152420
rect 195284 152220 195348 152284
rect 179092 151268 179156 151332
rect 196756 150180 196820 150244
rect 177620 150044 177684 150108
rect 177436 149908 177500 149972
rect 177804 149772 177868 149836
rect 170996 148412 171060 148476
rect 230980 148412 231044 148476
rect 168972 147596 169036 147660
rect 203932 147324 203996 147388
rect 264284 147324 264348 147388
rect 173388 147188 173452 147252
rect 174492 147188 174556 147252
rect 173204 147052 173268 147116
rect 162900 146916 162964 146980
rect 187372 146916 187436 146980
rect 168788 146236 168852 146300
rect 175228 146236 175292 146300
rect 184244 146236 184308 146300
rect 168604 146100 168668 146164
rect 201172 146100 201236 146164
rect 260052 146100 260116 146164
rect 180012 145964 180076 146028
rect 176516 145828 176580 145892
rect 205404 145692 205468 145756
rect 267780 145692 267844 145756
rect 204116 144740 204180 144804
rect 262444 144604 262508 144668
rect 191788 144332 191852 144396
rect 191236 144196 191300 144260
rect 164372 144060 164436 144124
rect 178908 144060 178972 144124
rect 174308 143380 174372 143444
rect 202092 143380 202156 143444
rect 200804 143244 200868 143308
rect 261708 143244 261772 143308
rect 173020 143108 173084 143172
rect 259684 142972 259748 143036
rect 202276 142836 202340 142900
rect 261524 142836 261588 142900
rect 264100 142836 264164 142900
rect 171732 142700 171796 142764
rect 172284 142700 172348 142764
rect 189948 142564 190012 142628
rect 201356 142292 201420 142356
rect 261340 142156 261404 142220
rect 232636 142020 232700 142084
rect 188844 141884 188908 141948
rect 249380 141884 249444 141948
rect 187556 141748 187620 141812
rect 187188 141612 187252 141676
rect 174492 141476 174556 141540
rect 191420 141476 191484 141540
rect 170260 141340 170324 141404
rect 188660 141340 188724 141404
rect 190316 141204 190380 141268
rect 191052 140796 191116 140860
rect 168420 140660 168484 140724
rect 181484 140660 181548 140724
rect 242204 140660 242268 140724
rect 177252 140524 177316 140588
rect 237972 140524 238036 140588
rect 189764 140388 189828 140452
rect 246436 140388 246500 140452
rect 240732 140252 240796 140316
rect 242020 140116 242084 140180
rect 188292 139980 188356 140044
rect 178724 139844 178788 139908
rect 184980 139708 185044 139772
rect 198412 139708 198476 139772
rect 234660 139300 234724 139364
rect 195652 139164 195716 139228
rect 230428 139028 230492 139092
rect 167132 138892 167196 138956
rect 168236 138892 168300 138956
rect 166948 138620 167012 138684
rect 177804 138620 177868 138684
rect 194180 137804 194244 137868
rect 193076 137668 193140 137732
rect 166212 137592 166276 137596
rect 166212 137536 166226 137592
rect 166226 137536 166276 137592
rect 166212 137532 166276 137536
rect 192708 137532 192772 137596
rect 251772 137532 251836 137596
rect 192524 137396 192588 137460
rect 250300 137396 250364 137460
rect 167132 137260 167196 137324
rect 194364 137260 194428 137324
rect 192892 137124 192956 137188
rect 236500 137124 236564 137188
rect 177436 136580 177500 136644
rect 271828 136580 271892 136644
rect 173388 135900 173452 135964
rect 180196 135900 180260 135964
rect 171732 134404 171796 134468
rect 166212 131684 166276 131748
rect 199332 131684 199396 131748
rect 175780 131140 175844 131204
rect 164372 130324 164436 130388
rect 180380 130324 180444 130388
rect 182956 127604 183020 127668
rect 181116 126924 181180 126988
rect 173204 126244 173268 126308
rect 199516 125428 199580 125492
rect 182588 124748 182652 124812
rect 180564 124068 180628 124132
rect 182772 122164 182836 122228
rect 193996 122028 194060 122092
rect 177620 120804 177684 120868
rect 195284 120668 195348 120732
rect 187188 119444 187252 119508
rect 203748 119308 203812 119372
rect 196940 117948 197004 118012
rect 189764 115228 189828 115292
rect 198044 115092 198108 115156
rect 188292 113868 188356 113932
rect 165844 113732 165908 113796
rect 199700 113732 199764 113796
rect 166028 112372 166092 112436
rect 181484 112372 181548 112436
rect 331812 111828 331876 111892
rect 173020 111012 173084 111076
rect 200988 109652 201052 109716
rect 200804 106796 200868 106860
rect 187372 105436 187436 105500
rect 202276 104076 202340 104140
rect 188476 102716 188540 102780
rect 202460 101356 202524 101420
rect 181300 98772 181364 98836
rect 198228 98636 198292 98700
rect 203932 95780 203996 95844
rect 179092 91700 179156 91764
rect 205220 90340 205284 90404
rect 205772 84764 205836 84828
rect 280660 71844 280724 71908
rect 202644 71028 202708 71092
rect 204116 69532 204180 69596
rect 187556 68172 187620 68236
rect 188660 66812 188724 66876
rect 188844 65452 188908 65516
rect 190132 64092 190196 64156
rect 189948 62732 190012 62796
rect 335860 59332 335924 59396
rect 194180 54436 194244 54500
rect 194364 51716 194428 51780
rect 197860 46140 197924 46204
rect 198412 44780 198476 44844
rect 199884 42060 199948 42124
rect 190316 40564 190380 40628
rect 201172 37844 201236 37908
rect 205404 35124 205468 35188
rect 195468 30908 195532 30972
rect 177252 24108 177316 24172
rect 201356 18532 201420 18596
rect 197124 11596 197188 11660
rect 192708 9420 192772 9484
rect 192892 9284 192956 9348
rect 192524 9148 192588 9212
rect 195652 9012 195716 9076
rect 195100 8876 195164 8940
rect 205956 7516 206020 7580
rect 184612 6836 184676 6900
rect 184980 6700 185044 6764
rect 185164 6564 185228 6628
rect 191604 6428 191668 6492
rect 191420 6292 191484 6356
rect 193076 6156 193140 6220
rect 184428 6020 184492 6084
rect 179276 3572 179340 3636
rect 184244 3436 184308 3500
rect 184060 3300 184124 3364
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 705798 6134 705830
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -1894 6134 -1862
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 705798 42134 705830
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -1894 42134 -1862
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 705798 78134 705830
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -1894 78134 -1862
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 705798 114134 705830
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -1894 114134 -1862
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 705798 150134 705830
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 175779 238100 175845 238101
rect 175779 238036 175780 238100
rect 175844 238036 175845 238100
rect 175779 238035 175845 238036
rect 165843 236740 165909 236741
rect 165843 236676 165844 236740
rect 165908 236676 165909 236740
rect 165843 236675 165909 236676
rect 162899 235516 162965 235517
rect 162899 235452 162900 235516
rect 162964 235452 162965 235516
rect 162899 235451 162965 235452
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 162715 160308 162781 160309
rect 162715 160244 162716 160308
rect 162780 160244 162781 160308
rect 162715 160243 162781 160244
rect 162718 159901 162778 160243
rect 162715 159900 162781 159901
rect 162715 159836 162716 159900
rect 162780 159836 162781 159900
rect 162715 159835 162781 159836
rect 162902 159765 162962 235451
rect 165475 233204 165541 233205
rect 165475 233140 165476 233204
rect 165540 233140 165541 233204
rect 165475 233139 165541 233140
rect 163819 232524 163885 232525
rect 163819 232460 163820 232524
rect 163884 232460 163885 232524
rect 163819 232459 163885 232460
rect 163635 220148 163701 220149
rect 163635 220084 163636 220148
rect 163700 220084 163701 220148
rect 163635 220083 163701 220084
rect 163451 209540 163517 209541
rect 163451 209476 163452 209540
rect 163516 209476 163517 209540
rect 163451 209475 163517 209476
rect 163454 159901 163514 209475
rect 163451 159900 163517 159901
rect 163451 159836 163452 159900
rect 163516 159836 163517 159900
rect 163451 159835 163517 159836
rect 162899 159764 162965 159765
rect 162899 159700 162900 159764
rect 162964 159700 162965 159764
rect 162899 159699 162965 159700
rect 163454 158677 163514 159835
rect 163638 159765 163698 220083
rect 163822 159901 163882 232459
rect 164739 232388 164805 232389
rect 164739 232324 164740 232388
rect 164804 232324 164805 232388
rect 164739 232323 164805 232324
rect 164208 183454 164528 183486
rect 164208 183218 164250 183454
rect 164486 183218 164528 183454
rect 164208 183134 164528 183218
rect 164208 182898 164250 183134
rect 164486 182898 164528 183134
rect 164208 182866 164528 182898
rect 164003 160444 164069 160445
rect 164003 160380 164004 160444
rect 164068 160380 164069 160444
rect 164003 160379 164069 160380
rect 164006 159901 164066 160379
rect 164742 159901 164802 232323
rect 165107 218924 165173 218925
rect 165107 218860 165108 218924
rect 165172 218860 165173 218924
rect 165107 218859 165173 218860
rect 164923 218652 164989 218653
rect 164923 218588 164924 218652
rect 164988 218588 164989 218652
rect 164923 218587 164989 218588
rect 163819 159900 163885 159901
rect 163819 159836 163820 159900
rect 163884 159836 163885 159900
rect 163819 159835 163885 159836
rect 164003 159900 164069 159901
rect 164003 159836 164004 159900
rect 164068 159836 164069 159900
rect 164003 159835 164069 159836
rect 164739 159900 164805 159901
rect 164739 159836 164740 159900
rect 164804 159836 164805 159900
rect 164739 159835 164805 159836
rect 163635 159764 163701 159765
rect 163635 159700 163636 159764
rect 163700 159700 163701 159764
rect 163635 159699 163701 159700
rect 164555 159764 164621 159765
rect 164555 159700 164556 159764
rect 164620 159700 164621 159764
rect 164555 159699 164621 159700
rect 163451 158676 163517 158677
rect 163451 158612 163452 158676
rect 163516 158612 163517 158676
rect 163451 158611 163517 158612
rect 164187 158676 164253 158677
rect 164187 158612 164188 158676
rect 164252 158612 164253 158676
rect 164187 158611 164253 158612
rect 162899 157180 162965 157181
rect 162899 157116 162900 157180
rect 162964 157116 162965 157180
rect 162899 157115 162965 157116
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 162902 146981 162962 157115
rect 162899 146980 162965 146981
rect 162899 146916 162900 146980
rect 162964 146916 162965 146980
rect 162899 146915 162965 146916
rect 164190 142170 164250 158611
rect 164558 157453 164618 159699
rect 164742 158677 164802 159835
rect 164739 158676 164805 158677
rect 164739 158612 164740 158676
rect 164804 158612 164805 158676
rect 164739 158611 164805 158612
rect 164926 158130 164986 218587
rect 165110 158405 165170 218859
rect 165478 159765 165538 233139
rect 165659 231164 165725 231165
rect 165659 231100 165660 231164
rect 165724 231100 165725 231164
rect 165659 231099 165725 231100
rect 165662 160037 165722 231099
rect 165659 160036 165725 160037
rect 165659 159972 165660 160036
rect 165724 159972 165725 160036
rect 165659 159971 165725 159972
rect 165475 159764 165541 159765
rect 165475 159700 165476 159764
rect 165540 159700 165541 159764
rect 165475 159699 165541 159700
rect 165662 158677 165722 159971
rect 165846 159901 165906 236675
rect 173755 236604 173821 236605
rect 173755 236540 173756 236604
rect 173820 236540 173821 236604
rect 173755 236539 173821 236540
rect 173571 233612 173637 233613
rect 173571 233548 173572 233612
rect 173636 233548 173637 233612
rect 173571 233547 173637 233548
rect 173019 233476 173085 233477
rect 173019 233412 173020 233476
rect 173084 233412 173085 233476
rect 173019 233411 173085 233412
rect 172283 231844 172349 231845
rect 172283 231780 172284 231844
rect 172348 231780 172349 231844
rect 172283 231779 172349 231780
rect 166395 231572 166461 231573
rect 166395 231508 166396 231572
rect 166460 231508 166461 231572
rect 166395 231507 166461 231508
rect 165843 159900 165909 159901
rect 165843 159836 165844 159900
rect 165908 159836 165909 159900
rect 165843 159835 165909 159836
rect 165291 158676 165357 158677
rect 165291 158612 165292 158676
rect 165356 158612 165357 158676
rect 165291 158611 165357 158612
rect 165659 158676 165725 158677
rect 165659 158612 165660 158676
rect 165724 158612 165725 158676
rect 165659 158611 165725 158612
rect 165107 158404 165173 158405
rect 165107 158340 165108 158404
rect 165172 158340 165173 158404
rect 165107 158339 165173 158340
rect 165294 158130 165354 158611
rect 164926 158070 165354 158130
rect 164555 157452 164621 157453
rect 164555 157388 164556 157452
rect 164620 157388 164621 157452
rect 164555 157387 164621 157388
rect 164371 157316 164437 157317
rect 164371 157252 164372 157316
rect 164436 157252 164437 157316
rect 164371 157251 164437 157252
rect 164374 144125 164434 157251
rect 164371 144124 164437 144125
rect 164371 144060 164372 144124
rect 164436 144060 164437 144124
rect 164371 144059 164437 144060
rect 164190 142110 164434 142170
rect 164374 130389 164434 142110
rect 164371 130388 164437 130389
rect 164371 130324 164372 130388
rect 164436 130324 164437 130388
rect 164371 130323 164437 130324
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 165846 113797 165906 159835
rect 166398 159765 166458 231507
rect 168235 231436 168301 231437
rect 168235 231372 168236 231436
rect 168300 231372 168301 231436
rect 168235 231371 168301 231372
rect 166579 231300 166645 231301
rect 166579 231236 166580 231300
rect 166644 231236 166645 231300
rect 166579 231235 166645 231236
rect 166582 159901 166642 231235
rect 168051 229804 168117 229805
rect 168051 229740 168052 229804
rect 168116 229740 168117 229804
rect 168051 229739 168117 229740
rect 167683 224364 167749 224365
rect 167683 224300 167684 224364
rect 167748 224300 167749 224364
rect 167683 224299 167749 224300
rect 166579 159900 166645 159901
rect 166579 159836 166580 159900
rect 166644 159836 166645 159900
rect 166579 159835 166645 159836
rect 166395 159764 166461 159765
rect 166395 159700 166396 159764
rect 166460 159700 166461 159764
rect 166395 159699 166461 159700
rect 167686 158677 167746 224299
rect 167867 218788 167933 218789
rect 167867 218724 167868 218788
rect 167932 218724 167933 218788
rect 167867 218723 167933 218724
rect 167870 159901 167930 218723
rect 168054 159901 168114 229739
rect 167867 159900 167933 159901
rect 167867 159836 167868 159900
rect 167932 159836 167933 159900
rect 167867 159835 167933 159836
rect 168051 159900 168117 159901
rect 168051 159836 168052 159900
rect 168116 159836 168117 159900
rect 168051 159835 168117 159836
rect 168238 159765 168298 231371
rect 168787 229940 168853 229941
rect 168787 229876 168788 229940
rect 168852 229876 168853 229940
rect 168787 229875 168853 229876
rect 168235 159764 168301 159765
rect 168235 159700 168236 159764
rect 168300 159700 168301 159764
rect 168235 159699 168301 159700
rect 168790 159629 168850 229875
rect 169339 224228 169405 224229
rect 169339 224164 169340 224228
rect 169404 224164 169405 224228
rect 169339 224163 169405 224164
rect 169155 220284 169221 220285
rect 169155 220220 169156 220284
rect 169220 220220 169221 220284
rect 169155 220219 169221 220220
rect 168971 217700 169037 217701
rect 168971 217636 168972 217700
rect 169036 217636 169037 217700
rect 168971 217635 169037 217636
rect 168974 159765 169034 217635
rect 169158 159901 169218 220219
rect 169342 160037 169402 224163
rect 170995 217836 171061 217837
rect 170995 217772 170996 217836
rect 171060 217772 171061 217836
rect 170995 217771 171061 217772
rect 170627 217428 170693 217429
rect 170627 217364 170628 217428
rect 170692 217364 170693 217428
rect 170627 217363 170693 217364
rect 170443 214572 170509 214573
rect 170443 214508 170444 214572
rect 170508 214508 170509 214572
rect 170443 214507 170509 214508
rect 169523 160716 169589 160717
rect 169523 160652 169524 160716
rect 169588 160652 169589 160716
rect 169523 160651 169589 160652
rect 169339 160036 169405 160037
rect 169339 159972 169340 160036
rect 169404 159972 169405 160036
rect 169339 159971 169405 159972
rect 169526 159901 169586 160651
rect 169155 159900 169221 159901
rect 169155 159836 169156 159900
rect 169220 159836 169221 159900
rect 169155 159835 169221 159836
rect 169523 159900 169589 159901
rect 169523 159836 169524 159900
rect 169588 159836 169589 159900
rect 169523 159835 169589 159836
rect 170259 159900 170325 159901
rect 170259 159836 170260 159900
rect 170324 159836 170325 159900
rect 170259 159835 170325 159836
rect 168971 159764 169037 159765
rect 168971 159700 168972 159764
rect 169036 159700 169037 159764
rect 168971 159699 169037 159700
rect 170075 159764 170141 159765
rect 170075 159700 170076 159764
rect 170140 159700 170141 159764
rect 170075 159699 170141 159700
rect 168787 159628 168853 159629
rect 168787 159564 168788 159628
rect 168852 159564 168853 159628
rect 168787 159563 168853 159564
rect 170078 158949 170138 159699
rect 170075 158948 170141 158949
rect 170075 158884 170076 158948
rect 170140 158884 170141 158948
rect 170075 158883 170141 158884
rect 170262 158677 170322 159835
rect 170446 159629 170506 214507
rect 170630 159765 170690 217363
rect 170811 217020 170877 217021
rect 170811 216956 170812 217020
rect 170876 216956 170877 217020
rect 170811 216955 170877 216956
rect 170814 159901 170874 216955
rect 170811 159900 170877 159901
rect 170811 159836 170812 159900
rect 170876 159836 170877 159900
rect 170811 159835 170877 159836
rect 170627 159764 170693 159765
rect 170627 159700 170628 159764
rect 170692 159700 170693 159764
rect 170627 159699 170693 159700
rect 170443 159628 170509 159629
rect 170443 159564 170444 159628
rect 170508 159564 170509 159628
rect 170443 159563 170509 159564
rect 170998 159357 171058 217771
rect 171731 217564 171797 217565
rect 171731 217500 171732 217564
rect 171796 217500 171797 217564
rect 171731 217499 171797 217500
rect 171363 160308 171429 160309
rect 171363 160244 171364 160308
rect 171428 160244 171429 160308
rect 171363 160243 171429 160244
rect 171179 159900 171245 159901
rect 171179 159836 171180 159900
rect 171244 159836 171245 159900
rect 171179 159835 171245 159836
rect 170995 159356 171061 159357
rect 170995 159292 170996 159356
rect 171060 159292 171061 159356
rect 170995 159291 171061 159292
rect 166027 158676 166093 158677
rect 166027 158612 166028 158676
rect 166092 158612 166093 158676
rect 166027 158611 166093 158612
rect 167683 158676 167749 158677
rect 167683 158612 167684 158676
rect 167748 158612 167749 158676
rect 167683 158611 167749 158612
rect 168419 158676 168485 158677
rect 168419 158612 168420 158676
rect 168484 158612 168485 158676
rect 168419 158611 168485 158612
rect 168971 158676 169037 158677
rect 168971 158612 168972 158676
rect 169036 158612 169037 158676
rect 168971 158611 169037 158612
rect 170259 158676 170325 158677
rect 170259 158612 170260 158676
rect 170324 158612 170325 158676
rect 170259 158611 170325 158612
rect 165843 113796 165909 113797
rect 165843 113732 165844 113796
rect 165908 113732 165909 113796
rect 165843 113731 165909 113732
rect 166030 112437 166090 158611
rect 168235 157860 168301 157861
rect 168235 157796 168236 157860
rect 168300 157796 168301 157860
rect 168235 157795 168301 157796
rect 167131 156772 167197 156773
rect 167131 156708 167132 156772
rect 167196 156708 167197 156772
rect 167131 156707 167197 156708
rect 167134 147690 167194 156707
rect 166950 147630 167194 147690
rect 166950 138685 167010 147630
rect 168238 138957 168298 157795
rect 168422 140725 168482 158611
rect 168603 158540 168669 158541
rect 168603 158476 168604 158540
rect 168668 158476 168669 158540
rect 168603 158475 168669 158476
rect 168606 146165 168666 158475
rect 168787 158404 168853 158405
rect 168787 158340 168788 158404
rect 168852 158340 168853 158404
rect 168787 158339 168853 158340
rect 168790 146301 168850 158339
rect 168974 147661 169034 158611
rect 171182 153210 171242 159835
rect 171366 159765 171426 160243
rect 171734 159901 171794 217499
rect 171915 217292 171981 217293
rect 171915 217228 171916 217292
rect 171980 217228 171981 217292
rect 171915 217227 171981 217228
rect 171547 159900 171613 159901
rect 171547 159836 171548 159900
rect 171612 159836 171613 159900
rect 171547 159835 171613 159836
rect 171731 159900 171797 159901
rect 171731 159836 171732 159900
rect 171796 159836 171797 159900
rect 171731 159835 171797 159836
rect 171363 159764 171429 159765
rect 171363 159700 171364 159764
rect 171428 159700 171429 159764
rect 171363 159699 171429 159700
rect 171550 158949 171610 159835
rect 171547 158948 171613 158949
rect 171547 158884 171548 158948
rect 171612 158884 171613 158948
rect 171547 158883 171613 158884
rect 171734 158677 171794 159835
rect 171918 159765 171978 217227
rect 172099 217156 172165 217157
rect 172099 217092 172100 217156
rect 172164 217092 172165 217156
rect 172099 217091 172165 217092
rect 171915 159764 171981 159765
rect 171915 159700 171916 159764
rect 171980 159700 171981 159764
rect 171915 159699 171981 159700
rect 171731 158676 171797 158677
rect 171731 158612 171732 158676
rect 171796 158612 171797 158676
rect 171731 158611 171797 158612
rect 171918 158541 171978 159699
rect 172102 159629 172162 217091
rect 172286 160309 172346 231779
rect 172283 160308 172349 160309
rect 172283 160244 172284 160308
rect 172348 160244 172349 160308
rect 172283 160243 172349 160244
rect 173022 159901 173082 233411
rect 173203 221508 173269 221509
rect 173203 221444 173204 221508
rect 173268 221444 173269 221508
rect 173203 221443 173269 221444
rect 173206 159901 173266 221443
rect 172651 159900 172717 159901
rect 172651 159836 172652 159900
rect 172716 159836 172717 159900
rect 172651 159835 172717 159836
rect 173019 159900 173085 159901
rect 173019 159836 173020 159900
rect 173084 159836 173085 159900
rect 173019 159835 173085 159836
rect 173203 159900 173269 159901
rect 173203 159836 173204 159900
rect 173268 159836 173269 159900
rect 173203 159835 173269 159836
rect 172099 159628 172165 159629
rect 172099 159564 172100 159628
rect 172164 159564 172165 159628
rect 172099 159563 172165 159564
rect 172102 158541 172162 159563
rect 172467 159220 172533 159221
rect 172467 159156 172468 159220
rect 172532 159156 172533 159220
rect 172467 159155 172533 159156
rect 172283 158676 172349 158677
rect 172283 158612 172284 158676
rect 172348 158612 172349 158676
rect 172283 158611 172349 158612
rect 171915 158540 171981 158541
rect 171915 158476 171916 158540
rect 171980 158476 171981 158540
rect 171915 158475 171981 158476
rect 172099 158540 172165 158541
rect 172099 158476 172100 158540
rect 172164 158476 172165 158540
rect 172099 158475 172165 158476
rect 170998 153150 171242 153210
rect 170998 148477 171058 153150
rect 170995 148476 171061 148477
rect 170995 148412 170996 148476
rect 171060 148412 171061 148476
rect 170995 148411 171061 148412
rect 170998 147690 171058 148411
rect 168971 147660 169037 147661
rect 168971 147596 168972 147660
rect 169036 147596 169037 147660
rect 168971 147595 169037 147596
rect 170262 147630 171058 147690
rect 168787 146300 168853 146301
rect 168787 146236 168788 146300
rect 168852 146236 168853 146300
rect 168787 146235 168853 146236
rect 168603 146164 168669 146165
rect 168603 146100 168604 146164
rect 168668 146100 168669 146164
rect 168603 146099 168669 146100
rect 170262 141405 170322 147630
rect 172286 142765 172346 158611
rect 172470 158133 172530 159155
rect 172654 158269 172714 159835
rect 173574 159765 173634 233547
rect 173758 159901 173818 236539
rect 174307 232796 174373 232797
rect 174307 232732 174308 232796
rect 174372 232732 174373 232796
rect 174307 232731 174373 232732
rect 174310 159901 174370 232731
rect 175043 232660 175109 232661
rect 175043 232596 175044 232660
rect 175108 232596 175109 232660
rect 175043 232595 175109 232596
rect 174675 231708 174741 231709
rect 174675 231644 174676 231708
rect 174740 231644 174741 231708
rect 174675 231643 174741 231644
rect 174491 213212 174557 213213
rect 174491 213148 174492 213212
rect 174556 213148 174557 213212
rect 174491 213147 174557 213148
rect 173755 159900 173821 159901
rect 173755 159836 173756 159900
rect 173820 159836 173821 159900
rect 173755 159835 173821 159836
rect 174307 159900 174373 159901
rect 174307 159836 174308 159900
rect 174372 159836 174373 159900
rect 174307 159835 174373 159836
rect 174494 159765 174554 213147
rect 174678 159901 174738 231643
rect 174675 159900 174741 159901
rect 174675 159836 174676 159900
rect 174740 159836 174741 159900
rect 174675 159835 174741 159836
rect 173571 159764 173637 159765
rect 173571 159700 173572 159764
rect 173636 159700 173637 159764
rect 173571 159699 173637 159700
rect 174491 159764 174557 159765
rect 174491 159700 174492 159764
rect 174556 159700 174557 159764
rect 174491 159699 174557 159700
rect 173203 158676 173269 158677
rect 173203 158612 173204 158676
rect 173268 158612 173269 158676
rect 173203 158611 173269 158612
rect 172651 158268 172717 158269
rect 172651 158204 172652 158268
rect 172716 158204 172717 158268
rect 172651 158203 172717 158204
rect 172467 158132 172533 158133
rect 172467 158068 172468 158132
rect 172532 158068 172533 158132
rect 172467 158067 172533 158068
rect 173019 157316 173085 157317
rect 173019 157252 173020 157316
rect 173084 157252 173085 157316
rect 173019 157251 173085 157252
rect 173022 143173 173082 157251
rect 173206 147117 173266 158611
rect 174678 158541 174738 159835
rect 175046 159629 175106 232595
rect 175227 159900 175293 159901
rect 175227 159836 175228 159900
rect 175292 159836 175293 159900
rect 175227 159835 175293 159836
rect 175043 159628 175109 159629
rect 175043 159564 175044 159628
rect 175108 159564 175109 159628
rect 175043 159563 175109 159564
rect 175043 158676 175109 158677
rect 175043 158612 175044 158676
rect 175108 158612 175109 158676
rect 175043 158611 175109 158612
rect 174675 158540 174741 158541
rect 174675 158476 174676 158540
rect 174740 158476 174741 158540
rect 174675 158475 174741 158476
rect 174307 158404 174373 158405
rect 174307 158340 174308 158404
rect 174372 158340 174373 158404
rect 174307 158339 174373 158340
rect 173387 147252 173453 147253
rect 173387 147188 173388 147252
rect 173452 147188 173453 147252
rect 173387 147187 173453 147188
rect 173203 147116 173269 147117
rect 173203 147052 173204 147116
rect 173268 147052 173269 147116
rect 173203 147051 173269 147052
rect 173019 143172 173085 143173
rect 173019 143108 173020 143172
rect 173084 143108 173085 143172
rect 173019 143107 173085 143108
rect 171731 142764 171797 142765
rect 171731 142700 171732 142764
rect 171796 142700 171797 142764
rect 171731 142699 171797 142700
rect 172283 142764 172349 142765
rect 172283 142700 172284 142764
rect 172348 142700 172349 142764
rect 172283 142699 172349 142700
rect 170259 141404 170325 141405
rect 170259 141340 170260 141404
rect 170324 141340 170325 141404
rect 170259 141339 170325 141340
rect 168419 140724 168485 140725
rect 168419 140660 168420 140724
rect 168484 140660 168485 140724
rect 168419 140659 168485 140660
rect 167131 138956 167197 138957
rect 167131 138892 167132 138956
rect 167196 138892 167197 138956
rect 167131 138891 167197 138892
rect 168235 138956 168301 138957
rect 168235 138892 168236 138956
rect 168300 138892 168301 138956
rect 168235 138891 168301 138892
rect 166947 138684 167013 138685
rect 166947 138620 166948 138684
rect 167012 138620 167013 138684
rect 166947 138619 167013 138620
rect 166211 137596 166277 137597
rect 166211 137532 166212 137596
rect 166276 137532 166277 137596
rect 166211 137531 166277 137532
rect 166214 131749 166274 137531
rect 167134 137325 167194 138891
rect 167131 137324 167197 137325
rect 167131 137260 167132 137324
rect 167196 137260 167197 137324
rect 167131 137259 167197 137260
rect 171734 134469 171794 142699
rect 171731 134468 171797 134469
rect 171731 134404 171732 134468
rect 171796 134404 171797 134468
rect 171731 134403 171797 134404
rect 166211 131748 166277 131749
rect 166211 131684 166212 131748
rect 166276 131684 166277 131748
rect 166211 131683 166277 131684
rect 166027 112436 166093 112437
rect 166027 112372 166028 112436
rect 166092 112372 166093 112436
rect 166027 112371 166093 112372
rect 173022 111077 173082 143107
rect 173206 126309 173266 147051
rect 173390 135965 173450 147187
rect 174310 143445 174370 158339
rect 175046 147690 175106 158611
rect 175230 158541 175290 159835
rect 175782 159493 175842 238035
rect 175963 237964 176029 237965
rect 175963 237900 175964 237964
rect 176028 237900 176029 237964
rect 175963 237899 176029 237900
rect 175966 160173 176026 237899
rect 177251 237692 177317 237693
rect 177251 237628 177252 237692
rect 177316 237628 177317 237692
rect 177251 237627 177317 237628
rect 176515 235380 176581 235381
rect 176515 235316 176516 235380
rect 176580 235316 176581 235380
rect 176515 235315 176581 235316
rect 176147 231028 176213 231029
rect 176147 230964 176148 231028
rect 176212 230964 176213 231028
rect 176147 230963 176213 230964
rect 175963 160172 176029 160173
rect 175963 160108 175964 160172
rect 176028 160108 176029 160172
rect 175963 160107 176029 160108
rect 175779 159492 175845 159493
rect 175779 159428 175780 159492
rect 175844 159428 175845 159492
rect 175779 159427 175845 159428
rect 175411 158676 175477 158677
rect 175411 158612 175412 158676
rect 175476 158612 175477 158676
rect 175411 158611 175477 158612
rect 175227 158540 175293 158541
rect 175227 158476 175228 158540
rect 175292 158476 175293 158540
rect 175227 158475 175293 158476
rect 175227 158268 175293 158269
rect 175227 158204 175228 158268
rect 175292 158204 175293 158268
rect 175227 158203 175293 158204
rect 174494 147630 175106 147690
rect 174494 147253 174554 147630
rect 174491 147252 174557 147253
rect 174491 147188 174492 147252
rect 174556 147188 174557 147252
rect 174491 147187 174557 147188
rect 174307 143444 174373 143445
rect 174307 143380 174308 143444
rect 174372 143380 174373 143444
rect 174307 143379 174373 143380
rect 174494 141541 174554 147187
rect 175230 146301 175290 158203
rect 175414 156909 175474 158611
rect 176150 157453 176210 230963
rect 176518 159901 176578 235315
rect 176515 159900 176581 159901
rect 176515 159836 176516 159900
rect 176580 159836 176581 159900
rect 176515 159835 176581 159836
rect 176331 159764 176397 159765
rect 176331 159700 176332 159764
rect 176396 159700 176397 159764
rect 176331 159699 176397 159700
rect 176334 158677 176394 159699
rect 177254 159493 177314 237627
rect 180379 234428 180445 234429
rect 180379 234364 180380 234428
rect 180444 234364 180445 234428
rect 180379 234363 180445 234364
rect 178539 220828 178605 220829
rect 178539 220764 178540 220828
rect 178604 220764 178605 220828
rect 178539 220763 178605 220764
rect 178542 159765 178602 220763
rect 179091 213892 179157 213893
rect 179091 213828 179092 213892
rect 179156 213828 179157 213892
rect 179091 213827 179157 213828
rect 178907 213756 178973 213757
rect 178907 213692 178908 213756
rect 178972 213692 178973 213756
rect 178907 213691 178973 213692
rect 178723 211852 178789 211853
rect 178723 211788 178724 211852
rect 178788 211788 178789 211852
rect 178723 211787 178789 211788
rect 178539 159764 178605 159765
rect 178539 159700 178540 159764
rect 178604 159700 178605 159764
rect 178539 159699 178605 159700
rect 177251 159492 177317 159493
rect 177251 159428 177252 159492
rect 177316 159428 177317 159492
rect 177251 159427 177317 159428
rect 178726 158677 178786 211787
rect 178910 159901 178970 213691
rect 178907 159900 178973 159901
rect 178907 159836 178908 159900
rect 178972 159836 178973 159900
rect 178907 159835 178973 159836
rect 176331 158676 176397 158677
rect 176331 158612 176332 158676
rect 176396 158612 176397 158676
rect 176331 158611 176397 158612
rect 178723 158676 178789 158677
rect 178723 158612 178724 158676
rect 178788 158612 178789 158676
rect 178723 158611 178789 158612
rect 176515 158540 176581 158541
rect 176515 158476 176516 158540
rect 176580 158476 176581 158540
rect 176515 158475 176581 158476
rect 176147 157452 176213 157453
rect 176147 157388 176148 157452
rect 176212 157388 176213 157452
rect 176147 157387 176213 157388
rect 175411 156908 175477 156909
rect 175411 156844 175412 156908
rect 175476 156844 175477 156908
rect 175411 156843 175477 156844
rect 175414 155957 175474 156843
rect 175411 155956 175477 155957
rect 175411 155892 175412 155956
rect 175476 155892 175477 155956
rect 175411 155891 175477 155892
rect 175227 146300 175293 146301
rect 175227 146236 175228 146300
rect 175292 146236 175293 146300
rect 175227 146235 175293 146236
rect 176518 145893 176578 158475
rect 177803 157860 177869 157861
rect 177803 157796 177804 157860
rect 177868 157796 177869 157860
rect 177803 157795 177869 157796
rect 177251 157724 177317 157725
rect 177251 157660 177252 157724
rect 177316 157660 177317 157724
rect 177251 157659 177317 157660
rect 176515 145892 176581 145893
rect 176515 145828 176516 145892
rect 176580 145828 176581 145892
rect 176515 145827 176581 145828
rect 176518 142170 176578 145827
rect 175782 142110 176578 142170
rect 174491 141540 174557 141541
rect 174491 141476 174492 141540
rect 174556 141476 174557 141540
rect 174491 141475 174557 141476
rect 173387 135964 173453 135965
rect 173387 135900 173388 135964
rect 173452 135900 173453 135964
rect 173387 135899 173453 135900
rect 175782 131205 175842 142110
rect 177254 140589 177314 157659
rect 177435 157452 177501 157453
rect 177435 157388 177436 157452
rect 177500 157388 177501 157452
rect 177435 157387 177501 157388
rect 177619 157452 177685 157453
rect 177619 157388 177620 157452
rect 177684 157388 177685 157452
rect 177619 157387 177685 157388
rect 177438 149973 177498 157387
rect 177622 150109 177682 157387
rect 177619 150108 177685 150109
rect 177619 150044 177620 150108
rect 177684 150044 177685 150108
rect 177619 150043 177685 150044
rect 177435 149972 177501 149973
rect 177435 149908 177436 149972
rect 177500 149908 177501 149972
rect 177435 149907 177501 149908
rect 177251 140588 177317 140589
rect 177251 140524 177252 140588
rect 177316 140524 177317 140588
rect 177251 140523 177317 140524
rect 175779 131204 175845 131205
rect 175779 131140 175780 131204
rect 175844 131140 175845 131204
rect 175779 131139 175845 131140
rect 173203 126308 173269 126309
rect 173203 126244 173204 126308
rect 173268 126244 173269 126308
rect 173203 126243 173269 126244
rect 173019 111076 173085 111077
rect 173019 111012 173020 111076
rect 173084 111012 173085 111076
rect 173019 111011 173085 111012
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 177254 24173 177314 140523
rect 177438 136645 177498 149907
rect 177435 136644 177501 136645
rect 177435 136580 177436 136644
rect 177500 136580 177501 136644
rect 177435 136579 177501 136580
rect 177622 120869 177682 150043
rect 177806 149837 177866 157795
rect 177803 149836 177869 149837
rect 177803 149772 177804 149836
rect 177868 149772 177869 149836
rect 177803 149771 177869 149772
rect 177806 138685 177866 149771
rect 178726 139909 178786 158611
rect 179094 157861 179154 213827
rect 180195 213484 180261 213485
rect 180195 213420 180196 213484
rect 180260 213420 180261 213484
rect 180195 213419 180261 213420
rect 180011 213076 180077 213077
rect 180011 213012 180012 213076
rect 180076 213012 180077 213076
rect 180011 213011 180077 213012
rect 179568 187174 179888 187206
rect 179568 186938 179610 187174
rect 179846 186938 179888 187174
rect 179568 186854 179888 186938
rect 179568 186618 179610 186854
rect 179846 186618 179888 186854
rect 179568 186586 179888 186618
rect 179275 157996 179341 157997
rect 179275 157932 179276 157996
rect 179340 157932 179341 157996
rect 179275 157931 179341 157932
rect 179091 157860 179157 157861
rect 179091 157796 179092 157860
rect 179156 157796 179157 157860
rect 179091 157795 179157 157796
rect 178907 157724 178973 157725
rect 178907 157660 178908 157724
rect 178972 157660 178973 157724
rect 178907 157659 178973 157660
rect 178910 144125 178970 157659
rect 179091 157452 179157 157453
rect 179091 157388 179092 157452
rect 179156 157388 179157 157452
rect 179091 157387 179157 157388
rect 179094 151333 179154 157387
rect 179278 155685 179338 157931
rect 180014 157725 180074 213011
rect 180198 158677 180258 213419
rect 180382 159901 180442 234363
rect 181483 234020 181549 234021
rect 181483 233956 181484 234020
rect 181548 233956 181549 234020
rect 181483 233955 181549 233956
rect 180563 233884 180629 233885
rect 180563 233820 180564 233884
rect 180628 233820 180629 233884
rect 180563 233819 180629 233820
rect 180566 159901 180626 233819
rect 181299 230076 181365 230077
rect 181299 230012 181300 230076
rect 181364 230012 181365 230076
rect 181299 230011 181365 230012
rect 181115 228580 181181 228581
rect 181115 228516 181116 228580
rect 181180 228516 181181 228580
rect 181115 228515 181181 228516
rect 180931 211988 180997 211989
rect 180931 211924 180932 211988
rect 180996 211924 180997 211988
rect 180931 211923 180997 211924
rect 180379 159900 180445 159901
rect 180379 159836 180380 159900
rect 180444 159836 180445 159900
rect 180379 159835 180445 159836
rect 180563 159900 180629 159901
rect 180563 159836 180564 159900
rect 180628 159836 180629 159900
rect 180563 159835 180629 159836
rect 180195 158676 180261 158677
rect 180195 158612 180196 158676
rect 180260 158612 180261 158676
rect 180195 158611 180261 158612
rect 180011 157724 180077 157725
rect 180011 157660 180012 157724
rect 180076 157660 180077 157724
rect 180011 157659 180077 157660
rect 180011 157452 180077 157453
rect 180011 157388 180012 157452
rect 180076 157388 180077 157452
rect 180011 157387 180077 157388
rect 179275 155684 179341 155685
rect 179275 155620 179276 155684
rect 179340 155620 179341 155684
rect 179275 155619 179341 155620
rect 179091 151332 179157 151333
rect 179091 151268 179092 151332
rect 179156 151268 179157 151332
rect 179091 151267 179157 151268
rect 178907 144124 178973 144125
rect 178907 144060 178908 144124
rect 178972 144060 178973 144124
rect 178907 144059 178973 144060
rect 178723 139908 178789 139909
rect 178723 139844 178724 139908
rect 178788 139844 178789 139908
rect 178723 139843 178789 139844
rect 177803 138684 177869 138685
rect 177803 138620 177804 138684
rect 177868 138620 177869 138684
rect 177803 138619 177869 138620
rect 177619 120868 177685 120869
rect 177619 120804 177620 120868
rect 177684 120804 177685 120868
rect 177619 120803 177685 120804
rect 179094 91765 179154 151267
rect 179091 91764 179157 91765
rect 179091 91700 179092 91764
rect 179156 91700 179157 91764
rect 179091 91699 179157 91700
rect 177251 24172 177317 24173
rect 177251 24108 177252 24172
rect 177316 24108 177317 24172
rect 177251 24107 177317 24108
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 179278 3637 179338 155619
rect 180014 146029 180074 157387
rect 180011 146028 180077 146029
rect 180011 145964 180012 146028
rect 180076 145964 180077 146028
rect 180011 145963 180077 145964
rect 180198 135965 180258 158611
rect 180195 135964 180261 135965
rect 180195 135900 180196 135964
rect 180260 135900 180261 135964
rect 180195 135899 180261 135900
rect 180382 130389 180442 159835
rect 180934 159765 180994 211923
rect 180931 159764 180997 159765
rect 180931 159700 180932 159764
rect 180996 159700 180997 159764
rect 180931 159699 180997 159700
rect 181118 159629 181178 228515
rect 181115 159628 181181 159629
rect 181115 159564 181116 159628
rect 181180 159564 181181 159628
rect 181115 159563 181181 159564
rect 181302 158677 181362 230011
rect 181486 159901 181546 233955
rect 181794 219454 182414 254898
rect 185514 705798 186134 705830
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 184427 234292 184493 234293
rect 184427 234228 184428 234292
rect 184492 234228 184493 234292
rect 184427 234227 184493 234228
rect 182587 233748 182653 233749
rect 182587 233684 182588 233748
rect 182652 233684 182653 233748
rect 182587 233683 182653 233684
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181483 159900 181549 159901
rect 181483 159836 181484 159900
rect 181548 159836 181549 159900
rect 181483 159835 181549 159836
rect 181299 158676 181365 158677
rect 181299 158612 181300 158676
rect 181364 158612 181365 158676
rect 181299 158611 181365 158612
rect 181115 157724 181181 157725
rect 181115 157660 181116 157724
rect 181180 157660 181181 157724
rect 181115 157659 181181 157660
rect 180563 157452 180629 157453
rect 180563 157388 180564 157452
rect 180628 157388 180629 157452
rect 180563 157387 180629 157388
rect 180379 130388 180445 130389
rect 180379 130324 180380 130388
rect 180444 130324 180445 130388
rect 180379 130323 180445 130324
rect 180566 124133 180626 157387
rect 181118 126989 181178 157659
rect 181115 126988 181181 126989
rect 181115 126924 181116 126988
rect 181180 126924 181181 126988
rect 181115 126923 181181 126924
rect 180563 124132 180629 124133
rect 180563 124068 180564 124132
rect 180628 124068 180629 124132
rect 180563 124067 180629 124068
rect 181302 98837 181362 158611
rect 181483 157452 181549 157453
rect 181483 157388 181484 157452
rect 181548 157388 181549 157452
rect 181483 157387 181549 157388
rect 181486 140725 181546 157387
rect 181794 147454 182414 182898
rect 182590 159901 182650 233683
rect 183139 226948 183205 226949
rect 183139 226884 183140 226948
rect 183204 226884 183205 226948
rect 183139 226883 183205 226884
rect 182955 219060 183021 219061
rect 182955 218996 182956 219060
rect 183020 218996 183021 219060
rect 182955 218995 183021 218996
rect 182771 213348 182837 213349
rect 182771 213284 182772 213348
rect 182836 213284 182837 213348
rect 182771 213283 182837 213284
rect 182587 159900 182653 159901
rect 182587 159836 182588 159900
rect 182652 159836 182653 159900
rect 182587 159835 182653 159836
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181483 140724 181549 140725
rect 181483 140660 181484 140724
rect 181548 140660 181549 140724
rect 181483 140659 181549 140660
rect 181486 112437 181546 140659
rect 181483 112436 181549 112437
rect 181483 112372 181484 112436
rect 181548 112372 181549 112436
rect 181483 112371 181549 112372
rect 181794 111454 182414 146898
rect 182590 124813 182650 159835
rect 182774 159765 182834 213283
rect 182771 159764 182837 159765
rect 182771 159700 182772 159764
rect 182836 159700 182837 159764
rect 182771 159699 182837 159700
rect 182587 124812 182653 124813
rect 182587 124748 182588 124812
rect 182652 124748 182653 124812
rect 182587 124747 182653 124748
rect 182774 122229 182834 159699
rect 182958 158677 183018 218995
rect 183142 159901 183202 226883
rect 184059 209540 184125 209541
rect 184059 209476 184060 209540
rect 184124 209476 184125 209540
rect 184059 209475 184125 209476
rect 184062 159901 184122 209475
rect 183139 159900 183205 159901
rect 183139 159836 183140 159900
rect 183204 159836 183205 159900
rect 183139 159835 183205 159836
rect 184059 159900 184125 159901
rect 184059 159836 184060 159900
rect 184124 159836 184125 159900
rect 184059 159835 184125 159836
rect 182955 158676 183021 158677
rect 182955 158612 182956 158676
rect 183020 158612 183021 158676
rect 182955 158611 183021 158612
rect 182958 127669 183018 158611
rect 182955 127668 183021 127669
rect 182955 127604 182956 127668
rect 183020 127604 183021 127668
rect 182955 127603 183021 127604
rect 182771 122228 182837 122229
rect 182771 122164 182772 122228
rect 182836 122164 182837 122228
rect 182771 122163 182837 122164
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181299 98836 181365 98837
rect 181299 98772 181300 98836
rect 181364 98772 181365 98836
rect 181299 98771 181365 98772
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 179275 3636 179341 3637
rect 179275 3572 179276 3636
rect 179340 3572 179341 3636
rect 179275 3571 179341 3572
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -1894 150134 -1862
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 184062 3365 184122 159835
rect 184430 159765 184490 234227
rect 184611 230212 184677 230213
rect 184611 230148 184612 230212
rect 184676 230148 184677 230212
rect 184611 230147 184677 230148
rect 184614 159901 184674 230147
rect 185514 223174 186134 258618
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 221514 705798 222134 705830
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 220675 373420 220741 373421
rect 220675 373356 220676 373420
rect 220740 373356 220741 373420
rect 220675 373355 220741 373356
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 220123 291548 220189 291549
rect 220123 291484 220124 291548
rect 220188 291484 220189 291548
rect 220123 291483 220189 291484
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 219939 291412 220005 291413
rect 219939 291348 219940 291412
rect 220004 291348 220005 291412
rect 219939 291347 220005 291348
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 188291 238508 188357 238509
rect 188291 238444 188292 238508
rect 188356 238444 188357 238508
rect 188291 238443 188357 238444
rect 186819 238236 186885 238237
rect 186819 238172 186820 238236
rect 186884 238172 186885 238236
rect 186819 238171 186885 238172
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185163 213620 185229 213621
rect 185163 213556 185164 213620
rect 185228 213556 185229 213620
rect 185163 213555 185229 213556
rect 185166 159901 185226 213555
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 184611 159900 184677 159901
rect 184611 159836 184612 159900
rect 184676 159836 184677 159900
rect 184611 159835 184677 159836
rect 185163 159900 185229 159901
rect 185163 159836 185164 159900
rect 185228 159836 185229 159900
rect 185163 159835 185229 159836
rect 184427 159764 184493 159765
rect 184427 159700 184428 159764
rect 184492 159700 184493 159764
rect 184427 159699 184493 159700
rect 184243 157452 184309 157453
rect 184243 157388 184244 157452
rect 184308 157388 184309 157452
rect 184243 157387 184309 157388
rect 184246 146301 184306 157387
rect 184243 146300 184309 146301
rect 184243 146236 184244 146300
rect 184308 146236 184309 146300
rect 184243 146235 184309 146236
rect 184246 3501 184306 146235
rect 184430 6085 184490 159699
rect 184614 6901 184674 159835
rect 184979 157452 185045 157453
rect 184979 157388 184980 157452
rect 185044 157388 185045 157452
rect 184979 157387 185045 157388
rect 184982 139773 185042 157387
rect 184979 139772 185045 139773
rect 184979 139708 184980 139772
rect 185044 139708 185045 139772
rect 184979 139707 185045 139708
rect 184611 6900 184677 6901
rect 184611 6836 184612 6900
rect 184676 6836 184677 6900
rect 184611 6835 184677 6836
rect 184982 6765 185042 139707
rect 184979 6764 185045 6765
rect 184979 6700 184980 6764
rect 185044 6700 185045 6764
rect 184979 6699 185045 6700
rect 185166 6629 185226 159835
rect 185514 151174 186134 186618
rect 186822 160717 186882 238171
rect 186819 160716 186885 160717
rect 186819 160652 186820 160716
rect 186884 160652 186885 160716
rect 186819 160651 186885 160652
rect 188294 158813 188354 238443
rect 191603 232932 191669 232933
rect 191603 232868 191604 232932
rect 191668 232868 191669 232932
rect 191603 232867 191669 232868
rect 188843 225588 188909 225589
rect 188843 225524 188844 225588
rect 188908 225524 188909 225588
rect 188843 225523 188909 225524
rect 188846 159901 188906 225523
rect 190315 210356 190381 210357
rect 190315 210292 190316 210356
rect 190380 210292 190381 210356
rect 190315 210291 190381 210292
rect 189579 209540 189645 209541
rect 189579 209476 189580 209540
rect 189644 209476 189645 209540
rect 189579 209475 189645 209476
rect 189582 208997 189642 209475
rect 189579 208996 189645 208997
rect 189579 208932 189580 208996
rect 189644 208932 189645 208996
rect 189579 208931 189645 208932
rect 190318 159901 190378 210291
rect 188475 159900 188541 159901
rect 188475 159836 188476 159900
rect 188540 159836 188541 159900
rect 188475 159835 188541 159836
rect 188843 159900 188909 159901
rect 188843 159836 188844 159900
rect 188908 159836 188909 159900
rect 188843 159835 188909 159836
rect 190315 159900 190381 159901
rect 190315 159836 190316 159900
rect 190380 159836 190381 159900
rect 190315 159835 190381 159836
rect 188291 158812 188357 158813
rect 188291 158748 188292 158812
rect 188356 158748 188357 158812
rect 188291 158747 188357 158748
rect 187003 158676 187069 158677
rect 187003 158612 187004 158676
rect 187068 158612 187069 158676
rect 187003 158611 187069 158612
rect 187187 158676 187253 158677
rect 187187 158612 187188 158676
rect 187252 158612 187253 158676
rect 187187 158611 187253 158612
rect 187555 158676 187621 158677
rect 187555 158612 187556 158676
rect 187620 158612 187621 158676
rect 187555 158611 187621 158612
rect 188291 158676 188357 158677
rect 188291 158612 188292 158676
rect 188356 158612 188357 158676
rect 188291 158611 188357 158612
rect 187006 153645 187066 158611
rect 187003 153644 187069 153645
rect 187003 153580 187004 153644
rect 187068 153580 187069 153644
rect 187003 153579 187069 153580
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 187190 141677 187250 158611
rect 187371 158540 187437 158541
rect 187371 158476 187372 158540
rect 187436 158476 187437 158540
rect 187371 158475 187437 158476
rect 187374 146981 187434 158475
rect 187371 146980 187437 146981
rect 187371 146916 187372 146980
rect 187436 146916 187437 146980
rect 187371 146915 187437 146916
rect 187187 141676 187253 141677
rect 187187 141612 187188 141676
rect 187252 141612 187253 141676
rect 187187 141611 187253 141612
rect 187190 119509 187250 141611
rect 187187 119508 187253 119509
rect 187187 119444 187188 119508
rect 187252 119444 187253 119508
rect 187187 119443 187253 119444
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 187374 105501 187434 146915
rect 187558 141813 187618 158611
rect 187555 141812 187621 141813
rect 187555 141748 187556 141812
rect 187620 141748 187621 141812
rect 187555 141747 187621 141748
rect 187371 105500 187437 105501
rect 187371 105436 187372 105500
rect 187436 105436 187437 105500
rect 187371 105435 187437 105436
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 187558 68237 187618 141747
rect 188294 140045 188354 158611
rect 188291 140044 188357 140045
rect 188291 139980 188292 140044
rect 188356 139980 188357 140044
rect 188291 139979 188357 139980
rect 188294 113933 188354 139979
rect 188291 113932 188357 113933
rect 188291 113868 188292 113932
rect 188356 113868 188357 113932
rect 188291 113867 188357 113868
rect 188478 102781 188538 159835
rect 190318 159490 190378 159835
rect 191606 159765 191666 232867
rect 193075 232524 193141 232525
rect 193075 232460 193076 232524
rect 193140 232460 193141 232524
rect 193075 232459 193141 232460
rect 193078 159901 193138 232459
rect 194363 231980 194429 231981
rect 194363 231916 194364 231980
rect 194428 231916 194429 231980
rect 194363 231915 194429 231916
rect 193811 209540 193877 209541
rect 193811 209476 193812 209540
rect 193876 209476 193877 209540
rect 193811 209475 193877 209476
rect 193814 167010 193874 209475
rect 193630 166950 193874 167010
rect 193630 159901 193690 166950
rect 194366 159901 194426 231915
rect 197123 225724 197189 225725
rect 197123 225660 197124 225724
rect 197188 225660 197189 225724
rect 197123 225659 197189 225660
rect 196939 214980 197005 214981
rect 196939 214916 196940 214980
rect 197004 214916 197005 214980
rect 196939 214915 197005 214916
rect 195651 214844 195717 214845
rect 195651 214780 195652 214844
rect 195716 214780 195717 214844
rect 195651 214779 195717 214780
rect 195467 209540 195533 209541
rect 195467 209476 195468 209540
rect 195532 209476 195533 209540
rect 195467 209475 195533 209476
rect 194928 183454 195248 183486
rect 194928 183218 194970 183454
rect 195206 183218 195248 183454
rect 194928 183134 195248 183218
rect 194928 182898 194970 183134
rect 195206 182898 195248 183134
rect 194928 182866 195248 182898
rect 195470 160850 195530 209475
rect 195286 160790 195530 160850
rect 195286 159901 195346 160790
rect 193075 159900 193141 159901
rect 193075 159836 193076 159900
rect 193140 159836 193141 159900
rect 193075 159835 193141 159836
rect 193627 159900 193693 159901
rect 193627 159836 193628 159900
rect 193692 159836 193693 159900
rect 193627 159835 193693 159836
rect 194363 159900 194429 159901
rect 194363 159836 194364 159900
rect 194428 159836 194429 159900
rect 194363 159835 194429 159836
rect 195283 159900 195349 159901
rect 195283 159836 195284 159900
rect 195348 159836 195349 159900
rect 195283 159835 195349 159836
rect 191603 159764 191669 159765
rect 191603 159700 191604 159764
rect 191668 159700 191669 159764
rect 191603 159699 191669 159700
rect 190134 159430 190378 159490
rect 188659 158676 188725 158677
rect 188659 158612 188660 158676
rect 188724 158612 188725 158676
rect 188659 158611 188725 158612
rect 188843 158676 188909 158677
rect 188843 158612 188844 158676
rect 188908 158612 188909 158676
rect 188843 158611 188909 158612
rect 189579 158676 189645 158677
rect 189579 158612 189580 158676
rect 189644 158612 189645 158676
rect 189579 158611 189645 158612
rect 189947 158676 190013 158677
rect 189947 158612 189948 158676
rect 190012 158612 190013 158676
rect 189947 158611 190013 158612
rect 188662 141405 188722 158611
rect 188846 141949 188906 158611
rect 189582 147690 189642 158611
rect 189582 147630 189826 147690
rect 188843 141948 188909 141949
rect 188843 141884 188844 141948
rect 188908 141884 188909 141948
rect 188843 141883 188909 141884
rect 188659 141404 188725 141405
rect 188659 141340 188660 141404
rect 188724 141340 188725 141404
rect 188659 141339 188725 141340
rect 188475 102780 188541 102781
rect 188475 102716 188476 102780
rect 188540 102716 188541 102780
rect 188475 102715 188541 102716
rect 187555 68236 187621 68237
rect 187555 68172 187556 68236
rect 187620 68172 187621 68236
rect 187555 68171 187621 68172
rect 188662 66877 188722 141339
rect 188659 66876 188725 66877
rect 188659 66812 188660 66876
rect 188724 66812 188725 66876
rect 188659 66811 188725 66812
rect 188846 65517 188906 141883
rect 189766 140453 189826 147630
rect 189950 142629 190010 158611
rect 189947 142628 190013 142629
rect 189947 142564 189948 142628
rect 190012 142564 190013 142628
rect 189947 142563 190013 142564
rect 189763 140452 189829 140453
rect 189763 140388 189764 140452
rect 189828 140388 189829 140452
rect 189763 140387 189829 140388
rect 189766 115293 189826 140387
rect 189763 115292 189829 115293
rect 189763 115228 189764 115292
rect 189828 115228 189829 115292
rect 189763 115227 189829 115228
rect 188843 65516 188909 65517
rect 188843 65452 188844 65516
rect 188908 65452 188909 65516
rect 188843 65451 188909 65452
rect 189950 62797 190010 142563
rect 190134 64157 190194 159430
rect 192523 159084 192589 159085
rect 192523 159020 192524 159084
rect 192588 159020 192589 159084
rect 192523 159019 192589 159020
rect 190315 158676 190381 158677
rect 190315 158612 190316 158676
rect 190380 158612 190381 158676
rect 190315 158611 190381 158612
rect 191235 158676 191301 158677
rect 191235 158612 191236 158676
rect 191300 158612 191301 158676
rect 191235 158611 191301 158612
rect 190318 141269 190378 158611
rect 191051 158540 191117 158541
rect 191051 158476 191052 158540
rect 191116 158476 191117 158540
rect 191051 158475 191117 158476
rect 190315 141268 190381 141269
rect 190315 141204 190316 141268
rect 190380 141204 190381 141268
rect 190315 141203 190381 141204
rect 190131 64156 190197 64157
rect 190131 64092 190132 64156
rect 190196 64092 190197 64156
rect 190131 64091 190197 64092
rect 189947 62796 190013 62797
rect 189947 62732 189948 62796
rect 190012 62732 190013 62796
rect 189947 62731 190013 62732
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 190318 40629 190378 141203
rect 191054 140861 191114 158475
rect 191238 144261 191298 158611
rect 191787 158404 191853 158405
rect 191787 158340 191788 158404
rect 191852 158340 191853 158404
rect 191787 158339 191853 158340
rect 191419 157316 191485 157317
rect 191419 157252 191420 157316
rect 191484 157252 191485 157316
rect 191419 157251 191485 157252
rect 191235 144260 191301 144261
rect 191235 144196 191236 144260
rect 191300 144196 191301 144260
rect 191235 144195 191301 144196
rect 191422 141541 191482 157251
rect 191790 144397 191850 158339
rect 191787 144396 191853 144397
rect 191787 144332 191788 144396
rect 191852 144332 191853 144396
rect 191787 144331 191853 144332
rect 191790 142170 191850 144331
rect 191606 142110 191850 142170
rect 191419 141540 191485 141541
rect 191419 141476 191420 141540
rect 191484 141476 191485 141540
rect 191419 141475 191485 141476
rect 191051 140860 191117 140861
rect 191051 140796 191052 140860
rect 191116 140796 191117 140860
rect 191051 140795 191117 140796
rect 190315 40628 190381 40629
rect 190315 40564 190316 40628
rect 190380 40564 190381 40628
rect 190315 40563 190381 40564
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185163 6628 185229 6629
rect 185163 6564 185164 6628
rect 185228 6564 185229 6628
rect 185163 6563 185229 6564
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 184427 6084 184493 6085
rect 184427 6020 184428 6084
rect 184492 6020 184493 6084
rect 184427 6019 184493 6020
rect 184243 3500 184309 3501
rect 184243 3436 184244 3500
rect 184308 3436 184309 3500
rect 184243 3435 184309 3436
rect 184059 3364 184125 3365
rect 184059 3300 184060 3364
rect 184124 3300 184125 3364
rect 184059 3299 184125 3300
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 -1306 186134 6618
rect 191422 6357 191482 141475
rect 191606 6493 191666 142110
rect 192526 137461 192586 159019
rect 193075 158676 193141 158677
rect 193075 158612 193076 158676
rect 193140 158612 193141 158676
rect 193075 158611 193141 158612
rect 192891 158540 192957 158541
rect 192891 158476 192892 158540
rect 192956 158476 192957 158540
rect 192891 158475 192957 158476
rect 192707 158268 192773 158269
rect 192707 158204 192708 158268
rect 192772 158204 192773 158268
rect 192707 158203 192773 158204
rect 192710 137597 192770 158203
rect 192707 137596 192773 137597
rect 192707 137532 192708 137596
rect 192772 137532 192773 137596
rect 192707 137531 192773 137532
rect 192523 137460 192589 137461
rect 192523 137396 192524 137460
rect 192588 137396 192589 137460
rect 192523 137395 192589 137396
rect 192526 9213 192586 137395
rect 192710 9485 192770 137531
rect 192894 137189 192954 158475
rect 193078 137733 193138 158611
rect 193630 158405 193690 159835
rect 195286 159490 195346 159835
rect 195654 159765 195714 214779
rect 195835 214708 195901 214709
rect 195835 214644 195836 214708
rect 195900 214644 195901 214708
rect 195835 214643 195901 214644
rect 195838 159901 195898 214643
rect 195835 159900 195901 159901
rect 195835 159836 195836 159900
rect 195900 159836 195901 159900
rect 195835 159835 195901 159836
rect 196942 159765 197002 214915
rect 197126 159901 197186 225659
rect 217794 219454 218414 254898
rect 219942 242181 220002 291347
rect 220126 272509 220186 291483
rect 220678 290325 220738 373355
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 236499 318476 236565 318477
rect 236499 318412 236500 318476
rect 236564 318412 236565 318476
rect 236499 318411 236565 318412
rect 223251 317116 223317 317117
rect 223251 317052 223252 317116
rect 223316 317052 223317 317116
rect 223251 317051 223317 317052
rect 222699 316028 222765 316029
rect 222699 315964 222700 316028
rect 222764 315964 222765 316028
rect 222699 315963 222765 315964
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221227 291276 221293 291277
rect 221227 291212 221228 291276
rect 221292 291212 221293 291276
rect 221227 291211 221293 291212
rect 220675 290324 220741 290325
rect 220675 290260 220676 290324
rect 220740 290260 220741 290324
rect 220675 290259 220741 290260
rect 221230 282165 221290 291211
rect 221227 282164 221293 282165
rect 221227 282100 221228 282164
rect 221292 282100 221293 282164
rect 221227 282099 221293 282100
rect 220123 272508 220189 272509
rect 220123 272444 220124 272508
rect 220188 272444 220189 272508
rect 220123 272443 220189 272444
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 219939 242180 220005 242181
rect 219939 242116 219940 242180
rect 220004 242116 220005 242180
rect 219939 242115 220005 242116
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 203195 212124 203261 212125
rect 203195 212060 203196 212124
rect 203260 212060 203261 212124
rect 203195 212059 203261 212060
rect 198411 210492 198477 210493
rect 198411 210428 198412 210492
rect 198476 210428 198477 210492
rect 198411 210427 198477 210428
rect 198043 210084 198109 210085
rect 198043 210020 198044 210084
rect 198108 210020 198109 210084
rect 198043 210019 198109 210020
rect 197859 209540 197925 209541
rect 197859 209476 197860 209540
rect 197924 209476 197925 209540
rect 197859 209475 197925 209476
rect 197862 159901 197922 209475
rect 198046 167010 198106 210019
rect 198046 166950 198290 167010
rect 198043 160988 198109 160989
rect 198043 160924 198044 160988
rect 198108 160924 198109 160988
rect 198043 160923 198109 160924
rect 197123 159900 197189 159901
rect 197123 159836 197124 159900
rect 197188 159836 197189 159900
rect 197123 159835 197189 159836
rect 197859 159900 197925 159901
rect 197859 159836 197860 159900
rect 197924 159836 197925 159900
rect 197859 159835 197925 159836
rect 195651 159764 195717 159765
rect 195651 159700 195652 159764
rect 195716 159700 195717 159764
rect 195651 159699 195717 159700
rect 196387 159764 196453 159765
rect 196387 159700 196388 159764
rect 196452 159700 196453 159764
rect 196387 159699 196453 159700
rect 196939 159764 197005 159765
rect 196939 159700 196940 159764
rect 197004 159700 197005 159764
rect 196939 159699 197005 159700
rect 195102 159430 195346 159490
rect 194179 158676 194245 158677
rect 194179 158612 194180 158676
rect 194244 158612 194245 158676
rect 194179 158611 194245 158612
rect 194363 158676 194429 158677
rect 194363 158612 194364 158676
rect 194428 158612 194429 158676
rect 194363 158611 194429 158612
rect 193995 158540 194061 158541
rect 193995 158476 193996 158540
rect 194060 158476 194061 158540
rect 193995 158475 194061 158476
rect 193627 158404 193693 158405
rect 193627 158340 193628 158404
rect 193692 158340 193693 158404
rect 193627 158339 193693 158340
rect 193998 152421 194058 158475
rect 193995 152420 194061 152421
rect 193995 152356 193996 152420
rect 194060 152356 194061 152420
rect 193995 152355 194061 152356
rect 193075 137732 193141 137733
rect 193075 137668 193076 137732
rect 193140 137668 193141 137732
rect 193075 137667 193141 137668
rect 192891 137188 192957 137189
rect 192891 137124 192892 137188
rect 192956 137124 192957 137188
rect 192891 137123 192957 137124
rect 192707 9484 192773 9485
rect 192707 9420 192708 9484
rect 192772 9420 192773 9484
rect 192707 9419 192773 9420
rect 192894 9349 192954 137123
rect 192891 9348 192957 9349
rect 192891 9284 192892 9348
rect 192956 9284 192957 9348
rect 192891 9283 192957 9284
rect 192523 9212 192589 9213
rect 192523 9148 192524 9212
rect 192588 9148 192589 9212
rect 192523 9147 192589 9148
rect 191603 6492 191669 6493
rect 191603 6428 191604 6492
rect 191668 6428 191669 6492
rect 191603 6427 191669 6428
rect 191419 6356 191485 6357
rect 191419 6292 191420 6356
rect 191484 6292 191485 6356
rect 191419 6291 191485 6292
rect 193078 6221 193138 137667
rect 193998 122093 194058 152355
rect 194182 137869 194242 158611
rect 194179 137868 194245 137869
rect 194179 137804 194180 137868
rect 194244 137804 194245 137868
rect 194179 137803 194245 137804
rect 193995 122092 194061 122093
rect 193995 122028 193996 122092
rect 194060 122028 194061 122092
rect 193995 122027 194061 122028
rect 194182 54501 194242 137803
rect 194366 137325 194426 158611
rect 194547 158268 194613 158269
rect 194547 158204 194548 158268
rect 194612 158204 194613 158268
rect 194547 158203 194613 158204
rect 194550 152693 194610 158203
rect 194547 152692 194613 152693
rect 194547 152628 194548 152692
rect 194612 152628 194613 152692
rect 194547 152627 194613 152628
rect 194363 137324 194429 137325
rect 194363 137260 194364 137324
rect 194428 137260 194429 137324
rect 194363 137259 194429 137260
rect 194179 54500 194245 54501
rect 194179 54436 194180 54500
rect 194244 54436 194245 54500
rect 194179 54435 194245 54436
rect 194366 51781 194426 137259
rect 194363 51780 194429 51781
rect 194363 51716 194364 51780
rect 194428 51716 194429 51780
rect 194363 51715 194429 51716
rect 195102 8941 195162 159430
rect 195283 158676 195349 158677
rect 195283 158612 195284 158676
rect 195348 158612 195349 158676
rect 195283 158611 195349 158612
rect 195286 152285 195346 158611
rect 195467 158540 195533 158541
rect 195467 158476 195468 158540
rect 195532 158476 195533 158540
rect 195467 158475 195533 158476
rect 195470 152965 195530 158475
rect 195651 158404 195717 158405
rect 195651 158340 195652 158404
rect 195716 158340 195717 158404
rect 195651 158339 195717 158340
rect 195467 152964 195533 152965
rect 195467 152900 195468 152964
rect 195532 152900 195533 152964
rect 195467 152899 195533 152900
rect 195283 152284 195349 152285
rect 195283 152220 195284 152284
rect 195348 152220 195349 152284
rect 195283 152219 195349 152220
rect 195286 120733 195346 152219
rect 195283 120732 195349 120733
rect 195283 120668 195284 120732
rect 195348 120668 195349 120732
rect 195283 120667 195349 120668
rect 195470 30973 195530 152899
rect 195654 139229 195714 158339
rect 196390 153237 196450 159699
rect 196755 158676 196821 158677
rect 196755 158612 196756 158676
rect 196820 158612 196821 158676
rect 196755 158611 196821 158612
rect 196939 158676 197005 158677
rect 196939 158612 196940 158676
rect 197004 158612 197005 158676
rect 196939 158611 197005 158612
rect 196387 153236 196453 153237
rect 196387 153172 196388 153236
rect 196452 153172 196453 153236
rect 196387 153171 196453 153172
rect 196758 150245 196818 158611
rect 196942 153101 197002 158611
rect 196939 153100 197005 153101
rect 196939 153036 196940 153100
rect 197004 153036 197005 153100
rect 196939 153035 197005 153036
rect 196755 150244 196821 150245
rect 196755 150180 196756 150244
rect 196820 150180 196821 150244
rect 196755 150179 196821 150180
rect 195651 139228 195717 139229
rect 195651 139164 195652 139228
rect 195716 139164 195717 139228
rect 195651 139163 195717 139164
rect 195467 30972 195533 30973
rect 195467 30908 195468 30972
rect 195532 30908 195533 30972
rect 195467 30907 195533 30908
rect 195654 9077 195714 139163
rect 196942 118013 197002 153035
rect 196939 118012 197005 118013
rect 196939 117948 196940 118012
rect 197004 117948 197005 118012
rect 196939 117947 197005 117948
rect 197126 11661 197186 159835
rect 197862 46205 197922 159835
rect 198046 159629 198106 160923
rect 198230 159901 198290 166950
rect 198227 159900 198293 159901
rect 198227 159836 198228 159900
rect 198292 159836 198293 159900
rect 198227 159835 198293 159836
rect 198414 159765 198474 210427
rect 199331 209812 199397 209813
rect 199331 209748 199332 209812
rect 199396 209748 199397 209812
rect 199331 209747 199397 209748
rect 199147 209540 199213 209541
rect 199147 209476 199148 209540
rect 199212 209476 199213 209540
rect 199147 209475 199213 209476
rect 198779 161124 198845 161125
rect 198779 161060 198780 161124
rect 198844 161060 198845 161124
rect 198779 161059 198845 161060
rect 198782 160173 198842 161059
rect 198779 160172 198845 160173
rect 198779 160108 198780 160172
rect 198844 160108 198845 160172
rect 198779 160107 198845 160108
rect 199150 159901 199210 209475
rect 199147 159900 199213 159901
rect 199147 159836 199148 159900
rect 199212 159836 199213 159900
rect 199147 159835 199213 159836
rect 199334 159765 199394 209747
rect 199883 209540 199949 209541
rect 199883 209476 199884 209540
rect 199948 209476 199949 209540
rect 199883 209475 199949 209476
rect 199886 159901 199946 209475
rect 201355 207636 201421 207637
rect 201355 207572 201356 207636
rect 201420 207572 201421 207636
rect 201355 207571 201421 207572
rect 201358 159901 201418 207571
rect 203198 206277 203258 212059
rect 203195 206276 203261 206277
rect 203195 206212 203196 206276
rect 203260 206212 203261 206276
rect 203195 206211 203261 206212
rect 208899 204916 208965 204917
rect 208899 204852 208900 204916
rect 208964 204852 208965 204916
rect 208899 204851 208965 204852
rect 207795 182884 207861 182885
rect 207795 182820 207796 182884
rect 207860 182820 207861 182884
rect 207795 182819 207861 182820
rect 205771 180028 205837 180029
rect 205771 179964 205772 180028
rect 205836 179964 205837 180028
rect 205771 179963 205837 179964
rect 204851 170372 204917 170373
rect 204851 170308 204852 170372
rect 204916 170308 204917 170372
rect 204851 170307 204917 170308
rect 204667 167652 204733 167653
rect 204667 167588 204668 167652
rect 204732 167588 204733 167652
rect 204667 167587 204733 167588
rect 204115 164932 204181 164933
rect 204115 164868 204116 164932
rect 204180 164868 204181 164932
rect 204115 164867 204181 164868
rect 203563 163572 203629 163573
rect 203563 163508 203564 163572
rect 203628 163508 203629 163572
rect 203563 163507 203629 163508
rect 203379 162348 203445 162349
rect 203379 162284 203380 162348
rect 203444 162284 203445 162348
rect 203379 162283 203445 162284
rect 203195 162212 203261 162213
rect 203195 162148 203196 162212
rect 203260 162148 203261 162212
rect 203195 162147 203261 162148
rect 202643 161940 202709 161941
rect 202643 161876 202644 161940
rect 202708 161876 202709 161940
rect 202643 161875 202709 161876
rect 199883 159900 199949 159901
rect 199883 159836 199884 159900
rect 199948 159836 199949 159900
rect 199883 159835 199949 159836
rect 200987 159900 201053 159901
rect 200987 159836 200988 159900
rect 201052 159836 201053 159900
rect 200987 159835 201053 159836
rect 201355 159900 201421 159901
rect 201355 159836 201356 159900
rect 201420 159836 201421 159900
rect 201355 159835 201421 159836
rect 198411 159764 198477 159765
rect 198411 159762 198412 159764
rect 198230 159702 198412 159762
rect 198043 159628 198109 159629
rect 198043 159564 198044 159628
rect 198108 159564 198109 159628
rect 198043 159563 198109 159564
rect 198043 152556 198109 152557
rect 198043 152492 198044 152556
rect 198108 152492 198109 152556
rect 198043 152491 198109 152492
rect 198046 115157 198106 152491
rect 198043 115156 198109 115157
rect 198043 115092 198044 115156
rect 198108 115092 198109 115156
rect 198043 115091 198109 115092
rect 198230 98701 198290 159702
rect 198411 159700 198412 159702
rect 198476 159700 198477 159764
rect 198411 159699 198477 159700
rect 199331 159764 199397 159765
rect 199331 159700 199332 159764
rect 199396 159700 199397 159764
rect 199331 159699 199397 159700
rect 199147 158948 199213 158949
rect 199147 158884 199148 158948
rect 199212 158884 199213 158948
rect 199147 158883 199213 158884
rect 198411 158676 198477 158677
rect 198411 158612 198412 158676
rect 198476 158612 198477 158676
rect 198411 158611 198477 158612
rect 198595 158676 198661 158677
rect 198595 158612 198596 158676
rect 198660 158612 198661 158676
rect 198595 158611 198661 158612
rect 198414 139773 198474 158611
rect 198598 152557 198658 158611
rect 199150 154590 199210 158883
rect 199334 158405 199394 159699
rect 199699 158676 199765 158677
rect 199699 158612 199700 158676
rect 199764 158612 199765 158676
rect 199699 158611 199765 158612
rect 199515 158540 199581 158541
rect 199515 158476 199516 158540
rect 199580 158476 199581 158540
rect 199515 158475 199581 158476
rect 199331 158404 199397 158405
rect 199331 158340 199332 158404
rect 199396 158340 199397 158404
rect 199331 158339 199397 158340
rect 199150 154530 199394 154590
rect 198595 152556 198661 152557
rect 198595 152492 198596 152556
rect 198660 152492 198661 152556
rect 198595 152491 198661 152492
rect 198411 139772 198477 139773
rect 198411 139708 198412 139772
rect 198476 139708 198477 139772
rect 198411 139707 198477 139708
rect 198227 98700 198293 98701
rect 198227 98636 198228 98700
rect 198292 98636 198293 98700
rect 198227 98635 198293 98636
rect 197859 46204 197925 46205
rect 197859 46140 197860 46204
rect 197924 46140 197925 46204
rect 197859 46139 197925 46140
rect 198414 44845 198474 139707
rect 199334 131749 199394 154530
rect 199331 131748 199397 131749
rect 199331 131684 199332 131748
rect 199396 131684 199397 131748
rect 199331 131683 199397 131684
rect 199518 125493 199578 158475
rect 199702 154053 199762 158611
rect 199699 154052 199765 154053
rect 199699 153988 199700 154052
rect 199764 153988 199765 154052
rect 199699 153987 199765 153988
rect 199515 125492 199581 125493
rect 199515 125428 199516 125492
rect 199580 125428 199581 125492
rect 199515 125427 199581 125428
rect 199702 113797 199762 153987
rect 199699 113796 199765 113797
rect 199699 113732 199700 113796
rect 199764 113732 199765 113796
rect 199699 113731 199765 113732
rect 198411 44844 198477 44845
rect 198411 44780 198412 44844
rect 198476 44780 198477 44844
rect 198411 44779 198477 44780
rect 199886 42125 199946 159835
rect 200803 158676 200869 158677
rect 200803 158612 200804 158676
rect 200868 158612 200869 158676
rect 200803 158611 200869 158612
rect 200806 143309 200866 158611
rect 200803 143308 200869 143309
rect 200803 143244 200804 143308
rect 200868 143244 200869 143308
rect 200803 143243 200869 143244
rect 200806 106861 200866 143243
rect 200990 109717 201050 159835
rect 202646 159765 202706 161875
rect 202459 159764 202525 159765
rect 202459 159700 202460 159764
rect 202524 159700 202525 159764
rect 202459 159699 202525 159700
rect 202643 159764 202709 159765
rect 202643 159700 202644 159764
rect 202708 159700 202709 159764
rect 202643 159699 202709 159700
rect 202091 158676 202157 158677
rect 202091 158612 202092 158676
rect 202156 158612 202157 158676
rect 202091 158611 202157 158612
rect 201171 158540 201237 158541
rect 201171 158476 201172 158540
rect 201236 158476 201237 158540
rect 201171 158475 201237 158476
rect 201174 146165 201234 158475
rect 201355 158404 201421 158405
rect 201355 158340 201356 158404
rect 201420 158340 201421 158404
rect 201355 158339 201421 158340
rect 201171 146164 201237 146165
rect 201171 146100 201172 146164
rect 201236 146100 201237 146164
rect 201171 146099 201237 146100
rect 200987 109716 201053 109717
rect 200987 109652 200988 109716
rect 201052 109652 201053 109716
rect 200987 109651 201053 109652
rect 200803 106860 200869 106861
rect 200803 106796 200804 106860
rect 200868 106796 200869 106860
rect 200803 106795 200869 106796
rect 199883 42124 199949 42125
rect 199883 42060 199884 42124
rect 199948 42060 199949 42124
rect 199883 42059 199949 42060
rect 201174 37909 201234 146099
rect 201358 142357 201418 158339
rect 202094 143445 202154 158611
rect 202275 158540 202341 158541
rect 202275 158476 202276 158540
rect 202340 158476 202341 158540
rect 202275 158475 202341 158476
rect 202091 143444 202157 143445
rect 202091 143380 202092 143444
rect 202156 143380 202157 143444
rect 202091 143379 202157 143380
rect 202278 142901 202338 158475
rect 202462 157589 202522 159699
rect 202459 157588 202525 157589
rect 202459 157524 202460 157588
rect 202524 157524 202525 157588
rect 202459 157523 202525 157524
rect 202275 142900 202341 142901
rect 202275 142836 202276 142900
rect 202340 142836 202341 142900
rect 202275 142835 202341 142836
rect 201355 142356 201421 142357
rect 201355 142292 201356 142356
rect 201420 142292 201421 142356
rect 201355 142291 201421 142292
rect 201171 37908 201237 37909
rect 201171 37844 201172 37908
rect 201236 37844 201237 37908
rect 201171 37843 201237 37844
rect 201358 18597 201418 142291
rect 202278 104141 202338 142835
rect 202275 104140 202341 104141
rect 202275 104076 202276 104140
rect 202340 104076 202341 104140
rect 202275 104075 202341 104076
rect 202462 101421 202522 157523
rect 202459 101420 202525 101421
rect 202459 101356 202460 101420
rect 202524 101356 202525 101420
rect 202459 101355 202525 101356
rect 202646 71093 202706 159699
rect 203198 157997 203258 162147
rect 203382 159221 203442 162283
rect 203566 161261 203626 163507
rect 203563 161260 203629 161261
rect 203563 161196 203564 161260
rect 203628 161196 203629 161260
rect 203563 161195 203629 161196
rect 203563 160308 203629 160309
rect 203563 160244 203564 160308
rect 203628 160244 203629 160308
rect 203563 160243 203629 160244
rect 203379 159220 203445 159221
rect 203379 159156 203380 159220
rect 203444 159156 203445 159220
rect 203379 159155 203445 159156
rect 203566 158133 203626 160243
rect 204118 159901 204178 164867
rect 204670 159901 204730 167587
rect 204115 159900 204181 159901
rect 204115 159836 204116 159900
rect 204180 159836 204181 159900
rect 204115 159835 204181 159836
rect 204667 159900 204733 159901
rect 204667 159836 204668 159900
rect 204732 159836 204733 159900
rect 204667 159835 204733 159836
rect 204118 158677 204178 159835
rect 204854 159765 204914 170307
rect 205403 165068 205469 165069
rect 205403 165004 205404 165068
rect 205468 165004 205469 165068
rect 205403 165003 205469 165004
rect 205219 163436 205285 163437
rect 205219 163372 205220 163436
rect 205284 163372 205285 163436
rect 205219 163371 205285 163372
rect 205222 159901 205282 163371
rect 205406 159901 205466 165003
rect 205774 159901 205834 179963
rect 205955 175948 206021 175949
rect 205955 175884 205956 175948
rect 206020 175884 206021 175948
rect 205955 175883 206021 175884
rect 205219 159900 205285 159901
rect 205219 159836 205220 159900
rect 205284 159836 205285 159900
rect 205219 159835 205285 159836
rect 205403 159900 205469 159901
rect 205403 159836 205404 159900
rect 205468 159836 205469 159900
rect 205403 159835 205469 159836
rect 205771 159900 205837 159901
rect 205771 159836 205772 159900
rect 205836 159836 205837 159900
rect 205771 159835 205837 159836
rect 204851 159764 204917 159765
rect 204851 159700 204852 159764
rect 204916 159700 204917 159764
rect 204851 159699 204917 159700
rect 203931 158676 203997 158677
rect 203931 158612 203932 158676
rect 203996 158612 203997 158676
rect 203931 158611 203997 158612
rect 204115 158676 204181 158677
rect 204115 158612 204116 158676
rect 204180 158612 204181 158676
rect 204115 158611 204181 158612
rect 203747 158540 203813 158541
rect 203747 158476 203748 158540
rect 203812 158476 203813 158540
rect 203747 158475 203813 158476
rect 203563 158132 203629 158133
rect 203563 158068 203564 158132
rect 203628 158068 203629 158132
rect 203563 158067 203629 158068
rect 203195 157996 203261 157997
rect 203195 157932 203196 157996
rect 203260 157932 203261 157996
rect 203195 157931 203261 157932
rect 203750 155821 203810 158475
rect 203747 155820 203813 155821
rect 203747 155756 203748 155820
rect 203812 155756 203813 155820
rect 203747 155755 203813 155756
rect 203750 119373 203810 155755
rect 203934 147389 203994 158611
rect 204115 158404 204181 158405
rect 204115 158340 204116 158404
rect 204180 158340 204181 158404
rect 204115 158339 204181 158340
rect 203931 147388 203997 147389
rect 203931 147324 203932 147388
rect 203996 147324 203997 147388
rect 203931 147323 203997 147324
rect 203747 119372 203813 119373
rect 203747 119308 203748 119372
rect 203812 119308 203813 119372
rect 203747 119307 203813 119308
rect 203934 95845 203994 147323
rect 204118 144805 204178 158339
rect 204115 144804 204181 144805
rect 204115 144740 204116 144804
rect 204180 144740 204181 144804
rect 204115 144739 204181 144740
rect 203931 95844 203997 95845
rect 203931 95780 203932 95844
rect 203996 95780 203997 95844
rect 203931 95779 203997 95780
rect 202643 71092 202709 71093
rect 202643 71028 202644 71092
rect 202708 71028 202709 71092
rect 202643 71027 202709 71028
rect 204118 69597 204178 144739
rect 205222 90405 205282 159835
rect 205403 158676 205469 158677
rect 205403 158612 205404 158676
rect 205468 158612 205469 158676
rect 205403 158611 205469 158612
rect 205406 145757 205466 158611
rect 205403 145756 205469 145757
rect 205403 145692 205404 145756
rect 205468 145692 205469 145756
rect 205403 145691 205469 145692
rect 205219 90404 205285 90405
rect 205219 90340 205220 90404
rect 205284 90340 205285 90404
rect 205219 90339 205285 90340
rect 204115 69596 204181 69597
rect 204115 69532 204116 69596
rect 204180 69532 204181 69596
rect 204115 69531 204181 69532
rect 205406 35189 205466 145691
rect 205774 84829 205834 159835
rect 205958 159765 206018 175883
rect 206139 166292 206205 166293
rect 206139 166228 206140 166292
rect 206204 166228 206205 166292
rect 206139 166227 206205 166228
rect 205955 159764 206021 159765
rect 205955 159700 205956 159764
rect 206020 159700 206021 159764
rect 205955 159699 206021 159700
rect 205771 84828 205837 84829
rect 205771 84764 205772 84828
rect 205836 84764 205837 84828
rect 205771 84763 205837 84764
rect 205403 35188 205469 35189
rect 205403 35124 205404 35188
rect 205468 35124 205469 35188
rect 205403 35123 205469 35124
rect 201355 18596 201421 18597
rect 201355 18532 201356 18596
rect 201420 18532 201421 18596
rect 201355 18531 201421 18532
rect 197123 11660 197189 11661
rect 197123 11596 197124 11660
rect 197188 11596 197189 11660
rect 197123 11595 197189 11596
rect 195651 9076 195717 9077
rect 195651 9012 195652 9076
rect 195716 9012 195717 9076
rect 195651 9011 195717 9012
rect 195099 8940 195165 8941
rect 195099 8876 195100 8940
rect 195164 8876 195165 8940
rect 195099 8875 195165 8876
rect 205958 7581 206018 159699
rect 206142 159221 206202 166227
rect 206875 162076 206941 162077
rect 206875 162012 206876 162076
rect 206940 162012 206941 162076
rect 206875 162011 206941 162012
rect 206139 159220 206205 159221
rect 206139 159156 206140 159220
rect 206204 159156 206205 159220
rect 206139 159155 206205 159156
rect 206878 158677 206938 162011
rect 207798 159765 207858 182819
rect 207979 171732 208045 171733
rect 207979 171668 207980 171732
rect 208044 171668 208045 171732
rect 207979 171667 208045 171668
rect 207982 159901 208042 171667
rect 207979 159900 208045 159901
rect 207979 159836 207980 159900
rect 208044 159836 208045 159900
rect 207979 159835 208045 159836
rect 207795 159764 207861 159765
rect 207795 159700 207796 159764
rect 207860 159700 207861 159764
rect 207795 159699 207861 159700
rect 206875 158676 206941 158677
rect 206875 158612 206876 158676
rect 206940 158612 206941 158676
rect 206875 158611 206941 158612
rect 206878 157589 206938 158611
rect 208902 158541 208962 204851
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 208899 158540 208965 158541
rect 208899 158476 208900 158540
rect 208964 158476 208965 158540
rect 208899 158475 208965 158476
rect 206875 157588 206941 157589
rect 206875 157524 206876 157588
rect 206940 157524 206941 157588
rect 206875 157523 206941 157524
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 205955 7580 206021 7581
rect 205955 7516 205956 7580
rect 206020 7516 206021 7580
rect 205955 7515 206021 7516
rect 193075 6220 193141 6221
rect 193075 6156 193076 6220
rect 193140 6156 193141 6220
rect 193075 6155 193141 6156
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -1894 186134 -1862
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 223174 222134 258618
rect 222702 247050 222762 315963
rect 223067 295084 223133 295085
rect 223067 295020 223068 295084
rect 223132 295020 223133 295084
rect 223067 295019 223133 295020
rect 222702 246990 222946 247050
rect 222886 241773 222946 246990
rect 222883 241772 222949 241773
rect 222883 241708 222884 241772
rect 222948 241708 222949 241772
rect 222883 241707 222949 241708
rect 222699 240412 222765 240413
rect 222699 240348 222700 240412
rect 222764 240348 222765 240412
rect 222699 240347 222765 240348
rect 222702 238781 222762 240347
rect 222886 239322 222946 241707
rect 223070 239461 223130 295019
rect 223254 239733 223314 317051
rect 223435 316980 223501 316981
rect 223435 316916 223436 316980
rect 223500 316916 223501 316980
rect 223435 316915 223501 316916
rect 223438 240413 223498 316915
rect 224723 315212 224789 315213
rect 224723 315148 224724 315212
rect 224788 315148 224789 315212
rect 224723 315147 224789 315148
rect 223987 305828 224053 305829
rect 223987 305764 223988 305828
rect 224052 305764 224053 305828
rect 223987 305763 224053 305764
rect 223803 298076 223869 298077
rect 223803 298012 223804 298076
rect 223868 298012 223869 298076
rect 223803 298011 223869 298012
rect 223619 294676 223685 294677
rect 223619 294612 223620 294676
rect 223684 294612 223685 294676
rect 223619 294611 223685 294612
rect 223435 240412 223501 240413
rect 223435 240348 223436 240412
rect 223500 240348 223501 240412
rect 223435 240347 223501 240348
rect 223251 239732 223317 239733
rect 223251 239668 223252 239732
rect 223316 239668 223317 239732
rect 223251 239667 223317 239668
rect 223435 239732 223501 239733
rect 223435 239668 223436 239732
rect 223500 239668 223501 239732
rect 223435 239667 223501 239668
rect 223067 239460 223133 239461
rect 223067 239396 223068 239460
rect 223132 239396 223133 239460
rect 223067 239395 223133 239396
rect 223438 239322 223498 239667
rect 223622 239461 223682 294611
rect 223806 239733 223866 298011
rect 223803 239732 223869 239733
rect 223803 239668 223804 239732
rect 223868 239668 223869 239732
rect 223803 239667 223869 239668
rect 223990 239730 224050 305763
rect 224726 239869 224786 315147
rect 232267 314532 232333 314533
rect 232267 314468 232268 314532
rect 232332 314468 232333 314532
rect 232267 314467 232333 314468
rect 231531 311404 231597 311405
rect 231531 311340 231532 311404
rect 231596 311340 231597 311404
rect 231531 311339 231597 311340
rect 231163 311132 231229 311133
rect 231163 311068 231164 311132
rect 231228 311068 231229 311132
rect 231163 311067 231229 311068
rect 227483 310452 227549 310453
rect 227483 310388 227484 310452
rect 227548 310388 227549 310452
rect 227483 310387 227549 310388
rect 226195 310180 226261 310181
rect 226195 310116 226196 310180
rect 226260 310116 226261 310180
rect 226195 310115 226261 310116
rect 225827 296444 225893 296445
rect 225827 296380 225828 296444
rect 225892 296380 225893 296444
rect 225827 296379 225893 296380
rect 225459 289644 225525 289645
rect 225459 289580 225460 289644
rect 225524 289580 225525 289644
rect 225459 289579 225525 289580
rect 225275 241092 225341 241093
rect 225275 241028 225276 241092
rect 225340 241028 225341 241092
rect 225275 241027 225341 241028
rect 225278 240277 225338 241027
rect 225275 240276 225341 240277
rect 225275 240212 225276 240276
rect 225340 240212 225341 240276
rect 225275 240211 225341 240212
rect 225278 239869 225338 240211
rect 225462 239869 225522 289579
rect 225830 240005 225890 296379
rect 226011 241772 226077 241773
rect 226011 241708 226012 241772
rect 226076 241708 226077 241772
rect 226011 241707 226077 241708
rect 225827 240004 225893 240005
rect 225827 239940 225828 240004
rect 225892 239940 225893 240004
rect 225827 239939 225893 239940
rect 224723 239868 224789 239869
rect 224723 239804 224724 239868
rect 224788 239804 224789 239868
rect 224723 239803 224789 239804
rect 225275 239868 225341 239869
rect 225275 239804 225276 239868
rect 225340 239804 225341 239868
rect 225275 239803 225341 239804
rect 225459 239868 225525 239869
rect 225459 239804 225460 239868
rect 225524 239804 225525 239868
rect 225459 239803 225525 239804
rect 224171 239732 224237 239733
rect 224171 239730 224172 239732
rect 223990 239670 224172 239730
rect 223619 239460 223685 239461
rect 223619 239396 223620 239460
rect 223684 239396 223685 239460
rect 223619 239395 223685 239396
rect 222886 239262 223498 239322
rect 222699 238780 222765 238781
rect 222699 238716 222700 238780
rect 222764 238716 222765 238780
rect 222699 238715 222765 238716
rect 223806 238509 223866 239667
rect 223990 238781 224050 239670
rect 224171 239668 224172 239670
rect 224236 239668 224237 239732
rect 224171 239667 224237 239668
rect 225459 239052 225525 239053
rect 225459 238988 225460 239052
rect 225524 238988 225525 239052
rect 225459 238987 225525 238988
rect 223987 238780 224053 238781
rect 223987 238716 223988 238780
rect 224052 238716 224053 238780
rect 223987 238715 224053 238716
rect 223803 238508 223869 238509
rect 223803 238444 223804 238508
rect 223868 238444 223869 238508
rect 223803 238443 223869 238444
rect 224355 236060 224421 236061
rect 224355 235996 224356 236060
rect 224420 235996 224421 236060
rect 224355 235995 224421 235996
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 224358 220693 224418 235995
rect 225462 228445 225522 238987
rect 226014 238509 226074 241707
rect 226198 239461 226258 310115
rect 227299 296580 227365 296581
rect 227299 296516 227300 296580
rect 227364 296516 227365 296580
rect 227299 296515 227365 296516
rect 227115 296308 227181 296309
rect 227115 296244 227116 296308
rect 227180 296244 227181 296308
rect 227115 296243 227181 296244
rect 226931 296036 226997 296037
rect 226931 295972 226932 296036
rect 226996 295972 226997 296036
rect 226931 295971 226997 295972
rect 226747 241228 226813 241229
rect 226747 241164 226748 241228
rect 226812 241164 226813 241228
rect 226747 241163 226813 241164
rect 226379 240140 226445 240141
rect 226379 240076 226380 240140
rect 226444 240076 226445 240140
rect 226379 240075 226445 240076
rect 226195 239460 226261 239461
rect 226195 239396 226196 239460
rect 226260 239396 226261 239460
rect 226195 239395 226261 239396
rect 226382 239053 226442 240075
rect 226563 239868 226629 239869
rect 226563 239804 226564 239868
rect 226628 239804 226629 239868
rect 226563 239803 226629 239804
rect 226566 239461 226626 239803
rect 226750 239461 226810 241163
rect 226563 239460 226629 239461
rect 226563 239396 226564 239460
rect 226628 239396 226629 239460
rect 226563 239395 226629 239396
rect 226747 239460 226813 239461
rect 226747 239396 226748 239460
rect 226812 239396 226813 239460
rect 226747 239395 226813 239396
rect 226379 239052 226445 239053
rect 226379 238988 226380 239052
rect 226444 238988 226445 239052
rect 226379 238987 226445 238988
rect 226934 238645 226994 295971
rect 227118 239869 227178 296243
rect 227115 239868 227181 239869
rect 227115 239804 227116 239868
rect 227180 239804 227181 239868
rect 227115 239803 227181 239804
rect 227118 239053 227178 239803
rect 227302 239325 227362 296515
rect 227486 239461 227546 310387
rect 230243 309772 230309 309773
rect 230243 309708 230244 309772
rect 230308 309708 230309 309772
rect 230243 309707 230309 309708
rect 228955 309636 229021 309637
rect 228955 309572 228956 309636
rect 229020 309572 229021 309636
rect 228955 309571 229021 309572
rect 228771 296172 228837 296173
rect 228771 296108 228772 296172
rect 228836 296108 228837 296172
rect 228771 296107 228837 296108
rect 227851 294948 227917 294949
rect 227851 294884 227852 294948
rect 227916 294884 227917 294948
rect 227851 294883 227917 294884
rect 227854 240005 227914 294883
rect 228219 294404 228285 294405
rect 228219 294340 228220 294404
rect 228284 294340 228285 294404
rect 228219 294339 228285 294340
rect 228222 241637 228282 294339
rect 228219 241636 228285 241637
rect 228219 241572 228220 241636
rect 228284 241572 228285 241636
rect 228219 241571 228285 241572
rect 228035 240276 228101 240277
rect 228035 240212 228036 240276
rect 228100 240212 228101 240276
rect 228035 240211 228101 240212
rect 227851 240004 227917 240005
rect 227851 239940 227852 240004
rect 227916 239940 227917 240004
rect 227851 239939 227917 239940
rect 228038 239869 228098 240211
rect 227851 239868 227917 239869
rect 227851 239804 227852 239868
rect 227916 239804 227917 239868
rect 227851 239803 227917 239804
rect 228035 239868 228101 239869
rect 228035 239804 228036 239868
rect 228100 239804 228101 239868
rect 228035 239803 228101 239804
rect 227483 239460 227549 239461
rect 227483 239396 227484 239460
rect 227548 239396 227549 239460
rect 227483 239395 227549 239396
rect 227299 239324 227365 239325
rect 227299 239260 227300 239324
rect 227364 239260 227365 239324
rect 227299 239259 227365 239260
rect 227115 239052 227181 239053
rect 227115 238988 227116 239052
rect 227180 238988 227181 239052
rect 227115 238987 227181 238988
rect 226931 238644 226997 238645
rect 226931 238580 226932 238644
rect 226996 238580 226997 238644
rect 226931 238579 226997 238580
rect 226011 238508 226077 238509
rect 226011 238444 226012 238508
rect 226076 238444 226077 238508
rect 226011 238443 226077 238444
rect 227854 237554 227914 239803
rect 228222 239461 228282 241571
rect 228774 239733 228834 296107
rect 228771 239732 228837 239733
rect 228771 239668 228772 239732
rect 228836 239668 228837 239732
rect 228771 239667 228837 239668
rect 228219 239460 228285 239461
rect 228219 239396 228220 239460
rect 228284 239396 228285 239460
rect 228219 239395 228285 239396
rect 228035 239052 228101 239053
rect 228035 238988 228036 239052
rect 228100 238988 228101 239052
rect 228035 238987 228101 238988
rect 227486 237494 227914 237554
rect 227486 236333 227546 237494
rect 228038 237390 228098 238987
rect 228958 238645 229018 309571
rect 229691 295220 229757 295221
rect 229691 295156 229692 295220
rect 229756 295156 229757 295220
rect 229691 295155 229757 295156
rect 229139 239868 229205 239869
rect 229139 239804 229140 239868
rect 229204 239804 229205 239868
rect 229139 239803 229205 239804
rect 228955 238644 229021 238645
rect 228955 238580 228956 238644
rect 229020 238580 229021 238644
rect 228955 238579 229021 238580
rect 227670 237330 228098 237390
rect 227483 236332 227549 236333
rect 227483 236268 227484 236332
rect 227548 236268 227549 236332
rect 227483 236267 227549 236268
rect 225459 228444 225525 228445
rect 225459 228380 225460 228444
rect 225524 228380 225525 228444
rect 225459 228379 225525 228380
rect 224355 220692 224421 220693
rect 224355 220628 224356 220692
rect 224420 220628 224421 220692
rect 224355 220627 224421 220628
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 227670 159493 227730 237330
rect 229142 233205 229202 239803
rect 229694 239461 229754 295155
rect 229875 294812 229941 294813
rect 229875 294748 229876 294812
rect 229940 294748 229941 294812
rect 229875 294747 229941 294748
rect 229878 239869 229938 294747
rect 230059 294540 230125 294541
rect 230059 294476 230060 294540
rect 230124 294476 230125 294540
rect 230059 294475 230125 294476
rect 229875 239868 229941 239869
rect 229875 239804 229876 239868
rect 229940 239804 229941 239868
rect 229875 239803 229941 239804
rect 229691 239460 229757 239461
rect 229691 239396 229692 239460
rect 229756 239396 229757 239460
rect 229691 239395 229757 239396
rect 229878 239189 229938 239803
rect 230062 239189 230122 294475
rect 229875 239188 229941 239189
rect 229875 239124 229876 239188
rect 229940 239124 229941 239188
rect 229875 239123 229941 239124
rect 230059 239188 230125 239189
rect 230059 239124 230060 239188
rect 230124 239124 230125 239188
rect 230059 239123 230125 239124
rect 230246 238645 230306 309707
rect 230427 240004 230493 240005
rect 230427 239940 230428 240004
rect 230492 239940 230493 240004
rect 230427 239939 230493 239940
rect 230243 238644 230309 238645
rect 230243 238580 230244 238644
rect 230308 238580 230309 238644
rect 230243 238579 230309 238580
rect 229139 233204 229205 233205
rect 229139 233140 229140 233204
rect 229204 233140 229205 233204
rect 229139 233139 229205 233140
rect 227667 159492 227733 159493
rect 227667 159428 227668 159492
rect 227732 159428 227733 159492
rect 227667 159427 227733 159428
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 230430 139093 230490 239939
rect 230611 239868 230677 239869
rect 230611 239804 230612 239868
rect 230676 239866 230677 239868
rect 230676 239806 230858 239866
rect 230676 239804 230677 239806
rect 230611 239803 230677 239804
rect 230611 239732 230677 239733
rect 230611 239668 230612 239732
rect 230676 239668 230677 239732
rect 230611 239667 230677 239668
rect 230614 238645 230674 239667
rect 230611 238644 230677 238645
rect 230611 238580 230612 238644
rect 230676 238580 230677 238644
rect 230611 238579 230677 238580
rect 230798 231845 230858 239806
rect 231166 239733 231226 311067
rect 231347 309908 231413 309909
rect 231347 309844 231348 309908
rect 231412 309844 231413 309908
rect 231347 309843 231413 309844
rect 231350 239733 231410 309843
rect 231163 239732 231229 239733
rect 231163 239668 231164 239732
rect 231228 239668 231229 239732
rect 231163 239667 231229 239668
rect 231347 239732 231413 239733
rect 231347 239668 231348 239732
rect 231412 239668 231413 239732
rect 231347 239667 231413 239668
rect 230979 238372 231045 238373
rect 230979 238308 230980 238372
rect 231044 238308 231045 238372
rect 230979 238307 231045 238308
rect 230795 231844 230861 231845
rect 230795 231780 230796 231844
rect 230860 231780 230861 231844
rect 230795 231779 230861 231780
rect 230982 216477 231042 238307
rect 231166 237829 231226 239667
rect 231163 237828 231229 237829
rect 231163 237764 231164 237828
rect 231228 237764 231229 237828
rect 231163 237763 231229 237764
rect 231350 237421 231410 239667
rect 231534 239461 231594 311339
rect 231715 311268 231781 311269
rect 231715 311204 231716 311268
rect 231780 311204 231781 311268
rect 231715 311203 231781 311204
rect 231718 239869 231778 311203
rect 231899 241636 231965 241637
rect 231899 241572 231900 241636
rect 231964 241572 231965 241636
rect 231899 241571 231965 241572
rect 231715 239868 231781 239869
rect 231715 239804 231716 239868
rect 231780 239804 231781 239868
rect 231715 239803 231781 239804
rect 231902 239461 231962 241571
rect 232083 241364 232149 241365
rect 232083 241300 232084 241364
rect 232148 241300 232149 241364
rect 232083 241299 232149 241300
rect 232086 239733 232146 241299
rect 232270 239733 232330 314467
rect 232819 314396 232885 314397
rect 232819 314332 232820 314396
rect 232884 314332 232885 314396
rect 232819 314331 232885 314332
rect 232635 311812 232701 311813
rect 232635 311748 232636 311812
rect 232700 311748 232701 311812
rect 232635 311747 232701 311748
rect 232451 294268 232517 294269
rect 232451 294204 232452 294268
rect 232516 294204 232517 294268
rect 232451 294203 232517 294204
rect 232454 239869 232514 294203
rect 232638 241365 232698 311747
rect 232635 241364 232701 241365
rect 232635 241300 232636 241364
rect 232700 241300 232701 241364
rect 232635 241299 232701 241300
rect 232635 240956 232701 240957
rect 232635 240892 232636 240956
rect 232700 240892 232701 240956
rect 232635 240891 232701 240892
rect 232638 240413 232698 240891
rect 232635 240412 232701 240413
rect 232635 240348 232636 240412
rect 232700 240348 232701 240412
rect 232635 240347 232701 240348
rect 232822 239869 232882 314331
rect 234107 313172 234173 313173
rect 234107 313108 234108 313172
rect 234172 313108 234173 313172
rect 234107 313107 234173 313108
rect 233555 312628 233621 312629
rect 233555 312564 233556 312628
rect 233620 312564 233621 312628
rect 233555 312563 233621 312564
rect 233003 241500 233069 241501
rect 233003 241436 233004 241500
rect 233068 241436 233069 241500
rect 233003 241435 233069 241436
rect 232451 239868 232517 239869
rect 232451 239804 232452 239868
rect 232516 239804 232517 239868
rect 232451 239803 232517 239804
rect 232819 239868 232885 239869
rect 232819 239804 232820 239868
rect 232884 239804 232885 239868
rect 232819 239803 232885 239804
rect 232083 239732 232149 239733
rect 232083 239668 232084 239732
rect 232148 239668 232149 239732
rect 232083 239667 232149 239668
rect 232267 239732 232333 239733
rect 232267 239668 232268 239732
rect 232332 239668 232333 239732
rect 232267 239667 232333 239668
rect 232086 239461 232146 239667
rect 231531 239460 231597 239461
rect 231531 239396 231532 239460
rect 231596 239396 231597 239460
rect 231531 239395 231597 239396
rect 231899 239460 231965 239461
rect 231899 239396 231900 239460
rect 231964 239396 231965 239460
rect 231899 239395 231965 239396
rect 232083 239460 232149 239461
rect 232083 239396 232084 239460
rect 232148 239396 232149 239460
rect 232083 239395 232149 239396
rect 231347 237420 231413 237421
rect 231347 237356 231348 237420
rect 231412 237356 231413 237420
rect 231347 237355 231413 237356
rect 231902 235109 231962 239395
rect 231899 235108 231965 235109
rect 231899 235044 231900 235108
rect 231964 235044 231965 235108
rect 231899 235043 231965 235044
rect 232270 233477 232330 239667
rect 232454 239189 232514 239803
rect 232635 239460 232701 239461
rect 232635 239396 232636 239460
rect 232700 239396 232701 239460
rect 232635 239395 232701 239396
rect 232451 239188 232517 239189
rect 232451 239124 232452 239188
rect 232516 239124 232517 239188
rect 232451 239123 232517 239124
rect 232267 233476 232333 233477
rect 232267 233412 232268 233476
rect 232332 233412 232333 233476
rect 232267 233411 232333 233412
rect 230979 216476 231045 216477
rect 230979 216412 230980 216476
rect 231044 216412 231045 216476
rect 230979 216411 231045 216412
rect 230982 148477 231042 216411
rect 230979 148476 231045 148477
rect 230979 148412 230980 148476
rect 231044 148412 231045 148476
rect 230979 148411 231045 148412
rect 232638 142085 232698 239395
rect 232822 233613 232882 239803
rect 233006 239461 233066 241435
rect 233371 240956 233437 240957
rect 233371 240892 233372 240956
rect 233436 240892 233437 240956
rect 233371 240891 233437 240892
rect 233374 239869 233434 240891
rect 233371 239868 233437 239869
rect 233371 239804 233372 239868
rect 233436 239804 233437 239868
rect 233371 239803 233437 239804
rect 233003 239460 233069 239461
rect 233003 239396 233004 239460
rect 233068 239396 233069 239460
rect 233003 239395 233069 239396
rect 233558 239325 233618 312563
rect 233739 312492 233805 312493
rect 233739 312428 233740 312492
rect 233804 312428 233805 312492
rect 233739 312427 233805 312428
rect 233742 240005 233802 312427
rect 233923 240684 233989 240685
rect 233923 240620 233924 240684
rect 233988 240620 233989 240684
rect 233923 240619 233989 240620
rect 233739 240004 233805 240005
rect 233739 239940 233740 240004
rect 233804 239940 233805 240004
rect 233739 239939 233805 239940
rect 233926 239461 233986 240619
rect 234110 239869 234170 313107
rect 234475 312764 234541 312765
rect 234475 312700 234476 312764
rect 234540 312700 234541 312764
rect 234475 312699 234541 312700
rect 234291 240684 234357 240685
rect 234291 240620 234292 240684
rect 234356 240620 234357 240684
rect 234291 240619 234357 240620
rect 234107 239868 234173 239869
rect 234107 239804 234108 239868
rect 234172 239804 234173 239868
rect 234107 239803 234173 239804
rect 234294 239733 234354 240619
rect 234478 239733 234538 312699
rect 235211 301612 235277 301613
rect 235211 301548 235212 301612
rect 235276 301548 235277 301612
rect 235211 301547 235277 301548
rect 234843 241636 234909 241637
rect 234843 241572 234844 241636
rect 234908 241572 234909 241636
rect 234843 241571 234909 241572
rect 234659 239868 234725 239869
rect 234659 239804 234660 239868
rect 234724 239804 234725 239868
rect 234659 239803 234725 239804
rect 234291 239732 234357 239733
rect 234291 239668 234292 239732
rect 234356 239668 234357 239732
rect 234291 239667 234357 239668
rect 234475 239732 234541 239733
rect 234475 239668 234476 239732
rect 234540 239668 234541 239732
rect 234475 239667 234541 239668
rect 233923 239460 233989 239461
rect 233923 239396 233924 239460
rect 233988 239396 233989 239460
rect 233923 239395 233989 239396
rect 233555 239324 233621 239325
rect 233555 239260 233556 239324
rect 233620 239260 233621 239324
rect 233555 239259 233621 239260
rect 233187 239188 233253 239189
rect 233187 239124 233188 239188
rect 233252 239124 233253 239188
rect 233187 239123 233253 239124
rect 232819 233612 232885 233613
rect 232819 233548 232820 233612
rect 232884 233548 232885 233612
rect 232819 233547 232885 233548
rect 233190 155413 233250 239123
rect 234478 237390 234538 239667
rect 234662 239325 234722 239803
rect 234659 239324 234725 239325
rect 234659 239260 234660 239324
rect 234724 239260 234725 239324
rect 234659 239259 234725 239260
rect 234846 239050 234906 241571
rect 235027 240548 235093 240549
rect 235027 240484 235028 240548
rect 235092 240484 235093 240548
rect 235027 240483 235093 240484
rect 235030 239733 235090 240483
rect 235214 240277 235274 301547
rect 235211 240276 235277 240277
rect 235211 240212 235212 240276
rect 235276 240212 235277 240276
rect 235211 240211 235277 240212
rect 236315 240276 236381 240277
rect 236315 240212 236316 240276
rect 236380 240212 236381 240276
rect 236315 240211 236381 240212
rect 236318 239869 236378 240211
rect 236315 239868 236381 239869
rect 236315 239804 236316 239868
rect 236380 239804 236381 239868
rect 236315 239803 236381 239804
rect 235027 239732 235093 239733
rect 235027 239668 235028 239732
rect 235092 239668 235093 239732
rect 235027 239667 235093 239668
rect 235395 239460 235461 239461
rect 235395 239396 235396 239460
rect 235460 239396 235461 239460
rect 235395 239395 235461 239396
rect 234662 238990 234906 239050
rect 234662 238645 234722 238990
rect 234659 238644 234725 238645
rect 234659 238580 234660 238644
rect 234724 238580 234725 238644
rect 234659 238579 234725 238580
rect 234294 237330 234538 237390
rect 234294 231709 234354 237330
rect 234475 234700 234541 234701
rect 234475 234636 234476 234700
rect 234540 234636 234541 234700
rect 234475 234635 234541 234636
rect 234291 231708 234357 231709
rect 234291 231644 234292 231708
rect 234356 231644 234357 231708
rect 234291 231643 234357 231644
rect 234478 224909 234538 234635
rect 234475 224908 234541 224909
rect 234475 224844 234476 224908
rect 234540 224844 234541 224908
rect 234475 224843 234541 224844
rect 233187 155412 233253 155413
rect 233187 155348 233188 155412
rect 233252 155348 233253 155412
rect 233187 155347 233253 155348
rect 232635 142084 232701 142085
rect 232635 142020 232636 142084
rect 232700 142020 232701 142084
rect 232635 142019 232701 142020
rect 234662 139365 234722 238579
rect 234843 236332 234909 236333
rect 234843 236268 234844 236332
rect 234908 236268 234909 236332
rect 234843 236267 234909 236268
rect 234846 222869 234906 236267
rect 235398 223005 235458 239395
rect 235579 236060 235645 236061
rect 235579 235996 235580 236060
rect 235644 235996 235645 236060
rect 235579 235995 235645 235996
rect 235582 228309 235642 235995
rect 236318 235653 236378 239803
rect 236502 238781 236562 318411
rect 237971 318340 238037 318341
rect 237971 318276 237972 318340
rect 238036 318276 238037 318340
rect 237971 318275 238037 318276
rect 236683 315620 236749 315621
rect 236683 315556 236684 315620
rect 236748 315556 236749 315620
rect 236683 315555 236749 315556
rect 236686 239733 236746 315555
rect 237051 315484 237117 315485
rect 237051 315420 237052 315484
rect 237116 315420 237117 315484
rect 237051 315419 237117 315420
rect 236867 293316 236933 293317
rect 236867 293252 236868 293316
rect 236932 293252 236933 293316
rect 236867 293251 236933 293252
rect 236870 240277 236930 293251
rect 236867 240276 236933 240277
rect 236867 240212 236868 240276
rect 236932 240212 236933 240276
rect 236867 240211 236933 240212
rect 236683 239732 236749 239733
rect 236683 239668 236684 239732
rect 236748 239668 236749 239732
rect 236683 239667 236749 239668
rect 237054 239461 237114 315419
rect 237787 299436 237853 299437
rect 237787 299372 237788 299436
rect 237852 299372 237853 299436
rect 237787 299371 237853 299372
rect 237790 239869 237850 299371
rect 237974 241773 238034 318275
rect 244779 314668 244845 314669
rect 244779 314604 244780 314668
rect 244844 314604 244845 314668
rect 244779 314603 244845 314604
rect 242571 314124 242637 314125
rect 242571 314060 242572 314124
rect 242636 314060 242637 314124
rect 242571 314059 242637 314060
rect 241283 313988 241349 313989
rect 241283 313924 241284 313988
rect 241348 313924 241349 313988
rect 241283 313923 241349 313924
rect 239995 310316 240061 310317
rect 239995 310252 239996 310316
rect 240060 310252 240061 310316
rect 239995 310251 240061 310252
rect 239443 302836 239509 302837
rect 239443 302772 239444 302836
rect 239508 302772 239509 302836
rect 239443 302771 239509 302772
rect 239259 297532 239325 297533
rect 239259 297468 239260 297532
rect 239324 297468 239325 297532
rect 239259 297467 239325 297468
rect 238339 297396 238405 297397
rect 238339 297332 238340 297396
rect 238404 297332 238405 297396
rect 238339 297331 238405 297332
rect 238155 293452 238221 293453
rect 238155 293388 238156 293452
rect 238220 293388 238221 293452
rect 238155 293387 238221 293388
rect 237971 241772 238037 241773
rect 237971 241708 237972 241772
rect 238036 241708 238037 241772
rect 237971 241707 238037 241708
rect 237603 239868 237669 239869
rect 237603 239804 237604 239868
rect 237668 239804 237669 239868
rect 237603 239803 237669 239804
rect 237787 239868 237853 239869
rect 237787 239804 237788 239868
rect 237852 239804 237853 239868
rect 237787 239803 237853 239804
rect 237051 239460 237117 239461
rect 237051 239396 237052 239460
rect 237116 239396 237117 239460
rect 237051 239395 237117 239396
rect 237235 239324 237301 239325
rect 237235 239260 237236 239324
rect 237300 239260 237301 239324
rect 237235 239259 237301 239260
rect 237238 239053 237298 239259
rect 237235 239052 237301 239053
rect 237235 238988 237236 239052
rect 237300 238988 237301 239052
rect 237235 238987 237301 238988
rect 236499 238780 236565 238781
rect 236499 238716 236500 238780
rect 236564 238716 236565 238780
rect 236499 238715 236565 238716
rect 237235 238780 237301 238781
rect 237235 238716 237236 238780
rect 237300 238716 237301 238780
rect 237235 238715 237301 238716
rect 236499 236604 236565 236605
rect 236499 236540 236500 236604
rect 236564 236540 236565 236604
rect 236499 236539 236565 236540
rect 236315 235652 236381 235653
rect 236315 235588 236316 235652
rect 236380 235588 236381 235652
rect 236315 235587 236381 235588
rect 235579 228308 235645 228309
rect 235579 228244 235580 228308
rect 235644 228244 235645 228308
rect 235579 228243 235645 228244
rect 235395 223004 235461 223005
rect 235395 222940 235396 223004
rect 235460 222940 235461 223004
rect 235395 222939 235461 222940
rect 234843 222868 234909 222869
rect 234843 222804 234844 222868
rect 234908 222804 234909 222868
rect 234843 222803 234909 222804
rect 234659 139364 234725 139365
rect 234659 139300 234660 139364
rect 234724 139300 234725 139364
rect 234659 139299 234725 139300
rect 230427 139092 230493 139093
rect 230427 139028 230428 139092
rect 230492 139028 230493 139092
rect 230427 139027 230493 139028
rect 236502 137189 236562 236539
rect 237238 232797 237298 238715
rect 237606 237829 237666 239803
rect 238158 239461 238218 293387
rect 238342 239733 238402 297331
rect 239075 293180 239141 293181
rect 239075 293116 239076 293180
rect 239140 293116 239141 293180
rect 239075 293115 239141 293116
rect 238891 240412 238957 240413
rect 238891 240348 238892 240412
rect 238956 240348 238957 240412
rect 238891 240347 238957 240348
rect 238894 239733 238954 240347
rect 238339 239732 238405 239733
rect 238339 239668 238340 239732
rect 238404 239668 238405 239732
rect 238339 239667 238405 239668
rect 238891 239732 238957 239733
rect 238891 239668 238892 239732
rect 238956 239668 238957 239732
rect 238891 239667 238957 239668
rect 239078 239461 239138 293115
rect 239262 239869 239322 297467
rect 239446 240138 239506 302771
rect 239446 240078 239874 240138
rect 239259 239868 239325 239869
rect 239259 239804 239260 239868
rect 239324 239804 239325 239868
rect 239259 239803 239325 239804
rect 239627 239868 239693 239869
rect 239627 239804 239628 239868
rect 239692 239804 239693 239868
rect 239627 239803 239693 239804
rect 238155 239460 238221 239461
rect 238155 239396 238156 239460
rect 238220 239396 238221 239460
rect 238155 239395 238221 239396
rect 239075 239460 239141 239461
rect 239075 239396 239076 239460
rect 239140 239396 239141 239460
rect 239075 239395 239141 239396
rect 239262 238781 239322 239803
rect 239259 238780 239325 238781
rect 239259 238716 239260 238780
rect 239324 238716 239325 238780
rect 239259 238715 239325 238716
rect 237603 237828 237669 237829
rect 237603 237764 237604 237828
rect 237668 237764 237669 237828
rect 237603 237763 237669 237764
rect 238155 236740 238221 236741
rect 238155 236676 238156 236740
rect 238220 236676 238221 236740
rect 238155 236675 238221 236676
rect 237235 232796 237301 232797
rect 237235 232732 237236 232796
rect 237300 232732 237301 232796
rect 237235 232731 237301 232732
rect 237971 231844 238037 231845
rect 237971 231780 237972 231844
rect 238036 231780 238037 231844
rect 237971 231779 238037 231780
rect 237974 218925 238034 231779
rect 237971 218924 238037 218925
rect 237971 218860 237972 218924
rect 238036 218860 238037 218924
rect 237971 218859 238037 218860
rect 237974 140589 238034 218859
rect 238158 157861 238218 236675
rect 239630 235109 239690 239803
rect 239814 239733 239874 240078
rect 239811 239732 239877 239733
rect 239811 239668 239812 239732
rect 239876 239668 239877 239732
rect 239811 239667 239877 239668
rect 239627 235108 239693 235109
rect 239627 235044 239628 235108
rect 239692 235044 239693 235108
rect 239627 235043 239693 235044
rect 239814 230490 239874 239667
rect 239998 239461 240058 310251
rect 241099 310044 241165 310045
rect 241099 309980 241100 310044
rect 241164 309980 241165 310044
rect 241099 309979 241165 309980
rect 240915 301476 240981 301477
rect 240915 301412 240916 301476
rect 240980 301412 240981 301476
rect 240915 301411 240981 301412
rect 240731 289372 240797 289373
rect 240731 289308 240732 289372
rect 240796 289308 240797 289372
rect 240731 289307 240797 289308
rect 240734 288557 240794 289307
rect 240731 288556 240797 288557
rect 240731 288492 240732 288556
rect 240796 288492 240797 288556
rect 240731 288491 240797 288492
rect 240547 239868 240613 239869
rect 240547 239866 240548 239868
rect 240366 239806 240548 239866
rect 239995 239460 240061 239461
rect 239995 239396 239996 239460
rect 240060 239396 240061 239460
rect 239995 239395 240061 239396
rect 239995 235380 240061 235381
rect 239995 235316 239996 235380
rect 240060 235316 240061 235380
rect 239995 235315 240061 235316
rect 239446 230430 239874 230490
rect 239446 213485 239506 230430
rect 239998 218653 240058 235315
rect 240366 233885 240426 239806
rect 240547 239804 240548 239806
rect 240612 239804 240613 239868
rect 240547 239803 240613 239804
rect 240918 239733 240978 301411
rect 241102 239869 241162 309979
rect 241099 239868 241165 239869
rect 241099 239804 241100 239868
rect 241164 239804 241165 239868
rect 241099 239803 241165 239804
rect 240547 239732 240613 239733
rect 240547 239668 240548 239732
rect 240612 239668 240613 239732
rect 240547 239667 240613 239668
rect 240915 239732 240981 239733
rect 240915 239668 240916 239732
rect 240980 239668 240981 239732
rect 240915 239667 240981 239668
rect 241099 239732 241165 239733
rect 241099 239668 241100 239732
rect 241164 239668 241165 239732
rect 241099 239667 241165 239668
rect 240363 233884 240429 233885
rect 240363 233820 240364 233884
rect 240428 233820 240429 233884
rect 240363 233819 240429 233820
rect 240550 228581 240610 239667
rect 240731 238780 240797 238781
rect 240731 238716 240732 238780
rect 240796 238716 240797 238780
rect 240731 238715 240797 238716
rect 240547 228580 240613 228581
rect 240547 228516 240548 228580
rect 240612 228516 240613 228580
rect 240547 228515 240613 228516
rect 239995 218652 240061 218653
rect 239995 218588 239996 218652
rect 240060 218588 240061 218652
rect 239995 218587 240061 218588
rect 239998 218109 240058 218587
rect 239995 218108 240061 218109
rect 239995 218044 239996 218108
rect 240060 218044 240061 218108
rect 239995 218043 240061 218044
rect 239443 213484 239509 213485
rect 239443 213420 239444 213484
rect 239508 213420 239509 213484
rect 239443 213419 239509 213420
rect 238155 157860 238221 157861
rect 238155 157796 238156 157860
rect 238220 157796 238221 157860
rect 238155 157795 238221 157796
rect 237971 140588 238037 140589
rect 237971 140524 237972 140588
rect 238036 140524 238037 140588
rect 237971 140523 238037 140524
rect 240734 140317 240794 238715
rect 240915 235380 240981 235381
rect 240915 235316 240916 235380
rect 240980 235316 240981 235380
rect 240915 235315 240981 235316
rect 240918 154053 240978 235315
rect 241102 234837 241162 239667
rect 241286 239461 241346 313923
rect 242019 240820 242085 240821
rect 242019 240756 242020 240820
rect 242084 240756 242085 240820
rect 242019 240755 242085 240756
rect 242022 239869 242082 240755
rect 242574 239869 242634 314059
rect 242755 313852 242821 313853
rect 242755 313788 242756 313852
rect 242820 313788 242821 313852
rect 242755 313787 242821 313788
rect 242019 239868 242085 239869
rect 242019 239804 242020 239868
rect 242084 239804 242085 239868
rect 242019 239803 242085 239804
rect 242571 239868 242637 239869
rect 242571 239804 242572 239868
rect 242636 239804 242637 239868
rect 242571 239803 242637 239804
rect 241651 239732 241717 239733
rect 241651 239668 241652 239732
rect 241716 239668 241717 239732
rect 241651 239667 241717 239668
rect 241283 239460 241349 239461
rect 241283 239396 241284 239460
rect 241348 239396 241349 239460
rect 241283 239395 241349 239396
rect 241654 237965 241714 239667
rect 241651 237964 241717 237965
rect 241651 237900 241652 237964
rect 241716 237900 241717 237964
rect 241651 237899 241717 237900
rect 242019 237828 242085 237829
rect 242019 237764 242020 237828
rect 242084 237764 242085 237828
rect 242019 237763 242085 237764
rect 241099 234836 241165 234837
rect 241099 234772 241100 234836
rect 241164 234772 241165 234836
rect 241099 234771 241165 234772
rect 240915 154052 240981 154053
rect 240915 153988 240916 154052
rect 240980 153988 240981 154052
rect 240915 153987 240981 153988
rect 240731 140316 240797 140317
rect 240731 140252 240732 140316
rect 240796 140252 240797 140316
rect 240731 140251 240797 140252
rect 242022 140181 242082 237763
rect 242574 235789 242634 239803
rect 242758 239461 242818 313787
rect 244043 289372 244109 289373
rect 244043 289308 244044 289372
rect 244108 289308 244109 289372
rect 244043 289307 244109 289308
rect 244046 239733 244106 289307
rect 243491 239732 243557 239733
rect 243491 239668 243492 239732
rect 243556 239668 243557 239732
rect 243491 239667 243557 239668
rect 244043 239732 244109 239733
rect 244043 239668 244044 239732
rect 244108 239668 244109 239732
rect 244043 239667 244109 239668
rect 242755 239460 242821 239461
rect 242755 239396 242756 239460
rect 242820 239396 242821 239460
rect 242755 239395 242821 239396
rect 242755 236060 242821 236061
rect 242755 235996 242756 236060
rect 242820 235996 242821 236060
rect 242755 235995 242821 235996
rect 242571 235788 242637 235789
rect 242571 235724 242572 235788
rect 242636 235724 242637 235788
rect 242571 235723 242637 235724
rect 242758 229110 242818 235995
rect 243494 235109 243554 239667
rect 244782 239461 244842 314603
rect 245515 314260 245581 314261
rect 245515 314196 245516 314260
rect 245580 314196 245581 314260
rect 245515 314195 245581 314196
rect 245147 293588 245213 293589
rect 245147 293524 245148 293588
rect 245212 293524 245213 293588
rect 245147 293523 245213 293524
rect 244963 289100 245029 289101
rect 244963 289036 244964 289100
rect 245028 289036 245029 289100
rect 244963 289035 245029 289036
rect 244779 239460 244845 239461
rect 244779 239396 244780 239460
rect 244844 239396 244845 239460
rect 244779 239395 244845 239396
rect 244966 239189 245026 289035
rect 244963 239188 245029 239189
rect 244963 239124 244964 239188
rect 245028 239124 245029 239188
rect 244963 239123 245029 239124
rect 245150 238645 245210 293523
rect 245518 239869 245578 314195
rect 249563 313036 249629 313037
rect 249563 312972 249564 313036
rect 249628 312972 249629 313036
rect 249563 312971 249629 312972
rect 246987 305012 247053 305013
rect 246987 304948 246988 305012
rect 247052 304948 247053 305012
rect 246987 304947 247053 304948
rect 246803 304196 246869 304197
rect 246803 304132 246804 304196
rect 246868 304132 246869 304196
rect 246803 304131 246869 304132
rect 246619 291820 246685 291821
rect 246619 291756 246620 291820
rect 246684 291756 246685 291820
rect 246619 291755 246685 291756
rect 245699 290324 245765 290325
rect 245699 290260 245700 290324
rect 245764 290260 245765 290324
rect 245699 290259 245765 290260
rect 245702 289917 245762 290259
rect 245699 289916 245765 289917
rect 245699 289852 245700 289916
rect 245764 289852 245765 289916
rect 245699 289851 245765 289852
rect 246435 289644 246501 289645
rect 246435 289580 246436 289644
rect 246500 289580 246501 289644
rect 246435 289579 246501 289580
rect 246251 289508 246317 289509
rect 246251 289444 246252 289508
rect 246316 289444 246317 289508
rect 246251 289443 246317 289444
rect 245515 239868 245581 239869
rect 245515 239804 245516 239868
rect 245580 239804 245581 239868
rect 245515 239803 245581 239804
rect 246067 239868 246133 239869
rect 246067 239804 246068 239868
rect 246132 239804 246133 239868
rect 246067 239803 246133 239804
rect 245518 238645 245578 239803
rect 245883 239732 245949 239733
rect 245883 239668 245884 239732
rect 245948 239668 245949 239732
rect 245883 239667 245949 239668
rect 245147 238644 245213 238645
rect 245147 238580 245148 238644
rect 245212 238580 245213 238644
rect 245147 238579 245213 238580
rect 245515 238644 245581 238645
rect 245515 238580 245516 238644
rect 245580 238580 245581 238644
rect 245515 238579 245581 238580
rect 244411 237012 244477 237013
rect 244411 236948 244412 237012
rect 244476 236948 244477 237012
rect 244411 236947 244477 236948
rect 243859 235652 243925 235653
rect 243859 235588 243860 235652
rect 243924 235588 243925 235652
rect 243859 235587 243925 235588
rect 243491 235108 243557 235109
rect 243491 235044 243492 235108
rect 243556 235044 243557 235108
rect 243491 235043 243557 235044
rect 242206 229050 242818 229110
rect 242206 219333 242266 229050
rect 242203 219332 242269 219333
rect 242203 219268 242204 219332
rect 242268 219268 242269 219332
rect 242203 219267 242269 219268
rect 242206 140725 242266 219267
rect 243862 219197 243922 235587
rect 244043 235516 244109 235517
rect 244043 235452 244044 235516
rect 244108 235452 244109 235516
rect 244043 235451 244109 235452
rect 243859 219196 243925 219197
rect 243859 219132 243860 219196
rect 243924 219132 243925 219196
rect 243859 219131 243925 219132
rect 243862 218109 243922 219131
rect 244046 219061 244106 235451
rect 244043 219060 244109 219061
rect 244043 218996 244044 219060
rect 244108 218996 244109 219060
rect 244043 218995 244109 218996
rect 244046 218245 244106 218995
rect 244043 218244 244109 218245
rect 244043 218180 244044 218244
rect 244108 218180 244109 218244
rect 244043 218179 244109 218180
rect 243859 218108 243925 218109
rect 243859 218044 243860 218108
rect 243924 218044 243925 218108
rect 243859 218043 243925 218044
rect 244414 213621 244474 236947
rect 244411 213620 244477 213621
rect 244411 213556 244412 213620
rect 244476 213556 244477 213620
rect 244411 213555 244477 213556
rect 245886 157997 245946 239667
rect 246070 239189 246130 239803
rect 246254 239597 246314 289443
rect 246438 288693 246498 289579
rect 246435 288692 246501 288693
rect 246435 288628 246436 288692
rect 246500 288628 246501 288692
rect 246435 288627 246501 288628
rect 246622 248430 246682 291755
rect 246438 248370 246682 248430
rect 246438 239869 246498 248370
rect 246435 239868 246501 239869
rect 246435 239804 246436 239868
rect 246500 239804 246501 239868
rect 246435 239803 246501 239804
rect 246251 239596 246317 239597
rect 246251 239532 246252 239596
rect 246316 239532 246317 239596
rect 246251 239531 246317 239532
rect 246067 239188 246133 239189
rect 246067 239124 246068 239188
rect 246132 239124 246133 239188
rect 246067 239123 246133 239124
rect 246254 237829 246314 239531
rect 246251 237828 246317 237829
rect 246251 237764 246252 237828
rect 246316 237764 246317 237828
rect 246251 237763 246317 237764
rect 245883 157996 245949 157997
rect 245883 157932 245884 157996
rect 245948 157932 245949 157996
rect 245883 157931 245949 157932
rect 242203 140724 242269 140725
rect 242203 140660 242204 140724
rect 242268 140660 242269 140724
rect 242203 140659 242269 140660
rect 246438 140453 246498 239803
rect 246806 239733 246866 304131
rect 246803 239732 246869 239733
rect 246803 239668 246804 239732
rect 246868 239668 246869 239732
rect 246803 239667 246869 239668
rect 246990 239594 247050 304947
rect 247171 289644 247237 289645
rect 247171 289580 247172 289644
rect 247236 289580 247237 289644
rect 247171 289579 247237 289580
rect 247174 247050 247234 289579
rect 247539 289508 247605 289509
rect 247539 289444 247540 289508
rect 247604 289444 247605 289508
rect 247539 289443 247605 289444
rect 247542 248430 247602 289443
rect 247542 248370 247970 248430
rect 247174 246990 247602 247050
rect 247542 239869 247602 246990
rect 247355 239868 247421 239869
rect 247355 239804 247356 239868
rect 247420 239804 247421 239868
rect 247355 239803 247421 239804
rect 247539 239868 247605 239869
rect 247539 239804 247540 239868
rect 247604 239804 247605 239868
rect 247539 239803 247605 239804
rect 247171 239596 247237 239597
rect 247171 239594 247172 239596
rect 246990 239534 247172 239594
rect 247171 239532 247172 239534
rect 247236 239532 247237 239596
rect 247171 239531 247237 239532
rect 247174 239325 247234 239531
rect 247171 239324 247237 239325
rect 247171 239260 247172 239324
rect 247236 239260 247237 239324
rect 247171 239259 247237 239260
rect 247171 238644 247237 238645
rect 247171 238580 247172 238644
rect 247236 238580 247237 238644
rect 247171 238579 247237 238580
rect 247174 236061 247234 238579
rect 247358 236877 247418 239803
rect 247542 238917 247602 239803
rect 247910 239597 247970 248370
rect 248827 239868 248893 239869
rect 248827 239804 248828 239868
rect 248892 239804 248893 239868
rect 248827 239803 248893 239804
rect 248830 239597 248890 239803
rect 249566 239597 249626 312971
rect 251035 312900 251101 312901
rect 251035 312836 251036 312900
rect 251100 312836 251101 312900
rect 251035 312835 251101 312836
rect 250851 312356 250917 312357
rect 250851 312292 250852 312356
rect 250916 312292 250917 312356
rect 250851 312291 250917 312292
rect 250667 287740 250733 287741
rect 250667 287676 250668 287740
rect 250732 287676 250733 287740
rect 250667 287675 250733 287676
rect 249931 239868 249997 239869
rect 249931 239804 249932 239868
rect 249996 239804 249997 239868
rect 249931 239803 249997 239804
rect 250115 239868 250181 239869
rect 250115 239804 250116 239868
rect 250180 239804 250181 239868
rect 250115 239803 250181 239804
rect 247907 239596 247973 239597
rect 247907 239532 247908 239596
rect 247972 239532 247973 239596
rect 247907 239531 247973 239532
rect 248827 239596 248893 239597
rect 248827 239532 248828 239596
rect 248892 239532 248893 239596
rect 248827 239531 248893 239532
rect 249563 239596 249629 239597
rect 249563 239532 249564 239596
rect 249628 239532 249629 239596
rect 249563 239531 249629 239532
rect 247539 238916 247605 238917
rect 247539 238852 247540 238916
rect 247604 238852 247605 238916
rect 247539 238851 247605 238852
rect 247910 237693 247970 239531
rect 249379 239460 249445 239461
rect 249379 239396 249380 239460
rect 249444 239396 249445 239460
rect 249379 239395 249445 239396
rect 249195 239188 249261 239189
rect 249195 239124 249196 239188
rect 249260 239124 249261 239188
rect 249195 239123 249261 239124
rect 248275 238644 248341 238645
rect 248275 238580 248276 238644
rect 248340 238580 248341 238644
rect 248275 238579 248341 238580
rect 247907 237692 247973 237693
rect 247907 237628 247908 237692
rect 247972 237628 247973 237692
rect 247907 237627 247973 237628
rect 247355 236876 247421 236877
rect 247355 236812 247356 236876
rect 247420 236812 247421 236876
rect 247355 236811 247421 236812
rect 247171 236060 247237 236061
rect 247171 235996 247172 236060
rect 247236 235996 247237 236060
rect 247171 235995 247237 235996
rect 247723 236060 247789 236061
rect 247723 235996 247724 236060
rect 247788 235996 247789 236060
rect 247723 235995 247789 235996
rect 247726 220557 247786 235995
rect 248278 227357 248338 238579
rect 249011 230076 249077 230077
rect 249011 230012 249012 230076
rect 249076 230012 249077 230076
rect 249011 230011 249077 230012
rect 248275 227356 248341 227357
rect 248275 227292 248276 227356
rect 248340 227292 248341 227356
rect 248275 227291 248341 227292
rect 249014 222597 249074 230011
rect 249011 222596 249077 222597
rect 249011 222532 249012 222596
rect 249076 222532 249077 222596
rect 249011 222531 249077 222532
rect 249198 220965 249258 239123
rect 249382 221917 249442 239395
rect 249566 237965 249626 239531
rect 249563 237964 249629 237965
rect 249563 237900 249564 237964
rect 249628 237900 249629 237964
rect 249563 237899 249629 237900
rect 249934 237390 249994 239803
rect 250118 239461 250178 239803
rect 250670 239597 250730 287675
rect 250667 239596 250733 239597
rect 250667 239532 250668 239596
rect 250732 239532 250733 239596
rect 250667 239531 250733 239532
rect 250854 239461 250914 312291
rect 251038 239597 251098 312835
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 251771 289508 251837 289509
rect 251771 289444 251772 289508
rect 251836 289444 251837 289508
rect 251771 289443 251837 289444
rect 252691 289508 252757 289509
rect 252691 289444 252692 289508
rect 252756 289444 252757 289508
rect 252691 289443 252757 289444
rect 251774 239597 251834 289443
rect 252694 239869 252754 289443
rect 253794 255454 254414 290898
rect 257514 705798 258134 705830
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 278635 451892 278701 451893
rect 278635 451828 278636 451892
rect 278700 451828 278701 451892
rect 278635 451827 278701 451828
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 277899 372196 277965 372197
rect 277899 372132 277900 372196
rect 277964 372132 277965 372196
rect 277899 372131 277965 372132
rect 276611 372060 276677 372061
rect 276611 371996 276612 372060
rect 276676 371996 276677 372060
rect 276611 371995 276677 371996
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 276614 330445 276674 371995
rect 276611 330444 276677 330445
rect 276611 330380 276612 330444
rect 276676 330380 276677 330444
rect 276611 330379 276677 330380
rect 277902 323645 277962 372131
rect 278638 369341 278698 451827
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289123 398988 289189 398989
rect 289123 398924 289124 398988
rect 289188 398924 289189 398988
rect 289123 398923 289189 398924
rect 283419 397220 283485 397221
rect 283419 397156 283420 397220
rect 283484 397156 283485 397220
rect 283419 397155 283485 397156
rect 282867 392052 282933 392053
rect 282867 391988 282868 392052
rect 282932 391988 282933 392052
rect 282867 391987 282933 391988
rect 281395 387156 281461 387157
rect 281395 387092 281396 387156
rect 281460 387092 281461 387156
rect 281395 387091 281461 387092
rect 279371 375460 279437 375461
rect 279371 375396 279372 375460
rect 279436 375396 279437 375460
rect 279371 375395 279437 375396
rect 278635 369340 278701 369341
rect 278635 369276 278636 369340
rect 278700 369276 278701 369340
rect 278635 369275 278701 369276
rect 278638 368661 278698 369275
rect 278635 368660 278701 368661
rect 278635 368596 278636 368660
rect 278700 368596 278701 368660
rect 278635 368595 278701 368596
rect 277899 323644 277965 323645
rect 277899 323580 277900 323644
rect 277964 323580 277965 323644
rect 277899 323579 277965 323580
rect 259315 311540 259381 311541
rect 259315 311476 259316 311540
rect 259380 311476 259381 311540
rect 259315 311475 259381 311476
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257107 286380 257173 286381
rect 257107 286316 257108 286380
rect 257172 286316 257173 286380
rect 257107 286315 257173 286316
rect 256923 267204 256989 267205
rect 256923 267140 256924 267204
rect 256988 267140 256989 267204
rect 256923 267139 256989 267140
rect 255819 267068 255885 267069
rect 255819 267004 255820 267068
rect 255884 267004 255885 267068
rect 255819 267003 255885 267004
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 251955 239868 252021 239869
rect 251955 239804 251956 239868
rect 252020 239804 252021 239868
rect 251955 239803 252021 239804
rect 252691 239868 252757 239869
rect 252691 239804 252692 239868
rect 252756 239804 252757 239868
rect 252691 239803 252757 239804
rect 253427 239868 253493 239869
rect 253427 239804 253428 239868
rect 253492 239804 253493 239868
rect 253427 239803 253493 239804
rect 251035 239596 251101 239597
rect 251035 239532 251036 239596
rect 251100 239532 251101 239596
rect 251035 239531 251101 239532
rect 251771 239596 251837 239597
rect 251771 239532 251772 239596
rect 251836 239532 251837 239596
rect 251771 239531 251837 239532
rect 250115 239460 250181 239461
rect 250115 239396 250116 239460
rect 250180 239396 250181 239460
rect 250115 239395 250181 239396
rect 250851 239460 250917 239461
rect 250851 239396 250852 239460
rect 250916 239396 250917 239460
rect 250851 239395 250917 239396
rect 250299 238644 250365 238645
rect 250299 238580 250300 238644
rect 250364 238580 250365 238644
rect 250299 238579 250365 238580
rect 249566 237330 249994 237390
rect 249379 221916 249445 221917
rect 249379 221852 249380 221916
rect 249444 221852 249445 221916
rect 249379 221851 249445 221852
rect 249195 220964 249261 220965
rect 249195 220900 249196 220964
rect 249260 220900 249261 220964
rect 249195 220899 249261 220900
rect 246987 220556 247053 220557
rect 246987 220492 246988 220556
rect 247052 220492 247053 220556
rect 246987 220491 247053 220492
rect 247723 220556 247789 220557
rect 247723 220492 247724 220556
rect 247788 220492 247789 220556
rect 247723 220491 247789 220492
rect 246990 220285 247050 220491
rect 246987 220284 247053 220285
rect 246987 220220 246988 220284
rect 247052 220220 247053 220284
rect 246987 220219 247053 220220
rect 249382 141949 249442 221851
rect 249566 220829 249626 237330
rect 249747 228580 249813 228581
rect 249747 228516 249748 228580
rect 249812 228516 249813 228580
rect 249747 228515 249813 228516
rect 249750 227085 249810 228515
rect 249747 227084 249813 227085
rect 249747 227020 249748 227084
rect 249812 227020 249813 227084
rect 249747 227019 249813 227020
rect 249747 222596 249813 222597
rect 249747 222532 249748 222596
rect 249812 222532 249813 222596
rect 249747 222531 249813 222532
rect 249750 221645 249810 222531
rect 249747 221644 249813 221645
rect 249747 221580 249748 221644
rect 249812 221580 249813 221644
rect 249747 221579 249813 221580
rect 249563 220828 249629 220829
rect 249563 220764 249564 220828
rect 249628 220764 249629 220828
rect 249563 220763 249629 220764
rect 249379 141948 249445 141949
rect 249379 141884 249380 141948
rect 249444 141884 249445 141948
rect 249379 141883 249445 141884
rect 246435 140452 246501 140453
rect 246435 140388 246436 140452
rect 246500 140388 246501 140452
rect 246435 140387 246501 140388
rect 242019 140180 242085 140181
rect 242019 140116 242020 140180
rect 242084 140116 242085 140180
rect 242019 140115 242085 140116
rect 250302 137461 250362 238579
rect 251035 237420 251101 237421
rect 251035 237356 251036 237420
rect 251100 237356 251101 237420
rect 251035 237355 251101 237356
rect 250667 236060 250733 236061
rect 250667 235996 250668 236060
rect 250732 235996 250733 236060
rect 250667 235995 250733 235996
rect 250670 231165 250730 235995
rect 250667 231164 250733 231165
rect 250667 231100 250668 231164
rect 250732 231100 250733 231164
rect 250667 231099 250733 231100
rect 251038 228581 251098 237355
rect 251774 236605 251834 239531
rect 251771 236604 251837 236605
rect 251771 236540 251772 236604
rect 251836 236540 251837 236604
rect 251771 236539 251837 236540
rect 251958 232661 252018 239803
rect 252694 238645 252754 239803
rect 252691 238644 252757 238645
rect 252691 238580 252692 238644
rect 252756 238580 252757 238644
rect 252691 238579 252757 238580
rect 252323 237692 252389 237693
rect 252323 237628 252324 237692
rect 252388 237628 252389 237692
rect 252323 237627 252389 237628
rect 252139 237012 252205 237013
rect 252139 236948 252140 237012
rect 252204 236948 252205 237012
rect 252139 236947 252205 236948
rect 251955 232660 252021 232661
rect 251955 232596 251956 232660
rect 252020 232596 252021 232660
rect 251955 232595 252021 232596
rect 251035 228580 251101 228581
rect 251035 228516 251036 228580
rect 251100 228516 251101 228580
rect 251035 228515 251101 228516
rect 251958 219450 252018 232595
rect 252142 223413 252202 236947
rect 252139 223412 252205 223413
rect 252139 223348 252140 223412
rect 252204 223348 252205 223412
rect 252139 223347 252205 223348
rect 252326 222730 252386 237627
rect 252691 237420 252757 237421
rect 252691 237356 252692 237420
rect 252756 237356 252757 237420
rect 252691 237355 252757 237356
rect 252694 233069 252754 237355
rect 252691 233068 252757 233069
rect 252691 233004 252692 233068
rect 252756 233004 252757 233068
rect 252691 233003 252757 233004
rect 252507 223412 252573 223413
rect 252507 223348 252508 223412
rect 252572 223348 252573 223412
rect 252507 223347 252573 223348
rect 252510 222869 252570 223347
rect 252507 222868 252573 222869
rect 252507 222804 252508 222868
rect 252572 222804 252573 222868
rect 252507 222803 252573 222804
rect 252507 222732 252573 222733
rect 252507 222730 252508 222732
rect 252326 222670 252508 222730
rect 252507 222668 252508 222670
rect 252572 222668 252573 222732
rect 252507 222667 252573 222668
rect 252510 221781 252570 222667
rect 253430 222189 253490 239803
rect 253427 222188 253493 222189
rect 253427 222124 253428 222188
rect 253492 222124 253493 222188
rect 253427 222123 253493 222124
rect 252507 221780 252573 221781
rect 252507 221716 252508 221780
rect 252572 221716 252573 221780
rect 252507 221715 252573 221716
rect 251774 219390 252018 219450
rect 253794 219454 254414 254898
rect 254715 239868 254781 239869
rect 254715 239804 254716 239868
rect 254780 239866 254781 239868
rect 254780 239806 254962 239866
rect 254780 239804 254781 239806
rect 254715 239803 254781 239804
rect 254902 225997 254962 239806
rect 255822 239733 255882 267003
rect 256371 265572 256437 265573
rect 256371 265508 256372 265572
rect 256436 265508 256437 265572
rect 256371 265507 256437 265508
rect 256187 257412 256253 257413
rect 256187 257348 256188 257412
rect 256252 257348 256253 257412
rect 256187 257347 256253 257348
rect 256003 239868 256069 239869
rect 256003 239804 256004 239868
rect 256068 239804 256069 239868
rect 256003 239803 256069 239804
rect 255819 239732 255885 239733
rect 255819 239668 255820 239732
rect 255884 239668 255885 239732
rect 255819 239667 255885 239668
rect 255635 238644 255701 238645
rect 255635 238580 255636 238644
rect 255700 238580 255701 238644
rect 255635 238579 255701 238580
rect 255451 237692 255517 237693
rect 255451 237628 255452 237692
rect 255516 237628 255517 237692
rect 255451 237627 255517 237628
rect 255267 236604 255333 236605
rect 255267 236540 255268 236604
rect 255332 236540 255333 236604
rect 255267 236539 255333 236540
rect 255270 230349 255330 236539
rect 255267 230348 255333 230349
rect 255267 230284 255268 230348
rect 255332 230284 255333 230348
rect 255267 230283 255333 230284
rect 254899 225996 254965 225997
rect 254899 225932 254900 225996
rect 254964 225932 254965 225996
rect 254899 225931 254965 225932
rect 255454 220149 255514 237627
rect 255638 225725 255698 238579
rect 255635 225724 255701 225725
rect 255635 225660 255636 225724
rect 255700 225660 255701 225724
rect 255635 225659 255701 225660
rect 255451 220148 255517 220149
rect 255451 220084 255452 220148
rect 255516 220084 255517 220148
rect 255451 220083 255517 220084
rect 251774 137597 251834 219390
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 255822 214981 255882 239667
rect 256006 236333 256066 239803
rect 256190 239461 256250 257347
rect 256187 239460 256253 239461
rect 256187 239396 256188 239460
rect 256252 239396 256253 239460
rect 256187 239395 256253 239396
rect 256374 239053 256434 265507
rect 256555 241636 256621 241637
rect 256555 241572 256556 241636
rect 256620 241572 256621 241636
rect 256555 241571 256621 241572
rect 256558 239733 256618 241571
rect 256926 239733 256986 267139
rect 257110 240005 257170 286315
rect 257514 259174 258134 294618
rect 259131 260132 259197 260133
rect 259131 260068 259132 260132
rect 259196 260068 259197 260132
rect 259131 260067 259197 260068
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257291 242316 257357 242317
rect 257291 242252 257292 242316
rect 257356 242252 257357 242316
rect 257291 242251 257357 242252
rect 257107 240004 257173 240005
rect 257107 239940 257108 240004
rect 257172 239940 257173 240004
rect 257107 239939 257173 239940
rect 256555 239732 256621 239733
rect 256555 239668 256556 239732
rect 256620 239668 256621 239732
rect 256555 239667 256621 239668
rect 256923 239732 256989 239733
rect 256923 239668 256924 239732
rect 256988 239668 256989 239732
rect 256923 239667 256989 239668
rect 257294 239461 257354 242251
rect 257291 239460 257357 239461
rect 257291 239396 257292 239460
rect 257356 239396 257357 239460
rect 257291 239395 257357 239396
rect 256371 239052 256437 239053
rect 256371 238988 256372 239052
rect 256436 238988 256437 239052
rect 256371 238987 256437 238988
rect 256003 236332 256069 236333
rect 256003 236268 256004 236332
rect 256068 236268 256069 236332
rect 256003 236267 256069 236268
rect 257107 233476 257173 233477
rect 257107 233412 257108 233476
rect 257172 233412 257173 233476
rect 257107 233411 257173 233412
rect 257110 221781 257170 233411
rect 257514 223174 258134 258618
rect 258395 240004 258461 240005
rect 258395 239940 258396 240004
rect 258460 240002 258461 240004
rect 258460 239942 258642 240002
rect 258460 239940 258461 239942
rect 258395 239939 258461 239940
rect 258395 236876 258461 236877
rect 258395 236812 258396 236876
rect 258460 236812 258461 236876
rect 258395 236811 258461 236812
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257107 221780 257173 221781
rect 257107 221716 257108 221780
rect 257172 221716 257173 221780
rect 257107 221715 257173 221716
rect 255819 214980 255885 214981
rect 255819 214916 255820 214980
rect 255884 214916 255885 214980
rect 255819 214915 255885 214916
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 251771 137596 251837 137597
rect 251771 137532 251772 137596
rect 251836 137532 251837 137596
rect 251771 137531 251837 137532
rect 250299 137460 250365 137461
rect 250299 137396 250300 137460
rect 250364 137396 250365 137460
rect 250299 137395 250365 137396
rect 236499 137188 236565 137189
rect 236499 137124 236500 137188
rect 236564 137124 236565 137188
rect 236499 137123 236565 137124
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -1894 222134 -1862
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 187174 258134 222618
rect 258398 222053 258458 236811
rect 258582 233613 258642 239942
rect 259134 239869 259194 260067
rect 259318 240005 259378 311475
rect 270355 308548 270421 308549
rect 270355 308484 270356 308548
rect 270420 308484 270421 308548
rect 270355 308483 270421 308484
rect 269619 300116 269685 300117
rect 269619 300052 269620 300116
rect 269684 300052 269685 300116
rect 269619 300051 269685 300052
rect 265019 271148 265085 271149
rect 265019 271084 265020 271148
rect 265084 271084 265085 271148
rect 265019 271083 265085 271084
rect 260603 264348 260669 264349
rect 260603 264284 260604 264348
rect 260668 264284 260669 264348
rect 260603 264283 260669 264284
rect 259867 242452 259933 242453
rect 259867 242388 259868 242452
rect 259932 242388 259933 242452
rect 259867 242387 259933 242388
rect 259315 240004 259381 240005
rect 259315 239940 259316 240004
rect 259380 239940 259381 240004
rect 259315 239939 259381 239940
rect 258763 239868 258829 239869
rect 258763 239804 258764 239868
rect 258828 239804 258829 239868
rect 258763 239803 258829 239804
rect 259131 239868 259197 239869
rect 259131 239804 259132 239868
rect 259196 239804 259197 239868
rect 259131 239803 259197 239804
rect 259683 239868 259749 239869
rect 259683 239804 259684 239868
rect 259748 239804 259749 239868
rect 259683 239803 259749 239804
rect 258766 237421 258826 239803
rect 259499 239732 259565 239733
rect 259499 239668 259500 239732
rect 259564 239668 259565 239732
rect 259499 239667 259565 239668
rect 259131 238236 259197 238237
rect 259131 238172 259132 238236
rect 259196 238172 259197 238236
rect 259131 238171 259197 238172
rect 258763 237420 258829 237421
rect 258763 237356 258764 237420
rect 258828 237356 258829 237420
rect 258763 237355 258829 237356
rect 258579 233612 258645 233613
rect 258579 233548 258580 233612
rect 258644 233548 258645 233612
rect 258579 233547 258645 233548
rect 259134 227629 259194 238171
rect 259502 229110 259562 239667
rect 259686 237829 259746 239803
rect 259870 239733 259930 242387
rect 260235 242180 260301 242181
rect 260235 242116 260236 242180
rect 260300 242116 260301 242180
rect 260235 242115 260301 242116
rect 260238 239869 260298 242115
rect 260235 239868 260301 239869
rect 260235 239804 260236 239868
rect 260300 239804 260301 239868
rect 260235 239803 260301 239804
rect 259867 239732 259933 239733
rect 259867 239668 259868 239732
rect 259932 239668 259933 239732
rect 259867 239667 259933 239668
rect 259683 237828 259749 237829
rect 259683 237764 259684 237828
rect 259748 237764 259749 237828
rect 259683 237763 259749 237764
rect 260238 229110 260298 239803
rect 260606 239461 260666 264283
rect 262811 258772 262877 258773
rect 262811 258708 262812 258772
rect 262876 258708 262877 258772
rect 262811 258707 262877 258708
rect 260971 253196 261037 253197
rect 260971 253132 260972 253196
rect 261036 253132 261037 253196
rect 260971 253131 261037 253132
rect 260787 243812 260853 243813
rect 260787 243748 260788 243812
rect 260852 243748 260853 243812
rect 260787 243747 260853 243748
rect 260790 239733 260850 243747
rect 260974 239733 261034 253131
rect 262259 249116 262325 249117
rect 262259 249052 262260 249116
rect 262324 249052 262325 249116
rect 262259 249051 262325 249052
rect 261523 240004 261589 240005
rect 261523 239940 261524 240004
rect 261588 239940 261589 240004
rect 261523 239939 261589 239940
rect 260787 239732 260853 239733
rect 260787 239668 260788 239732
rect 260852 239668 260853 239732
rect 260787 239667 260853 239668
rect 260971 239732 261037 239733
rect 260971 239668 260972 239732
rect 261036 239668 261037 239732
rect 260971 239667 261037 239668
rect 260603 239460 260669 239461
rect 260603 239396 260604 239460
rect 260668 239396 260669 239460
rect 260603 239395 260669 239396
rect 260974 238917 261034 239667
rect 261339 239460 261405 239461
rect 261339 239396 261340 239460
rect 261404 239396 261405 239460
rect 261339 239395 261405 239396
rect 260971 238916 261037 238917
rect 260971 238852 260972 238916
rect 261036 238852 261037 238916
rect 260971 238851 261037 238852
rect 260603 237828 260669 237829
rect 260603 237764 260604 237828
rect 260668 237764 260669 237828
rect 260603 237763 260669 237764
rect 260419 237420 260485 237421
rect 260419 237356 260420 237420
rect 260484 237356 260485 237420
rect 260419 237355 260485 237356
rect 259318 229050 259562 229110
rect 259686 229050 260298 229110
rect 259131 227628 259197 227629
rect 259131 227564 259132 227628
rect 259196 227564 259197 227628
rect 259131 227563 259197 227564
rect 259134 226405 259194 227563
rect 259131 226404 259197 226405
rect 259131 226340 259132 226404
rect 259196 226340 259197 226404
rect 259131 226339 259197 226340
rect 258395 222052 258461 222053
rect 258395 221988 258396 222052
rect 258460 221988 258461 222052
rect 258395 221987 258461 221988
rect 259131 222052 259197 222053
rect 259131 221988 259132 222052
rect 259196 221988 259197 222052
rect 259131 221987 259197 221988
rect 259134 221101 259194 221987
rect 259131 221100 259197 221101
rect 259131 221036 259132 221100
rect 259196 221036 259197 221100
rect 259131 221035 259197 221036
rect 259318 216341 259378 229050
rect 259315 216340 259381 216341
rect 259315 216276 259316 216340
rect 259380 216276 259381 216340
rect 259315 216275 259381 216276
rect 259318 215389 259378 216275
rect 259315 215388 259381 215389
rect 259315 215324 259316 215388
rect 259380 215324 259381 215388
rect 259315 215323 259381 215324
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 259686 143037 259746 229050
rect 260422 225861 260482 237355
rect 260419 225860 260485 225861
rect 260419 225796 260420 225860
rect 260484 225796 260485 225860
rect 260419 225795 260485 225796
rect 260422 219450 260482 225795
rect 260606 223549 260666 237763
rect 260603 223548 260669 223549
rect 260603 223484 260604 223548
rect 260668 223484 260669 223548
rect 260603 223483 260669 223484
rect 260054 219390 260482 219450
rect 260054 146165 260114 219390
rect 260051 146164 260117 146165
rect 260051 146100 260052 146164
rect 260116 146100 260117 146164
rect 260051 146099 260117 146100
rect 259683 143036 259749 143037
rect 259683 142972 259684 143036
rect 259748 142972 259749 143036
rect 259683 142971 259749 142972
rect 261342 142221 261402 239395
rect 261526 142901 261586 239939
rect 262262 239733 262322 249051
rect 262443 246260 262509 246261
rect 262443 246196 262444 246260
rect 262508 246196 262509 246260
rect 262443 246195 262509 246196
rect 262259 239732 262325 239733
rect 262259 239668 262260 239732
rect 262324 239668 262325 239732
rect 262259 239667 262325 239668
rect 262446 238917 262506 246195
rect 262814 240005 262874 258707
rect 264467 250476 264533 250477
rect 264467 250412 264468 250476
rect 264532 250412 264533 250476
rect 264467 250411 264533 250412
rect 263731 242724 263797 242725
rect 263731 242660 263732 242724
rect 263796 242660 263797 242724
rect 263731 242659 263797 242660
rect 262811 240004 262877 240005
rect 262811 239940 262812 240004
rect 262876 239940 262877 240004
rect 262811 239939 262877 239940
rect 262627 239868 262693 239869
rect 262627 239804 262628 239868
rect 262692 239804 262693 239868
rect 262627 239803 262693 239804
rect 262443 238916 262509 238917
rect 262443 238852 262444 238916
rect 262508 238852 262509 238916
rect 262443 238851 262509 238852
rect 262075 236876 262141 236877
rect 262075 236812 262076 236876
rect 262140 236812 262141 236876
rect 262075 236811 262141 236812
rect 262078 229110 262138 236811
rect 261710 229050 262138 229110
rect 261710 225997 261770 229050
rect 261707 225996 261773 225997
rect 261707 225932 261708 225996
rect 261772 225932 261773 225996
rect 261707 225931 261773 225932
rect 261710 143309 261770 225931
rect 262446 144669 262506 238851
rect 262630 237965 262690 239803
rect 263179 239460 263245 239461
rect 263179 239396 263180 239460
rect 263244 239396 263245 239460
rect 263179 239395 263245 239396
rect 262627 237964 262693 237965
rect 262627 237900 262628 237964
rect 262692 237900 262693 237964
rect 262627 237899 262693 237900
rect 262630 236741 262690 237899
rect 262627 236740 262693 236741
rect 262627 236676 262628 236740
rect 262692 236676 262693 236740
rect 262627 236675 262693 236676
rect 263182 229110 263242 239395
rect 263734 238237 263794 242659
rect 264470 239053 264530 250411
rect 264835 245036 264901 245037
rect 264835 244972 264836 245036
rect 264900 244972 264901 245036
rect 264835 244971 264901 244972
rect 264651 242044 264717 242045
rect 264651 241980 264652 242044
rect 264716 241980 264717 242044
rect 264651 241979 264717 241980
rect 264654 239869 264714 241979
rect 264651 239868 264717 239869
rect 264651 239804 264652 239868
rect 264716 239804 264717 239868
rect 264651 239803 264717 239804
rect 264099 239052 264165 239053
rect 264099 238988 264100 239052
rect 264164 238988 264165 239052
rect 264099 238987 264165 238988
rect 264467 239052 264533 239053
rect 264467 238988 264468 239052
rect 264532 238988 264533 239052
rect 264467 238987 264533 238988
rect 263731 238236 263797 238237
rect 263731 238172 263732 238236
rect 263796 238172 263797 238236
rect 263731 238171 263797 238172
rect 263182 229050 263426 229110
rect 263366 223277 263426 229050
rect 263363 223276 263429 223277
rect 263363 223212 263364 223276
rect 263428 223212 263429 223276
rect 263363 223211 263429 223212
rect 262443 144668 262509 144669
rect 262443 144604 262444 144668
rect 262508 144604 262509 144668
rect 262443 144603 262509 144604
rect 261707 143308 261773 143309
rect 261707 143244 261708 143308
rect 261772 143244 261773 143308
rect 261707 143243 261773 143244
rect 264102 142901 264162 238987
rect 264838 238645 264898 244971
rect 265022 244290 265082 271083
rect 267595 264212 267661 264213
rect 267595 264148 267596 264212
rect 267660 264148 267661 264212
rect 267595 264147 267661 264148
rect 266123 244900 266189 244901
rect 266123 244836 266124 244900
rect 266188 244836 266189 244900
rect 266123 244835 266189 244836
rect 265022 244230 265266 244290
rect 265019 243540 265085 243541
rect 265019 243476 265020 243540
rect 265084 243476 265085 243540
rect 265019 243475 265085 243476
rect 265022 239053 265082 243475
rect 265019 239052 265085 239053
rect 265019 238988 265020 239052
rect 265084 238988 265085 239052
rect 265019 238987 265085 238988
rect 265206 238781 265266 244230
rect 265939 242860 266005 242861
rect 265939 242796 265940 242860
rect 266004 242796 266005 242860
rect 265939 242795 266005 242796
rect 265755 241772 265821 241773
rect 265755 241708 265756 241772
rect 265820 241708 265821 241772
rect 265755 241707 265821 241708
rect 265387 240684 265453 240685
rect 265387 240620 265388 240684
rect 265452 240620 265453 240684
rect 265387 240619 265453 240620
rect 265390 239869 265450 240619
rect 265758 239869 265818 241707
rect 265387 239868 265453 239869
rect 265387 239804 265388 239868
rect 265452 239804 265453 239868
rect 265387 239803 265453 239804
rect 265755 239868 265821 239869
rect 265755 239804 265756 239868
rect 265820 239804 265821 239868
rect 265755 239803 265821 239804
rect 265203 238780 265269 238781
rect 265203 238716 265204 238780
rect 265268 238716 265269 238780
rect 265203 238715 265269 238716
rect 264835 238644 264901 238645
rect 264835 238580 264836 238644
rect 264900 238580 264901 238644
rect 264835 238579 264901 238580
rect 264283 238508 264349 238509
rect 264283 238444 264284 238508
rect 264348 238444 264349 238508
rect 264283 238443 264349 238444
rect 264286 147389 264346 238443
rect 265942 237693 266002 242795
rect 266126 239869 266186 244835
rect 267411 243132 267477 243133
rect 267411 243068 267412 243132
rect 267476 243068 267477 243132
rect 267411 243067 267477 243068
rect 266307 240004 266373 240005
rect 266307 239940 266308 240004
rect 266372 239940 266373 240004
rect 266307 239939 266373 239940
rect 266123 239868 266189 239869
rect 266123 239804 266124 239868
rect 266188 239804 266189 239868
rect 266123 239803 266189 239804
rect 266126 239325 266186 239803
rect 266310 239733 266370 239939
rect 266307 239732 266373 239733
rect 266307 239668 266308 239732
rect 266372 239668 266373 239732
rect 266307 239667 266373 239668
rect 267414 239325 267474 243067
rect 267598 239869 267658 264147
rect 269622 240413 269682 300051
rect 269619 240412 269685 240413
rect 269619 240348 269620 240412
rect 269684 240348 269685 240412
rect 269619 240347 269685 240348
rect 267595 239868 267661 239869
rect 267595 239804 267596 239868
rect 267660 239804 267661 239868
rect 267595 239803 267661 239804
rect 266123 239324 266189 239325
rect 266123 239260 266124 239324
rect 266188 239260 266189 239324
rect 266123 239259 266189 239260
rect 267411 239324 267477 239325
rect 267411 239260 267412 239324
rect 267476 239260 267477 239324
rect 267411 239259 267477 239260
rect 266307 238508 266373 238509
rect 266307 238444 266308 238508
rect 266372 238444 266373 238508
rect 266307 238443 266373 238444
rect 265939 237692 266005 237693
rect 265939 237628 265940 237692
rect 266004 237628 266005 237692
rect 265939 237627 266005 237628
rect 266310 175949 266370 238443
rect 267779 237828 267845 237829
rect 267779 237764 267780 237828
rect 267844 237764 267845 237828
rect 267779 237763 267845 237764
rect 266307 175948 266373 175949
rect 266307 175884 266308 175948
rect 266372 175884 266373 175948
rect 266307 175883 266373 175884
rect 264283 147388 264349 147389
rect 264283 147324 264284 147388
rect 264348 147324 264349 147388
rect 264283 147323 264349 147324
rect 267782 145757 267842 237763
rect 268331 237284 268397 237285
rect 268331 237220 268332 237284
rect 268396 237220 268397 237284
rect 268331 237219 268397 237220
rect 268334 155821 268394 237219
rect 270358 236741 270418 308483
rect 271091 307188 271157 307189
rect 271091 307124 271092 307188
rect 271156 307124 271157 307188
rect 271091 307123 271157 307124
rect 271094 240141 271154 307123
rect 271275 300252 271341 300253
rect 271275 300188 271276 300252
rect 271340 300188 271341 300252
rect 271275 300187 271341 300188
rect 271091 240140 271157 240141
rect 271091 240076 271092 240140
rect 271156 240076 271157 240140
rect 271091 240075 271157 240076
rect 270355 236740 270421 236741
rect 270355 236676 270356 236740
rect 270420 236676 270421 236740
rect 270355 236675 270421 236676
rect 271278 230213 271338 300187
rect 279374 290733 279434 375395
rect 280475 373012 280541 373013
rect 280475 372948 280476 373012
rect 280540 372948 280541 373012
rect 280475 372947 280541 372948
rect 279923 372740 279989 372741
rect 279923 372676 279924 372740
rect 279988 372676 279989 372740
rect 279923 372675 279989 372676
rect 279555 371516 279621 371517
rect 279555 371452 279556 371516
rect 279620 371452 279621 371516
rect 279555 371451 279621 371452
rect 279558 322285 279618 371451
rect 279926 359413 279986 372675
rect 280478 366349 280538 372947
rect 280659 372332 280725 372333
rect 280659 372268 280660 372332
rect 280724 372268 280725 372332
rect 280659 372267 280725 372268
rect 280475 366348 280541 366349
rect 280475 366284 280476 366348
rect 280540 366284 280541 366348
rect 280475 366283 280541 366284
rect 280662 361045 280722 372267
rect 280659 361044 280725 361045
rect 280659 360980 280660 361044
rect 280724 360980 280725 361044
rect 280659 360979 280725 360980
rect 279923 359412 279989 359413
rect 279923 359348 279924 359412
rect 279988 359348 279989 359412
rect 279923 359347 279989 359348
rect 280659 359412 280725 359413
rect 280659 359348 280660 359412
rect 280724 359348 280725 359412
rect 280659 359347 280725 359348
rect 279555 322284 279621 322285
rect 279555 322220 279556 322284
rect 279620 322220 279621 322284
rect 279555 322219 279621 322220
rect 279371 290732 279437 290733
rect 279371 290668 279372 290732
rect 279436 290668 279437 290732
rect 279371 290667 279437 290668
rect 273851 242044 273917 242045
rect 273851 241980 273852 242044
rect 273916 241980 273917 242044
rect 273851 241979 273917 241980
rect 273854 241773 273914 241979
rect 273851 241772 273917 241773
rect 273851 241708 273852 241772
rect 273916 241708 273917 241772
rect 273851 241707 273917 241708
rect 271827 241636 271893 241637
rect 271827 241572 271828 241636
rect 271892 241572 271893 241636
rect 271827 241571 271893 241572
rect 271830 239733 271890 241571
rect 271827 239732 271893 239733
rect 271827 239668 271828 239732
rect 271892 239668 271893 239732
rect 271827 239667 271893 239668
rect 271275 230212 271341 230213
rect 271275 230148 271276 230212
rect 271340 230148 271341 230212
rect 271275 230147 271341 230148
rect 268331 155820 268397 155821
rect 268331 155756 268332 155820
rect 268396 155756 268397 155820
rect 268331 155755 268397 155756
rect 267779 145756 267845 145757
rect 267779 145692 267780 145756
rect 267844 145692 267845 145756
rect 267779 145691 267845 145692
rect 261523 142900 261589 142901
rect 261523 142836 261524 142900
rect 261588 142836 261589 142900
rect 261523 142835 261589 142836
rect 264099 142900 264165 142901
rect 264099 142836 264100 142900
rect 264164 142836 264165 142900
rect 264099 142835 264165 142836
rect 261339 142220 261405 142221
rect 261339 142156 261340 142220
rect 261404 142156 261405 142220
rect 261339 142155 261405 142156
rect 271830 136645 271890 239667
rect 273854 154325 273914 241707
rect 273851 154324 273917 154325
rect 273851 154260 273852 154324
rect 273916 154260 273917 154324
rect 273851 154259 273917 154260
rect 271827 136644 271893 136645
rect 271827 136580 271828 136644
rect 271892 136580 271893 136644
rect 271827 136579 271893 136580
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 280662 71909 280722 359347
rect 281398 316981 281458 387091
rect 282870 379530 282930 391987
rect 282870 379470 283114 379530
rect 282683 371380 282749 371381
rect 282683 371316 282684 371380
rect 282748 371316 282749 371380
rect 282683 371315 282749 371316
rect 282131 369748 282197 369749
rect 282131 369684 282132 369748
rect 282196 369684 282197 369748
rect 282131 369683 282197 369684
rect 281579 369476 281645 369477
rect 281579 369412 281580 369476
rect 281644 369412 281645 369476
rect 281579 369411 281645 369412
rect 281582 361861 281642 369411
rect 281579 361860 281645 361861
rect 281579 361796 281580 361860
rect 281644 361796 281645 361860
rect 281579 361795 281645 361796
rect 282134 360909 282194 369683
rect 282686 369477 282746 371315
rect 282683 369476 282749 369477
rect 282683 369412 282684 369476
rect 282748 369412 282749 369476
rect 282683 369411 282749 369412
rect 282131 360908 282197 360909
rect 282131 360844 282132 360908
rect 282196 360844 282197 360908
rect 282131 360843 282197 360844
rect 283054 360210 283114 379470
rect 282870 360150 283114 360210
rect 282870 331230 282930 360150
rect 282686 331170 282930 331230
rect 282686 321877 282746 331170
rect 283422 328470 283482 397155
rect 288019 388924 288085 388925
rect 288019 388860 288020 388924
rect 288084 388860 288085 388924
rect 288019 388859 288085 388860
rect 287467 388788 287533 388789
rect 287467 388724 287468 388788
rect 287532 388724 287533 388788
rect 287467 388723 287533 388724
rect 286731 388244 286797 388245
rect 286731 388180 286732 388244
rect 286796 388180 286797 388244
rect 286731 388179 286797 388180
rect 286363 381716 286429 381717
rect 286363 381652 286364 381716
rect 286428 381652 286429 381716
rect 286363 381651 286429 381652
rect 285075 376820 285141 376821
rect 285075 376756 285076 376820
rect 285140 376756 285141 376820
rect 285075 376755 285141 376756
rect 283422 328410 284034 328470
rect 282683 321876 282749 321877
rect 282683 321812 282684 321876
rect 282748 321812 282749 321876
rect 282683 321811 282749 321812
rect 282683 321604 282749 321605
rect 282683 321540 282684 321604
rect 282748 321540 282749 321604
rect 282683 321539 282749 321540
rect 282686 320789 282746 321539
rect 283235 321060 283301 321061
rect 283235 320996 283236 321060
rect 283300 320996 283301 321060
rect 283235 320995 283301 320996
rect 282683 320788 282749 320789
rect 282683 320724 282684 320788
rect 282748 320724 282749 320788
rect 282683 320723 282749 320724
rect 283238 319021 283298 320995
rect 283974 320789 284034 328410
rect 284339 321876 284405 321877
rect 284339 321812 284340 321876
rect 284404 321812 284405 321876
rect 284339 321811 284405 321812
rect 283971 320788 284037 320789
rect 283971 320724 283972 320788
rect 284036 320724 284037 320788
rect 283971 320723 284037 320724
rect 283787 320108 283853 320109
rect 283787 320044 283788 320108
rect 283852 320044 283853 320108
rect 283787 320043 283853 320044
rect 283603 319972 283669 319973
rect 283603 319908 283604 319972
rect 283668 319908 283669 319972
rect 283603 319907 283669 319908
rect 283419 319292 283485 319293
rect 283419 319228 283420 319292
rect 283484 319228 283485 319292
rect 283419 319227 283485 319228
rect 283235 319020 283301 319021
rect 283235 318956 283236 319020
rect 283300 318956 283301 319020
rect 283235 318955 283301 318956
rect 283422 318749 283482 319227
rect 283606 319021 283666 319907
rect 283790 319429 283850 320043
rect 283787 319428 283853 319429
rect 283787 319364 283788 319428
rect 283852 319364 283853 319428
rect 283787 319363 283853 319364
rect 283974 319293 284034 320723
rect 284342 319973 284402 321811
rect 284523 321604 284589 321605
rect 284523 321540 284524 321604
rect 284588 321540 284589 321604
rect 284523 321539 284589 321540
rect 284526 320109 284586 321539
rect 285078 320789 285138 376755
rect 285259 369884 285325 369885
rect 285259 369820 285260 369884
rect 285324 369820 285325 369884
rect 285259 369819 285325 369820
rect 285262 368797 285322 369819
rect 285259 368796 285325 368797
rect 285259 368732 285260 368796
rect 285324 368732 285325 368796
rect 285259 368731 285325 368732
rect 286366 321605 286426 381651
rect 286547 369476 286613 369477
rect 286547 369412 286548 369476
rect 286612 369412 286613 369476
rect 286547 369411 286613 369412
rect 286363 321604 286429 321605
rect 286363 321540 286364 321604
rect 286428 321540 286429 321604
rect 286363 321539 286429 321540
rect 285075 320788 285141 320789
rect 285075 320724 285076 320788
rect 285140 320724 285141 320788
rect 285075 320723 285141 320724
rect 284707 320652 284773 320653
rect 284707 320588 284708 320652
rect 284772 320588 284773 320652
rect 284707 320587 284773 320588
rect 284891 320652 284957 320653
rect 284891 320588 284892 320652
rect 284956 320588 284957 320652
rect 284891 320587 284957 320588
rect 284523 320108 284589 320109
rect 284523 320044 284524 320108
rect 284588 320044 284589 320108
rect 284523 320043 284589 320044
rect 284339 319972 284405 319973
rect 284339 319908 284340 319972
rect 284404 319908 284405 319972
rect 284339 319907 284405 319908
rect 283971 319292 284037 319293
rect 283971 319228 283972 319292
rect 284036 319228 284037 319292
rect 283971 319227 284037 319228
rect 283603 319020 283669 319021
rect 283603 318956 283604 319020
rect 283668 318956 283669 319020
rect 283603 318955 283669 318956
rect 283419 318748 283485 318749
rect 283419 318684 283420 318748
rect 283484 318684 283485 318748
rect 283419 318683 283485 318684
rect 284526 317933 284586 320043
rect 284710 319021 284770 320587
rect 284894 319021 284954 320587
rect 285078 319701 285138 320723
rect 286550 320245 286610 369411
rect 286547 320244 286613 320245
rect 286547 320180 286548 320244
rect 286612 320180 286613 320244
rect 286547 320179 286613 320180
rect 285627 320108 285693 320109
rect 285627 320044 285628 320108
rect 285692 320044 285693 320108
rect 285627 320043 285693 320044
rect 285075 319700 285141 319701
rect 285075 319636 285076 319700
rect 285140 319636 285141 319700
rect 285075 319635 285141 319636
rect 285630 319293 285690 320043
rect 285627 319292 285693 319293
rect 285627 319228 285628 319292
rect 285692 319228 285693 319292
rect 285627 319227 285693 319228
rect 284707 319020 284773 319021
rect 284707 318956 284708 319020
rect 284772 318956 284773 319020
rect 284707 318955 284773 318956
rect 284891 319020 284957 319021
rect 284891 318956 284892 319020
rect 284956 318956 284957 319020
rect 284891 318955 284957 318956
rect 285811 318340 285877 318341
rect 285811 318276 285812 318340
rect 285876 318276 285877 318340
rect 285811 318275 285877 318276
rect 285627 318068 285693 318069
rect 285627 318004 285628 318068
rect 285692 318004 285693 318068
rect 285627 318003 285693 318004
rect 284523 317932 284589 317933
rect 284523 317868 284524 317932
rect 284588 317868 284589 317932
rect 284523 317867 284589 317868
rect 283051 317524 283117 317525
rect 283051 317460 283052 317524
rect 283116 317460 283117 317524
rect 283051 317459 283117 317460
rect 284339 317524 284405 317525
rect 284339 317460 284340 317524
rect 284404 317460 284405 317524
rect 284339 317459 284405 317460
rect 281395 316980 281461 316981
rect 281395 316916 281396 316980
rect 281460 316916 281461 316980
rect 281395 316915 281461 316916
rect 281398 307733 281458 316915
rect 283054 311910 283114 317459
rect 282870 311850 283114 311910
rect 281395 307732 281461 307733
rect 281395 307668 281396 307732
rect 281460 307668 281461 307732
rect 281395 307667 281461 307668
rect 282870 307597 282930 311850
rect 284342 309093 284402 317459
rect 284339 309092 284405 309093
rect 284339 309028 284340 309092
rect 284404 309028 284405 309092
rect 284339 309027 284405 309028
rect 282867 307596 282933 307597
rect 282867 307532 282868 307596
rect 282932 307532 282933 307596
rect 282867 307531 282933 307532
rect 285630 296581 285690 318003
rect 285627 296580 285693 296581
rect 285627 296516 285628 296580
rect 285692 296516 285693 296580
rect 285627 296515 285693 296516
rect 285814 296445 285874 318275
rect 286550 318069 286610 320179
rect 286734 320109 286794 388179
rect 287283 369476 287349 369477
rect 287283 369412 287284 369476
rect 287348 369412 287349 369476
rect 287283 369411 287349 369412
rect 287286 368525 287346 369411
rect 287283 368524 287349 368525
rect 287283 368460 287284 368524
rect 287348 368460 287349 368524
rect 287283 368459 287349 368460
rect 287470 320789 287530 388723
rect 287835 387564 287901 387565
rect 287835 387500 287836 387564
rect 287900 387500 287901 387564
rect 287835 387499 287901 387500
rect 287467 320788 287533 320789
rect 287467 320724 287468 320788
rect 287532 320724 287533 320788
rect 287467 320723 287533 320724
rect 287467 320652 287533 320653
rect 287467 320588 287468 320652
rect 287532 320588 287533 320652
rect 287467 320587 287533 320588
rect 287283 320244 287349 320245
rect 287283 320180 287284 320244
rect 287348 320180 287349 320244
rect 287283 320179 287349 320180
rect 286731 320108 286797 320109
rect 286731 320044 286732 320108
rect 286796 320044 286797 320108
rect 286731 320043 286797 320044
rect 286915 320108 286981 320109
rect 286915 320044 286916 320108
rect 286980 320044 286981 320108
rect 286915 320043 286981 320044
rect 286918 319293 286978 320043
rect 286915 319292 286981 319293
rect 286915 319228 286916 319292
rect 286980 319228 286981 319292
rect 286915 319227 286981 319228
rect 287286 319021 287346 320179
rect 287470 319701 287530 320587
rect 287651 320108 287717 320109
rect 287651 320044 287652 320108
rect 287716 320044 287717 320108
rect 287651 320043 287717 320044
rect 287467 319700 287533 319701
rect 287467 319636 287468 319700
rect 287532 319636 287533 319700
rect 287467 319635 287533 319636
rect 287283 319020 287349 319021
rect 287283 318956 287284 319020
rect 287348 318956 287349 319020
rect 287283 318955 287349 318956
rect 286547 318068 286613 318069
rect 286547 318004 286548 318068
rect 286612 318004 286613 318068
rect 286547 318003 286613 318004
rect 287099 317932 287165 317933
rect 287099 317868 287100 317932
rect 287164 317868 287165 317932
rect 287099 317867 287165 317868
rect 285811 296444 285877 296445
rect 285811 296380 285812 296444
rect 285876 296380 285877 296444
rect 285811 296379 285877 296380
rect 287102 257549 287162 317867
rect 287654 317389 287714 320043
rect 287838 318749 287898 387499
rect 288022 319701 288082 388859
rect 288755 378724 288821 378725
rect 288755 378660 288756 378724
rect 288820 378660 288821 378724
rect 288755 378659 288821 378660
rect 288571 321876 288637 321877
rect 288571 321812 288572 321876
rect 288636 321812 288637 321876
rect 288571 321811 288637 321812
rect 288574 321194 288634 321811
rect 288390 321134 288634 321194
rect 288390 320925 288450 321134
rect 288571 321060 288637 321061
rect 288571 320996 288572 321060
rect 288636 320996 288637 321060
rect 288571 320995 288637 320996
rect 288387 320924 288453 320925
rect 288387 320860 288388 320924
rect 288452 320860 288453 320924
rect 288387 320859 288453 320860
rect 288574 320789 288634 320995
rect 288203 320788 288269 320789
rect 288203 320724 288204 320788
rect 288268 320724 288269 320788
rect 288203 320723 288269 320724
rect 288571 320788 288637 320789
rect 288571 320724 288572 320788
rect 288636 320724 288637 320788
rect 288571 320723 288637 320724
rect 288019 319700 288085 319701
rect 288019 319636 288020 319700
rect 288084 319636 288085 319700
rect 288019 319635 288085 319636
rect 287835 318748 287901 318749
rect 287835 318684 287836 318748
rect 287900 318684 287901 318748
rect 287835 318683 287901 318684
rect 287651 317388 287717 317389
rect 287651 317324 287652 317388
rect 287716 317324 287717 317388
rect 287651 317323 287717 317324
rect 288206 314669 288266 320723
rect 288387 320244 288453 320245
rect 288387 320180 288388 320244
rect 288452 320180 288453 320244
rect 288387 320179 288453 320180
rect 288390 319293 288450 320179
rect 288571 319972 288637 319973
rect 288571 319908 288572 319972
rect 288636 319908 288637 319972
rect 288571 319907 288637 319908
rect 288574 319293 288634 319907
rect 288758 319701 288818 378659
rect 288939 369340 289005 369341
rect 288939 369276 288940 369340
rect 289004 369276 289005 369340
rect 288939 369275 289005 369276
rect 288942 368661 289002 369275
rect 288939 368660 289005 368661
rect 288939 368596 288940 368660
rect 289004 368596 289005 368660
rect 288939 368595 289005 368596
rect 288939 322012 289005 322013
rect 288939 321948 288940 322012
rect 289004 321948 289005 322012
rect 288939 321947 289005 321948
rect 288942 321333 289002 321947
rect 288939 321332 289005 321333
rect 288939 321268 288940 321332
rect 289004 321268 289005 321332
rect 288939 321267 289005 321268
rect 288939 320108 289005 320109
rect 288939 320044 288940 320108
rect 289004 320044 289005 320108
rect 288939 320043 289005 320044
rect 288755 319700 288821 319701
rect 288755 319636 288756 319700
rect 288820 319636 288821 319700
rect 288755 319635 288821 319636
rect 288387 319292 288453 319293
rect 288387 319228 288388 319292
rect 288452 319228 288453 319292
rect 288387 319227 288453 319228
rect 288571 319292 288637 319293
rect 288571 319228 288572 319292
rect 288636 319228 288637 319292
rect 288571 319227 288637 319228
rect 288387 317932 288453 317933
rect 288387 317868 288388 317932
rect 288452 317868 288453 317932
rect 288387 317867 288453 317868
rect 288203 314668 288269 314669
rect 288203 314604 288204 314668
rect 288268 314604 288269 314668
rect 288203 314603 288269 314604
rect 287099 257548 287165 257549
rect 287099 257484 287100 257548
rect 287164 257484 287165 257548
rect 287099 257483 287165 257484
rect 288390 241501 288450 317867
rect 288758 295221 288818 319635
rect 288942 319021 289002 320043
rect 288939 319020 289005 319021
rect 288939 318956 288940 319020
rect 289004 318956 289005 319020
rect 288939 318955 289005 318956
rect 289126 318069 289186 398923
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289491 388652 289557 388653
rect 289491 388588 289492 388652
rect 289556 388588 289557 388652
rect 289491 388587 289557 388588
rect 289307 378588 289373 378589
rect 289307 378524 289308 378588
rect 289372 378524 289373 378588
rect 289307 378523 289373 378524
rect 289310 320789 289370 378523
rect 289307 320788 289373 320789
rect 289307 320724 289308 320788
rect 289372 320724 289373 320788
rect 289307 320723 289373 320724
rect 289123 318068 289189 318069
rect 289123 318004 289124 318068
rect 289188 318004 289189 318068
rect 289123 318003 289189 318004
rect 288755 295220 288821 295221
rect 288755 295156 288756 295220
rect 288820 295156 288821 295220
rect 288755 295155 288821 295156
rect 289310 245445 289370 320723
rect 289494 320109 289554 388587
rect 289794 363454 290414 398898
rect 293514 705798 294134 705830
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 307707 404292 307773 404293
rect 307707 404228 307708 404292
rect 307772 404228 307773 404292
rect 307707 404227 307773 404228
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293171 392596 293237 392597
rect 293171 392532 293172 392596
rect 293236 392532 293237 392596
rect 293171 392531 293237 392532
rect 291699 389060 291765 389061
rect 291699 388996 291700 389060
rect 291764 388996 291765 389060
rect 291699 388995 291765 388996
rect 290963 379268 291029 379269
rect 290963 379204 290964 379268
rect 291028 379204 291029 379268
rect 290963 379203 291029 379204
rect 290779 378860 290845 378861
rect 290779 378796 290780 378860
rect 290844 378796 290845 378860
rect 290779 378795 290845 378796
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289491 320108 289557 320109
rect 289491 320044 289492 320108
rect 289556 320044 289557 320108
rect 289491 320043 289557 320044
rect 289794 291454 290414 326898
rect 290595 321604 290661 321605
rect 290595 321540 290596 321604
rect 290660 321540 290661 321604
rect 290595 321539 290661 321540
rect 290598 318885 290658 321539
rect 290782 319973 290842 378795
rect 290966 321197 291026 379203
rect 291331 379132 291397 379133
rect 291331 379068 291332 379132
rect 291396 379068 291397 379132
rect 291331 379067 291397 379068
rect 291147 321468 291213 321469
rect 291147 321404 291148 321468
rect 291212 321404 291213 321468
rect 291147 321403 291213 321404
rect 290963 321196 291029 321197
rect 290963 321132 290964 321196
rect 291028 321132 291029 321196
rect 290963 321131 291029 321132
rect 290779 319972 290845 319973
rect 290779 319908 290780 319972
rect 290844 319908 290845 319972
rect 290779 319907 290845 319908
rect 290779 319836 290845 319837
rect 290779 319772 290780 319836
rect 290844 319772 290845 319836
rect 290779 319771 290845 319772
rect 290595 318884 290661 318885
rect 290595 318820 290596 318884
rect 290660 318820 290661 318884
rect 290595 318819 290661 318820
rect 290595 318068 290661 318069
rect 290595 318004 290596 318068
rect 290660 318004 290661 318068
rect 290595 318003 290661 318004
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289307 245444 289373 245445
rect 289307 245380 289308 245444
rect 289372 245380 289373 245444
rect 289307 245379 289373 245380
rect 288387 241500 288453 241501
rect 288387 241436 288388 241500
rect 288452 241436 288453 241500
rect 288387 241435 288453 241436
rect 289794 219454 290414 254898
rect 290598 247893 290658 318003
rect 290782 317525 290842 319771
rect 290779 317524 290845 317525
rect 290779 317460 290780 317524
rect 290844 317460 290845 317524
rect 290779 317459 290845 317460
rect 290966 311910 291026 321131
rect 291150 320245 291210 321403
rect 291147 320244 291213 320245
rect 291147 320180 291148 320244
rect 291212 320180 291213 320244
rect 291147 320179 291213 320180
rect 291334 320109 291394 379067
rect 291331 320108 291397 320109
rect 291331 320044 291332 320108
rect 291396 320044 291397 320108
rect 291331 320043 291397 320044
rect 291147 319156 291213 319157
rect 291147 319092 291148 319156
rect 291212 319092 291213 319156
rect 291147 319091 291213 319092
rect 290782 311850 291026 311910
rect 290782 309773 290842 311850
rect 290779 309772 290845 309773
rect 290779 309708 290780 309772
rect 290844 309708 290845 309772
rect 290779 309707 290845 309708
rect 291150 294405 291210 319091
rect 291334 309909 291394 320043
rect 291702 317525 291762 388995
rect 292987 381580 293053 381581
rect 292987 381516 292988 381580
rect 293052 381516 293053 381580
rect 292987 381515 293053 381516
rect 291883 379404 291949 379405
rect 291883 379340 291884 379404
rect 291948 379340 291949 379404
rect 291883 379339 291949 379340
rect 291886 320789 291946 379339
rect 292251 378996 292317 378997
rect 292251 378932 292252 378996
rect 292316 378932 292317 378996
rect 292251 378931 292317 378932
rect 291883 320788 291949 320789
rect 291883 320724 291884 320788
rect 291948 320724 291949 320788
rect 291883 320723 291949 320724
rect 291699 317524 291765 317525
rect 291699 317460 291700 317524
rect 291764 317460 291765 317524
rect 291699 317459 291765 317460
rect 291699 311132 291765 311133
rect 291699 311068 291700 311132
rect 291764 311068 291765 311132
rect 291699 311067 291765 311068
rect 291331 309908 291397 309909
rect 291331 309844 291332 309908
rect 291396 309844 291397 309908
rect 291331 309843 291397 309844
rect 291147 294404 291213 294405
rect 291147 294340 291148 294404
rect 291212 294340 291213 294404
rect 291147 294339 291213 294340
rect 290595 247892 290661 247893
rect 290595 247828 290596 247892
rect 290660 247828 290661 247892
rect 290595 247827 290661 247828
rect 291702 220013 291762 311067
rect 291886 310997 291946 320723
rect 292254 320245 292314 378931
rect 292803 374780 292869 374781
rect 292803 374716 292804 374780
rect 292868 374716 292869 374780
rect 292803 374715 292869 374716
rect 292619 321332 292685 321333
rect 292619 321268 292620 321332
rect 292684 321268 292685 321332
rect 292619 321267 292685 321268
rect 292622 320789 292682 321267
rect 292619 320788 292685 320789
rect 292619 320724 292620 320788
rect 292684 320724 292685 320788
rect 292619 320723 292685 320724
rect 292435 320652 292501 320653
rect 292435 320588 292436 320652
rect 292500 320588 292501 320652
rect 292435 320587 292501 320588
rect 292251 320244 292317 320245
rect 292251 320180 292252 320244
rect 292316 320180 292317 320244
rect 292251 320179 292317 320180
rect 292067 320108 292133 320109
rect 292067 320044 292068 320108
rect 292132 320044 292133 320108
rect 292067 320043 292133 320044
rect 292070 318341 292130 320043
rect 292254 319157 292314 320179
rect 292251 319156 292317 319157
rect 292251 319092 292252 319156
rect 292316 319092 292317 319156
rect 292251 319091 292317 319092
rect 292067 318340 292133 318341
rect 292067 318276 292068 318340
rect 292132 318276 292133 318340
rect 292067 318275 292133 318276
rect 292438 318069 292498 320587
rect 292619 320108 292685 320109
rect 292619 320044 292620 320108
rect 292684 320044 292685 320108
rect 292619 320043 292685 320044
rect 292622 319293 292682 320043
rect 292619 319292 292685 319293
rect 292619 319228 292620 319292
rect 292684 319228 292685 319292
rect 292619 319227 292685 319228
rect 292806 318613 292866 374715
rect 292990 320245 293050 381515
rect 293174 320653 293234 392531
rect 293514 367174 294134 402618
rect 297219 394636 297285 394637
rect 297219 394572 297220 394636
rect 297284 394572 297285 394636
rect 297219 394571 297285 394572
rect 296483 394364 296549 394365
rect 296483 394300 296484 394364
rect 296548 394300 296549 394364
rect 296483 394299 296549 394300
rect 295011 391644 295077 391645
rect 295011 391580 295012 391644
rect 295076 391580 295077 391644
rect 295011 391579 295077 391580
rect 294643 390556 294709 390557
rect 294643 390492 294644 390556
rect 294708 390492 294709 390556
rect 294643 390491 294709 390492
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293355 322012 293421 322013
rect 293355 321948 293356 322012
rect 293420 321948 293421 322012
rect 293355 321947 293421 321948
rect 293358 321333 293418 321947
rect 293355 321332 293421 321333
rect 293355 321268 293356 321332
rect 293420 321268 293421 321332
rect 293355 321267 293421 321268
rect 293171 320652 293237 320653
rect 293171 320588 293172 320652
rect 293236 320588 293237 320652
rect 293171 320587 293237 320588
rect 292987 320244 293053 320245
rect 292987 320180 292988 320244
rect 293052 320180 293053 320244
rect 292987 320179 293053 320180
rect 292987 319972 293053 319973
rect 292987 319908 292988 319972
rect 293052 319908 293053 319972
rect 292987 319907 293053 319908
rect 292990 319293 293050 319907
rect 292987 319292 293053 319293
rect 292987 319228 292988 319292
rect 293052 319228 293053 319292
rect 292987 319227 293053 319228
rect 292803 318612 292869 318613
rect 292803 318548 292804 318612
rect 292868 318548 292869 318612
rect 292803 318547 292869 318548
rect 292435 318068 292501 318069
rect 292435 318004 292436 318068
rect 292500 318004 292501 318068
rect 292435 318003 292501 318004
rect 292435 317388 292501 317389
rect 292435 317324 292436 317388
rect 292500 317324 292501 317388
rect 292435 317323 292501 317324
rect 291883 310996 291949 310997
rect 291883 310932 291884 310996
rect 291948 310932 291949 310996
rect 291883 310931 291949 310932
rect 292438 299301 292498 317323
rect 292435 299300 292501 299301
rect 292435 299236 292436 299300
rect 292500 299236 292501 299300
rect 292435 299235 292501 299236
rect 293174 296730 293234 320587
rect 293355 320244 293421 320245
rect 293355 320180 293356 320244
rect 293420 320180 293421 320244
rect 293355 320179 293421 320180
rect 293358 313173 293418 320179
rect 293355 313172 293421 313173
rect 293355 313108 293356 313172
rect 293420 313108 293421 313172
rect 293355 313107 293421 313108
rect 292622 296670 293234 296730
rect 292622 240957 292682 296670
rect 293514 295174 294134 330618
rect 294275 321196 294341 321197
rect 294275 321132 294276 321196
rect 294340 321132 294341 321196
rect 294275 321131 294341 321132
rect 294278 320109 294338 321131
rect 294275 320108 294341 320109
rect 294275 320044 294276 320108
rect 294340 320044 294341 320108
rect 294275 320043 294341 320044
rect 294459 320108 294525 320109
rect 294459 320044 294460 320108
rect 294524 320044 294525 320108
rect 294459 320043 294525 320044
rect 294278 312629 294338 320043
rect 294275 312628 294341 312629
rect 294275 312564 294276 312628
rect 294340 312564 294341 312628
rect 294275 312563 294341 312564
rect 294462 312493 294522 320043
rect 294646 318749 294706 390491
rect 295014 321197 295074 391579
rect 295195 391100 295261 391101
rect 295195 391036 295196 391100
rect 295260 391036 295261 391100
rect 295195 391035 295261 391036
rect 295011 321196 295077 321197
rect 295011 321132 295012 321196
rect 295076 321132 295077 321196
rect 295011 321131 295077 321132
rect 294827 320244 294893 320245
rect 294827 320180 294828 320244
rect 294892 320180 294893 320244
rect 294827 320179 294893 320180
rect 295011 320244 295077 320245
rect 295011 320180 295012 320244
rect 295076 320180 295077 320244
rect 295011 320179 295077 320180
rect 294830 319429 294890 320179
rect 294827 319428 294893 319429
rect 294827 319364 294828 319428
rect 294892 319364 294893 319428
rect 294827 319363 294893 319364
rect 295014 319293 295074 320179
rect 295198 320109 295258 391035
rect 296299 376004 296365 376005
rect 296299 375940 296300 376004
rect 296364 375940 296365 376004
rect 296299 375939 296365 375940
rect 295563 320652 295629 320653
rect 295563 320588 295564 320652
rect 295628 320588 295629 320652
rect 295563 320587 295629 320588
rect 295195 320108 295261 320109
rect 295195 320044 295196 320108
rect 295260 320044 295261 320108
rect 295195 320043 295261 320044
rect 295379 320108 295445 320109
rect 295379 320044 295380 320108
rect 295444 320044 295445 320108
rect 295379 320043 295445 320044
rect 295195 319836 295261 319837
rect 295195 319772 295196 319836
rect 295260 319772 295261 319836
rect 295195 319771 295261 319772
rect 295011 319292 295077 319293
rect 295011 319228 295012 319292
rect 295076 319228 295077 319292
rect 295011 319227 295077 319228
rect 295198 318885 295258 319771
rect 295382 319293 295442 320043
rect 295566 319429 295626 320587
rect 296302 320245 296362 375939
rect 295747 320244 295813 320245
rect 295747 320180 295748 320244
rect 295812 320180 295813 320244
rect 295747 320179 295813 320180
rect 296299 320244 296365 320245
rect 296299 320180 296300 320244
rect 296364 320180 296365 320244
rect 296299 320179 296365 320180
rect 295563 319428 295629 319429
rect 295563 319364 295564 319428
rect 295628 319364 295629 319428
rect 295563 319363 295629 319364
rect 295379 319292 295445 319293
rect 295379 319228 295380 319292
rect 295444 319228 295445 319292
rect 295379 319227 295445 319228
rect 295750 319021 295810 320179
rect 295747 319020 295813 319021
rect 295747 318956 295748 319020
rect 295812 318956 295813 319020
rect 295747 318955 295813 318956
rect 295195 318884 295261 318885
rect 295195 318820 295196 318884
rect 295260 318820 295261 318884
rect 295195 318819 295261 318820
rect 294643 318748 294709 318749
rect 294643 318684 294644 318748
rect 294708 318684 294709 318748
rect 294643 318683 294709 318684
rect 294646 312765 294706 318683
rect 296302 315757 296362 320179
rect 296486 320109 296546 394299
rect 297222 320789 297282 394571
rect 297955 394500 298021 394501
rect 297955 394436 297956 394500
rect 298020 394436 298021 394500
rect 297955 394435 298021 394436
rect 297587 387428 297653 387429
rect 297587 387364 297588 387428
rect 297652 387364 297653 387428
rect 297587 387363 297653 387364
rect 297403 374644 297469 374645
rect 297403 374580 297404 374644
rect 297468 374580 297469 374644
rect 297403 374579 297469 374580
rect 297219 320788 297285 320789
rect 297219 320724 297220 320788
rect 297284 320724 297285 320788
rect 297219 320723 297285 320724
rect 296483 320108 296549 320109
rect 296483 320044 296484 320108
rect 296548 320044 296549 320108
rect 296483 320043 296549 320044
rect 296851 320108 296917 320109
rect 296851 320044 296852 320108
rect 296916 320044 296917 320108
rect 296851 320043 296917 320044
rect 296486 315893 296546 320043
rect 296667 318748 296733 318749
rect 296667 318684 296668 318748
rect 296732 318684 296733 318748
rect 296667 318683 296733 318684
rect 296483 315892 296549 315893
rect 296483 315828 296484 315892
rect 296548 315828 296549 315892
rect 296483 315827 296549 315828
rect 296299 315756 296365 315757
rect 296299 315692 296300 315756
rect 296364 315692 296365 315756
rect 296299 315691 296365 315692
rect 294643 312764 294709 312765
rect 294643 312700 294644 312764
rect 294708 312700 294709 312764
rect 294643 312699 294709 312700
rect 294459 312492 294525 312493
rect 294459 312428 294460 312492
rect 294524 312428 294525 312492
rect 294459 312427 294525 312428
rect 296670 311910 296730 318683
rect 296854 318477 296914 320043
rect 297222 318810 297282 320723
rect 297406 319021 297466 374579
rect 297590 320109 297650 387363
rect 297587 320108 297653 320109
rect 297587 320044 297588 320108
rect 297652 320044 297653 320108
rect 297587 320043 297653 320044
rect 297771 320108 297837 320109
rect 297771 320044 297772 320108
rect 297836 320044 297837 320108
rect 297771 320043 297837 320044
rect 297403 319020 297469 319021
rect 297403 318956 297404 319020
rect 297468 318956 297469 319020
rect 297403 318955 297469 318956
rect 297038 318750 297282 318810
rect 296851 318476 296917 318477
rect 296851 318412 296852 318476
rect 296916 318412 296917 318476
rect 296851 318411 296917 318412
rect 297038 315621 297098 318750
rect 297035 315620 297101 315621
rect 297035 315556 297036 315620
rect 297100 315556 297101 315620
rect 297035 315555 297101 315556
rect 297406 315485 297466 318955
rect 297403 315484 297469 315485
rect 297403 315420 297404 315484
rect 297468 315420 297469 315484
rect 297403 315419 297469 315420
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 292619 240956 292685 240957
rect 292619 240892 292620 240956
rect 292684 240892 292685 240956
rect 292619 240891 292685 240892
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 291699 220012 291765 220013
rect 291699 219948 291700 220012
rect 291764 219948 291765 220012
rect 291699 219947 291765 219948
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 280659 71908 280725 71909
rect 280659 71844 280660 71908
rect 280724 71844 280725 71908
rect 280659 71843 280725 71844
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -1894 258134 -1862
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 187174 294134 222618
rect 296486 311850 296730 311910
rect 296486 219450 296546 311850
rect 297590 310453 297650 320043
rect 297774 319021 297834 320043
rect 297958 319429 298018 394435
rect 299243 393276 299309 393277
rect 299243 393212 299244 393276
rect 299308 393212 299309 393276
rect 299243 393211 299309 393212
rect 298875 384436 298941 384437
rect 298875 384372 298876 384436
rect 298940 384372 298941 384436
rect 298875 384371 298941 384372
rect 298323 321876 298389 321877
rect 298323 321812 298324 321876
rect 298388 321812 298389 321876
rect 298323 321811 298389 321812
rect 298326 321061 298386 321811
rect 298323 321060 298389 321061
rect 298323 320996 298324 321060
rect 298388 320996 298389 321060
rect 298323 320995 298389 320996
rect 298323 320652 298389 320653
rect 298323 320588 298324 320652
rect 298388 320588 298389 320652
rect 298323 320587 298389 320588
rect 298507 320652 298573 320653
rect 298507 320588 298508 320652
rect 298572 320588 298573 320652
rect 298507 320587 298573 320588
rect 298139 320108 298205 320109
rect 298139 320044 298140 320108
rect 298204 320044 298205 320108
rect 298139 320043 298205 320044
rect 297955 319428 298021 319429
rect 297955 319364 297956 319428
rect 298020 319364 298021 319428
rect 297955 319363 298021 319364
rect 297771 319020 297837 319021
rect 297771 318956 297772 319020
rect 297836 318956 297837 319020
rect 297771 318955 297837 318956
rect 297958 318749 298018 319363
rect 297955 318748 298021 318749
rect 297955 318684 297956 318748
rect 298020 318684 298021 318748
rect 297955 318683 298021 318684
rect 297587 310452 297653 310453
rect 297587 310388 297588 310452
rect 297652 310388 297653 310452
rect 297587 310387 297653 310388
rect 298142 293453 298202 320043
rect 298326 297397 298386 320587
rect 298510 318885 298570 320587
rect 298691 320244 298757 320245
rect 298691 320180 298692 320244
rect 298756 320180 298757 320244
rect 298691 320179 298757 320180
rect 298694 319021 298754 320179
rect 298878 320109 298938 384371
rect 299059 321604 299125 321605
rect 299059 321540 299060 321604
rect 299124 321540 299125 321604
rect 299059 321539 299125 321540
rect 299062 320109 299122 321539
rect 299246 320789 299306 393211
rect 306235 393140 306301 393141
rect 306235 393076 306236 393140
rect 306300 393076 306301 393140
rect 306235 393075 306301 393076
rect 304763 393004 304829 393005
rect 304763 392940 304764 393004
rect 304828 392940 304829 393004
rect 304763 392939 304829 392940
rect 300715 392868 300781 392869
rect 300715 392804 300716 392868
rect 300780 392804 300781 392868
rect 300715 392803 300781 392804
rect 299243 320788 299309 320789
rect 299243 320724 299244 320788
rect 299308 320724 299309 320788
rect 299243 320723 299309 320724
rect 299243 320652 299309 320653
rect 299243 320588 299244 320652
rect 299308 320588 299309 320652
rect 299243 320587 299309 320588
rect 298875 320108 298941 320109
rect 298875 320044 298876 320108
rect 298940 320044 298941 320108
rect 298875 320043 298941 320044
rect 299059 320108 299125 320109
rect 299059 320044 299060 320108
rect 299124 320044 299125 320108
rect 299059 320043 299125 320044
rect 298875 319972 298941 319973
rect 298875 319908 298876 319972
rect 298940 319908 298941 319972
rect 298875 319907 298941 319908
rect 298691 319020 298757 319021
rect 298691 318956 298692 319020
rect 298756 318956 298757 319020
rect 298691 318955 298757 318956
rect 298507 318884 298573 318885
rect 298507 318820 298508 318884
rect 298572 318820 298573 318884
rect 298507 318819 298573 318820
rect 298510 316029 298570 318819
rect 298878 316301 298938 319907
rect 299246 316437 299306 320587
rect 300347 320516 300413 320517
rect 300347 320452 300348 320516
rect 300412 320452 300413 320516
rect 300347 320451 300413 320452
rect 299427 320244 299493 320245
rect 299427 320180 299428 320244
rect 299492 320180 299493 320244
rect 299427 320179 299493 320180
rect 300163 320244 300229 320245
rect 300163 320180 300164 320244
rect 300228 320180 300229 320244
rect 300163 320179 300229 320180
rect 299430 316573 299490 320179
rect 299795 320108 299861 320109
rect 299795 320044 299796 320108
rect 299860 320044 299861 320108
rect 299795 320043 299861 320044
rect 299798 318885 299858 320043
rect 300166 319429 300226 320179
rect 300163 319428 300229 319429
rect 300163 319364 300164 319428
rect 300228 319364 300229 319428
rect 300163 319363 300229 319364
rect 300350 319021 300410 320451
rect 300531 320108 300597 320109
rect 300531 320044 300532 320108
rect 300596 320044 300597 320108
rect 300531 320043 300597 320044
rect 300534 319429 300594 320043
rect 300531 319428 300597 319429
rect 300531 319364 300532 319428
rect 300596 319364 300597 319428
rect 300531 319363 300597 319364
rect 300347 319020 300413 319021
rect 300347 318956 300348 319020
rect 300412 318956 300413 319020
rect 300347 318955 300413 318956
rect 299795 318884 299861 318885
rect 299795 318820 299796 318884
rect 299860 318820 299861 318884
rect 299795 318819 299861 318820
rect 300718 318749 300778 392803
rect 304579 392732 304645 392733
rect 304579 392668 304580 392732
rect 304644 392668 304645 392732
rect 304579 392667 304645 392668
rect 303475 392460 303541 392461
rect 303475 392396 303476 392460
rect 303540 392396 303541 392460
rect 303475 392395 303541 392396
rect 302003 385932 302069 385933
rect 302003 385868 302004 385932
rect 302068 385868 302069 385932
rect 302003 385867 302069 385868
rect 301267 321740 301333 321741
rect 301267 321676 301268 321740
rect 301332 321676 301333 321740
rect 301267 321675 301333 321676
rect 301270 320789 301330 321675
rect 301267 320788 301333 320789
rect 301267 320724 301268 320788
rect 301332 320724 301333 320788
rect 301267 320723 301333 320724
rect 301635 320516 301701 320517
rect 301635 320452 301636 320516
rect 301700 320452 301701 320516
rect 301635 320451 301701 320452
rect 300899 320108 300965 320109
rect 300899 320044 300900 320108
rect 300964 320044 300965 320108
rect 300899 320043 300965 320044
rect 300715 318748 300781 318749
rect 300715 318684 300716 318748
rect 300780 318684 300781 318748
rect 300715 318683 300781 318684
rect 300715 318476 300781 318477
rect 300715 318412 300716 318476
rect 300780 318412 300781 318476
rect 300715 318411 300781 318412
rect 300531 317796 300597 317797
rect 300531 317732 300532 317796
rect 300596 317732 300597 317796
rect 300531 317731 300597 317732
rect 299611 317524 299677 317525
rect 299611 317460 299612 317524
rect 299676 317460 299677 317524
rect 299611 317459 299677 317460
rect 299427 316572 299493 316573
rect 299427 316508 299428 316572
rect 299492 316508 299493 316572
rect 299427 316507 299493 316508
rect 299243 316436 299309 316437
rect 299243 316372 299244 316436
rect 299308 316372 299309 316436
rect 299243 316371 299309 316372
rect 298875 316300 298941 316301
rect 298875 316236 298876 316300
rect 298940 316236 298941 316300
rect 298875 316235 298941 316236
rect 298507 316028 298573 316029
rect 298507 315964 298508 316028
rect 298572 315964 298573 316028
rect 298507 315963 298573 315964
rect 299614 310317 299674 317459
rect 299611 310316 299677 310317
rect 299611 310252 299612 310316
rect 299676 310252 299677 310316
rect 299611 310251 299677 310252
rect 300534 310045 300594 317731
rect 300531 310044 300597 310045
rect 300531 309980 300532 310044
rect 300596 309980 300597 310044
rect 300531 309979 300597 309980
rect 300718 301613 300778 318411
rect 299611 301612 299677 301613
rect 299611 301548 299612 301612
rect 299676 301548 299677 301612
rect 299611 301547 299677 301548
rect 300715 301612 300781 301613
rect 300715 301548 300716 301612
rect 300780 301548 300781 301612
rect 300715 301547 300781 301548
rect 298323 297396 298389 297397
rect 298323 297332 298324 297396
rect 298388 297332 298389 297396
rect 298323 297331 298389 297332
rect 298139 293452 298205 293453
rect 298139 293388 298140 293452
rect 298204 293388 298205 293452
rect 298139 293387 298205 293388
rect 296486 219390 296914 219450
rect 296854 218925 296914 219390
rect 296851 218924 296917 218925
rect 296851 218860 296852 218924
rect 296916 218860 296917 218924
rect 296851 218859 296917 218860
rect 299614 218789 299674 301547
rect 300902 301477 300962 320043
rect 301638 319429 301698 320451
rect 302006 320109 302066 385867
rect 303478 321570 303538 392395
rect 304582 328470 304642 392667
rect 303294 321510 303538 321570
rect 304030 328410 304642 328470
rect 302739 320244 302805 320245
rect 302739 320180 302740 320244
rect 302804 320180 302805 320244
rect 302739 320179 302805 320180
rect 302003 320108 302069 320109
rect 302003 320044 302004 320108
rect 302068 320044 302069 320108
rect 302003 320043 302069 320044
rect 302555 320108 302621 320109
rect 302555 320044 302556 320108
rect 302620 320044 302621 320108
rect 302555 320043 302621 320044
rect 301635 319428 301701 319429
rect 301635 319364 301636 319428
rect 301700 319364 301701 319428
rect 301635 319363 301701 319364
rect 301267 317796 301333 317797
rect 301267 317732 301268 317796
rect 301332 317732 301333 317796
rect 301267 317731 301333 317732
rect 301083 317524 301149 317525
rect 301083 317460 301084 317524
rect 301148 317460 301149 317524
rect 301083 317459 301149 317460
rect 301086 315213 301146 317459
rect 301083 315212 301149 315213
rect 301083 315148 301084 315212
rect 301148 315148 301149 315212
rect 301083 315147 301149 315148
rect 301270 314533 301330 317731
rect 302003 317524 302069 317525
rect 302003 317460 302004 317524
rect 302068 317460 302069 317524
rect 302003 317459 302069 317460
rect 301267 314532 301333 314533
rect 301267 314468 301268 314532
rect 301332 314468 301333 314532
rect 301267 314467 301333 314468
rect 302006 306390 302066 317459
rect 302558 314125 302618 320043
rect 302742 318069 302802 320179
rect 303294 320109 303354 321510
rect 304030 320653 304090 328410
rect 304766 320789 304826 392939
rect 304947 369476 305013 369477
rect 304947 369412 304948 369476
rect 305012 369412 305013 369476
rect 304947 369411 305013 369412
rect 304950 345030 305010 369411
rect 304950 344970 305194 345030
rect 305134 325710 305194 344970
rect 305134 325650 305378 325710
rect 304763 320788 304829 320789
rect 304763 320786 304764 320788
rect 304582 320726 304764 320786
rect 304027 320652 304093 320653
rect 304027 320588 304028 320652
rect 304092 320588 304093 320652
rect 304027 320587 304093 320588
rect 303291 320108 303357 320109
rect 303291 320044 303292 320108
rect 303356 320044 303357 320108
rect 303291 320043 303357 320044
rect 303659 320108 303725 320109
rect 303659 320044 303660 320108
rect 303724 320044 303725 320108
rect 303659 320043 303725 320044
rect 302739 318068 302805 318069
rect 302739 318004 302740 318068
rect 302804 318004 302805 318068
rect 302739 318003 302805 318004
rect 303291 317796 303357 317797
rect 303291 317732 303292 317796
rect 303356 317732 303357 317796
rect 303291 317731 303357 317732
rect 302739 317524 302805 317525
rect 302739 317460 302740 317524
rect 302804 317460 302805 317524
rect 302739 317459 302805 317460
rect 302555 314124 302621 314125
rect 302555 314060 302556 314124
rect 302620 314060 302621 314124
rect 302555 314059 302621 314060
rect 302742 307733 302802 317459
rect 302739 307732 302805 307733
rect 302739 307668 302740 307732
rect 302804 307668 302805 307732
rect 302739 307667 302805 307668
rect 301454 306330 302066 306390
rect 301454 304877 301514 306330
rect 301451 304876 301517 304877
rect 301451 304812 301452 304876
rect 301516 304812 301517 304876
rect 301451 304811 301517 304812
rect 300899 301476 300965 301477
rect 300899 301412 300900 301476
rect 300964 301412 300965 301476
rect 300899 301411 300965 301412
rect 301454 219333 301514 304811
rect 303294 297941 303354 317731
rect 303475 317524 303541 317525
rect 303475 317460 303476 317524
rect 303540 317460 303541 317524
rect 303475 317459 303541 317460
rect 303291 297940 303357 297941
rect 303291 297876 303292 297940
rect 303356 297876 303357 297940
rect 303291 297875 303357 297876
rect 303294 296730 303354 297875
rect 303478 297805 303538 317459
rect 303662 317253 303722 320043
rect 303659 317252 303725 317253
rect 303659 317188 303660 317252
rect 303724 317188 303725 317252
rect 303659 317187 303725 317188
rect 303475 297804 303541 297805
rect 303475 297740 303476 297804
rect 303540 297740 303541 297804
rect 303475 297739 303541 297740
rect 302742 296670 303354 296730
rect 301451 219332 301517 219333
rect 301451 219268 301452 219332
rect 301516 219268 301517 219332
rect 301451 219267 301517 219268
rect 302742 219061 302802 296670
rect 303478 277410 303538 297739
rect 304030 293589 304090 320587
rect 304582 314261 304642 320726
rect 304763 320724 304764 320726
rect 304828 320724 304829 320788
rect 304763 320723 304829 320724
rect 304763 320244 304829 320245
rect 304763 320180 304764 320244
rect 304828 320180 304829 320244
rect 304763 320179 304829 320180
rect 304766 319021 304826 320179
rect 305131 320108 305197 320109
rect 305131 320044 305132 320108
rect 305196 320044 305197 320108
rect 305131 320043 305197 320044
rect 304763 319020 304829 319021
rect 304763 318956 304764 319020
rect 304828 318956 304829 319020
rect 304763 318955 304829 318956
rect 304763 318068 304829 318069
rect 304763 318004 304764 318068
rect 304828 318004 304829 318068
rect 304763 318003 304829 318004
rect 304579 314260 304645 314261
rect 304579 314196 304580 314260
rect 304644 314196 304645 314260
rect 304579 314195 304645 314196
rect 304766 302973 304826 318003
rect 304763 302972 304829 302973
rect 304763 302908 304764 302972
rect 304828 302908 304829 302972
rect 304763 302907 304829 302908
rect 304027 293588 304093 293589
rect 304027 293524 304028 293588
rect 304092 293524 304093 293588
rect 304027 293523 304093 293524
rect 302926 277350 303538 277410
rect 302926 219197 302986 277350
rect 305134 245309 305194 320043
rect 305318 317797 305378 325650
rect 305867 320652 305933 320653
rect 305867 320588 305868 320652
rect 305932 320588 305933 320652
rect 305867 320587 305933 320588
rect 305683 320516 305749 320517
rect 305683 320452 305684 320516
rect 305748 320452 305749 320516
rect 305683 320451 305749 320452
rect 305499 320244 305565 320245
rect 305499 320180 305500 320244
rect 305564 320180 305565 320244
rect 305499 320179 305565 320180
rect 305502 319565 305562 320179
rect 305499 319564 305565 319565
rect 305499 319500 305500 319564
rect 305564 319500 305565 319564
rect 305499 319499 305565 319500
rect 305686 319021 305746 320451
rect 305870 319565 305930 320587
rect 306238 320109 306298 393075
rect 307523 387700 307589 387701
rect 307523 387636 307524 387700
rect 307588 387636 307589 387700
rect 307523 387635 307589 387636
rect 306971 369476 307037 369477
rect 306971 369412 306972 369476
rect 307036 369412 307037 369476
rect 306971 369411 307037 369412
rect 306974 320789 307034 369411
rect 306419 320788 306485 320789
rect 306419 320724 306420 320788
rect 306484 320724 306485 320788
rect 306419 320723 306485 320724
rect 306971 320788 307037 320789
rect 306971 320724 306972 320788
rect 307036 320724 307037 320788
rect 306971 320723 307037 320724
rect 306235 320108 306301 320109
rect 306235 320044 306236 320108
rect 306300 320044 306301 320108
rect 306235 320043 306301 320044
rect 306051 319972 306117 319973
rect 306051 319908 306052 319972
rect 306116 319908 306117 319972
rect 306051 319907 306117 319908
rect 306054 319565 306114 319907
rect 305867 319564 305933 319565
rect 305867 319500 305868 319564
rect 305932 319500 305933 319564
rect 305867 319499 305933 319500
rect 306051 319564 306117 319565
rect 306051 319500 306052 319564
rect 306116 319500 306117 319564
rect 306051 319499 306117 319500
rect 305683 319020 305749 319021
rect 305683 318956 305684 319020
rect 305748 318956 305749 319020
rect 305683 318955 305749 318956
rect 305315 317796 305381 317797
rect 305315 317732 305316 317796
rect 305380 317732 305381 317796
rect 305315 317731 305381 317732
rect 305499 317524 305565 317525
rect 305499 317460 305500 317524
rect 305564 317460 305565 317524
rect 305499 317459 305565 317460
rect 305502 304197 305562 317459
rect 305499 304196 305565 304197
rect 305499 304132 305500 304196
rect 305564 304132 305565 304196
rect 305499 304131 305565 304132
rect 305131 245308 305197 245309
rect 305131 245244 305132 245308
rect 305196 245244 305197 245308
rect 305131 245243 305197 245244
rect 306422 226133 306482 320723
rect 306787 320244 306853 320245
rect 306787 320180 306788 320244
rect 306852 320180 306853 320244
rect 306787 320179 306853 320180
rect 306790 319565 306850 320179
rect 306971 320108 307037 320109
rect 306971 320044 306972 320108
rect 307036 320044 307037 320108
rect 306971 320043 307037 320044
rect 307339 320108 307405 320109
rect 307339 320044 307340 320108
rect 307404 320044 307405 320108
rect 307339 320043 307405 320044
rect 306787 319564 306853 319565
rect 306787 319500 306788 319564
rect 306852 319500 306853 319564
rect 306787 319499 306853 319500
rect 306974 318477 307034 320043
rect 307342 319429 307402 320043
rect 307339 319428 307405 319429
rect 307339 319364 307340 319428
rect 307404 319364 307405 319428
rect 307339 319363 307405 319364
rect 307526 318749 307586 387635
rect 307710 371517 307770 404227
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 310283 398852 310349 398853
rect 310283 398788 310284 398852
rect 310348 398788 310349 398852
rect 310283 398787 310349 398788
rect 308995 377500 309061 377501
rect 308995 377436 308996 377500
rect 309060 377436 309061 377500
rect 308995 377435 309061 377436
rect 307707 371516 307773 371517
rect 307707 371452 307708 371516
rect 307772 371452 307773 371516
rect 307707 371451 307773 371452
rect 307710 367709 307770 371451
rect 307707 367708 307773 367709
rect 307707 367644 307708 367708
rect 307772 367644 307773 367708
rect 307707 367643 307773 367644
rect 308259 320380 308325 320381
rect 308259 320316 308260 320380
rect 308324 320316 308325 320380
rect 308259 320315 308325 320316
rect 308075 320108 308141 320109
rect 308075 320044 308076 320108
rect 308140 320044 308141 320108
rect 308075 320043 308141 320044
rect 307891 319564 307957 319565
rect 307891 319500 307892 319564
rect 307956 319500 307957 319564
rect 307891 319499 307957 319500
rect 307894 318885 307954 319499
rect 307891 318884 307957 318885
rect 307891 318820 307892 318884
rect 307956 318820 307957 318884
rect 307891 318819 307957 318820
rect 308078 318749 308138 320043
rect 308262 319021 308322 320315
rect 308443 320244 308509 320245
rect 308443 320180 308444 320244
rect 308508 320180 308509 320244
rect 308443 320179 308509 320180
rect 308627 320244 308693 320245
rect 308627 320180 308628 320244
rect 308692 320180 308693 320244
rect 308627 320179 308693 320180
rect 308446 319565 308506 320179
rect 308443 319564 308509 319565
rect 308443 319500 308444 319564
rect 308508 319500 308509 319564
rect 308443 319499 308509 319500
rect 308630 319429 308690 320179
rect 308998 320109 309058 377435
rect 310286 320381 310346 398787
rect 321323 394228 321389 394229
rect 321323 394164 321324 394228
rect 321388 394164 321389 394228
rect 321323 394163 321389 394164
rect 311755 391780 311821 391781
rect 311755 391716 311756 391780
rect 311820 391716 311821 391780
rect 311755 391715 311821 391716
rect 311019 369476 311085 369477
rect 311019 369412 311020 369476
rect 311084 369412 311085 369476
rect 311019 369411 311085 369412
rect 311022 321570 311082 369411
rect 310838 321510 311082 321570
rect 310651 320788 310717 320789
rect 310651 320724 310652 320788
rect 310716 320724 310717 320788
rect 310651 320723 310717 320724
rect 309179 320380 309245 320381
rect 309179 320316 309180 320380
rect 309244 320316 309245 320380
rect 309179 320315 309245 320316
rect 310283 320380 310349 320381
rect 310283 320316 310284 320380
rect 310348 320316 310349 320380
rect 310283 320315 310349 320316
rect 308995 320108 309061 320109
rect 308995 320044 308996 320108
rect 309060 320044 309061 320108
rect 308995 320043 309061 320044
rect 308627 319428 308693 319429
rect 308627 319364 308628 319428
rect 308692 319364 308693 319428
rect 308627 319363 308693 319364
rect 308259 319020 308325 319021
rect 308259 318956 308260 319020
rect 308324 318956 308325 319020
rect 308259 318955 308325 318956
rect 307523 318748 307589 318749
rect 307523 318684 307524 318748
rect 307588 318684 307589 318748
rect 307523 318683 307589 318684
rect 308075 318748 308141 318749
rect 308075 318684 308076 318748
rect 308140 318684 308141 318748
rect 308075 318683 308141 318684
rect 306971 318476 307037 318477
rect 306971 318412 306972 318476
rect 307036 318412 307037 318476
rect 306971 318411 307037 318412
rect 306603 317932 306669 317933
rect 306603 317868 306604 317932
rect 306668 317868 306669 317932
rect 306603 317867 306669 317868
rect 306606 291821 306666 317867
rect 307707 317796 307773 317797
rect 307707 317732 307708 317796
rect 307772 317732 307773 317796
rect 307707 317731 307773 317732
rect 306787 317524 306853 317525
rect 306787 317460 306788 317524
rect 306852 317460 306853 317524
rect 306787 317459 306853 317460
rect 306790 314669 306850 317459
rect 306787 314668 306853 314669
rect 306787 314604 306788 314668
rect 306852 314604 306853 314668
rect 306787 314603 306853 314604
rect 307710 297669 307770 317731
rect 308259 317524 308325 317525
rect 308259 317460 308260 317524
rect 308324 317460 308325 317524
rect 308259 317459 308325 317460
rect 308262 298077 308322 317459
rect 309182 313037 309242 320315
rect 309363 320244 309429 320245
rect 309363 320180 309364 320244
rect 309428 320180 309429 320244
rect 309363 320179 309429 320180
rect 309366 319565 309426 320179
rect 309547 320108 309613 320109
rect 309547 320044 309548 320108
rect 309612 320044 309613 320108
rect 309547 320043 309613 320044
rect 310099 320108 310165 320109
rect 310099 320044 310100 320108
rect 310164 320044 310165 320108
rect 310099 320043 310165 320044
rect 309550 319565 309610 320043
rect 309363 319564 309429 319565
rect 309363 319500 309364 319564
rect 309428 319500 309429 319564
rect 309363 319499 309429 319500
rect 309547 319564 309613 319565
rect 309547 319500 309548 319564
rect 309612 319500 309613 319564
rect 309547 319499 309613 319500
rect 309731 319428 309797 319429
rect 309731 319364 309732 319428
rect 309796 319364 309797 319428
rect 309731 319363 309797 319364
rect 309734 317797 309794 319363
rect 309731 317796 309797 317797
rect 309731 317732 309732 317796
rect 309796 317732 309797 317796
rect 309731 317731 309797 317732
rect 309731 317524 309797 317525
rect 309731 317460 309732 317524
rect 309796 317460 309797 317524
rect 309731 317459 309797 317460
rect 309915 317524 309981 317525
rect 309915 317460 309916 317524
rect 309980 317460 309981 317524
rect 309915 317459 309981 317460
rect 309734 313173 309794 317459
rect 309731 313172 309797 313173
rect 309731 313108 309732 313172
rect 309796 313108 309797 313172
rect 309731 313107 309797 313108
rect 309179 313036 309245 313037
rect 309179 312972 309180 313036
rect 309244 312972 309245 313036
rect 309179 312971 309245 312972
rect 309918 311910 309978 317459
rect 310102 315757 310162 320043
rect 310283 317796 310349 317797
rect 310283 317732 310284 317796
rect 310348 317732 310349 317796
rect 310283 317731 310349 317732
rect 310099 315756 310165 315757
rect 310099 315692 310100 315756
rect 310164 315692 310165 315756
rect 310099 315691 310165 315692
rect 309734 311850 309978 311910
rect 309734 299437 309794 311850
rect 309731 299436 309797 299437
rect 309731 299372 309732 299436
rect 309796 299372 309797 299436
rect 309731 299371 309797 299372
rect 308259 298076 308325 298077
rect 308259 298012 308260 298076
rect 308324 298012 308325 298076
rect 308259 298011 308325 298012
rect 307707 297668 307773 297669
rect 307707 297604 307708 297668
rect 307772 297604 307773 297668
rect 307707 297603 307773 297604
rect 306603 291820 306669 291821
rect 306603 291756 306604 291820
rect 306668 291756 306669 291820
rect 306603 291755 306669 291756
rect 308262 277410 308322 298011
rect 309734 296730 309794 299371
rect 310286 297669 310346 317731
rect 310283 297668 310349 297669
rect 310283 297604 310284 297668
rect 310348 297604 310349 297668
rect 310283 297603 310349 297604
rect 309550 296670 309794 296730
rect 309550 277410 309610 296670
rect 310286 277410 310346 297603
rect 307710 277350 308322 277410
rect 309182 277350 309610 277410
rect 309734 277350 310346 277410
rect 306419 226132 306485 226133
rect 306419 226068 306420 226132
rect 306484 226068 306485 226132
rect 306419 226067 306485 226068
rect 307710 220557 307770 277350
rect 309182 228581 309242 277350
rect 309179 228580 309245 228581
rect 309179 228516 309180 228580
rect 309244 228516 309245 228580
rect 309179 228515 309245 228516
rect 309734 220693 309794 277350
rect 310654 238101 310714 320723
rect 310838 320109 310898 321510
rect 311758 320789 311818 391715
rect 314147 390964 314213 390965
rect 314147 390900 314148 390964
rect 314212 390900 314213 390964
rect 314147 390899 314213 390900
rect 312491 370156 312557 370157
rect 312491 370092 312492 370156
rect 312556 370092 312557 370156
rect 312491 370091 312557 370092
rect 311755 320788 311821 320789
rect 311755 320724 311756 320788
rect 311820 320724 311821 320788
rect 311755 320723 311821 320724
rect 312307 320516 312373 320517
rect 312307 320452 312308 320516
rect 312372 320452 312373 320516
rect 312307 320451 312373 320452
rect 311203 320380 311269 320381
rect 311203 320316 311204 320380
rect 311268 320316 311269 320380
rect 311203 320315 311269 320316
rect 310835 320108 310901 320109
rect 310835 320044 310836 320108
rect 310900 320044 310901 320108
rect 310835 320043 310901 320044
rect 310651 238100 310717 238101
rect 310651 238036 310652 238100
rect 310716 238036 310717 238100
rect 310651 238035 310717 238036
rect 309731 220692 309797 220693
rect 309731 220628 309732 220692
rect 309796 220628 309797 220692
rect 309731 220627 309797 220628
rect 307707 220556 307773 220557
rect 307707 220492 307708 220556
rect 307772 220492 307773 220556
rect 307707 220491 307773 220492
rect 310838 220421 310898 320043
rect 311206 319429 311266 320315
rect 312123 320108 312189 320109
rect 312123 320044 312124 320108
rect 312188 320044 312189 320108
rect 312123 320043 312189 320044
rect 311203 319428 311269 319429
rect 311203 319364 311204 319428
rect 311268 319364 311269 319428
rect 311203 319363 311269 319364
rect 312126 319021 312186 320043
rect 312310 319429 312370 320451
rect 312494 320109 312554 370091
rect 313779 369476 313845 369477
rect 313779 369412 313780 369476
rect 313844 369412 313845 369476
rect 313779 369411 313845 369412
rect 313595 320652 313661 320653
rect 313595 320588 313596 320652
rect 313660 320588 313661 320652
rect 313595 320587 313661 320588
rect 312675 320244 312741 320245
rect 312675 320180 312676 320244
rect 312740 320180 312741 320244
rect 312675 320179 312741 320180
rect 312491 320108 312557 320109
rect 312491 320044 312492 320108
rect 312556 320044 312557 320108
rect 312491 320043 312557 320044
rect 312307 319428 312373 319429
rect 312307 319364 312308 319428
rect 312372 319364 312373 319428
rect 312307 319363 312373 319364
rect 312123 319020 312189 319021
rect 312123 318956 312124 319020
rect 312188 318956 312189 319020
rect 312123 318955 312189 318956
rect 312494 314669 312554 320043
rect 312491 314668 312557 314669
rect 312491 314604 312492 314668
rect 312556 314604 312557 314668
rect 312491 314603 312557 314604
rect 312678 314533 312738 320179
rect 313598 319429 313658 320587
rect 313782 320245 313842 369411
rect 313963 320516 314029 320517
rect 313963 320452 313964 320516
rect 314028 320452 314029 320516
rect 313963 320451 314029 320452
rect 313779 320244 313845 320245
rect 313779 320180 313780 320244
rect 313844 320180 313845 320244
rect 313779 320179 313845 320180
rect 313595 319428 313661 319429
rect 313595 319364 313596 319428
rect 313660 319364 313661 319428
rect 313595 319363 313661 319364
rect 312859 317796 312925 317797
rect 312859 317732 312860 317796
rect 312924 317732 312925 317796
rect 312859 317731 312925 317732
rect 312862 314669 312922 317731
rect 313043 317524 313109 317525
rect 313043 317460 313044 317524
rect 313108 317460 313109 317524
rect 313043 317459 313109 317460
rect 313411 317524 313477 317525
rect 313411 317460 313412 317524
rect 313476 317460 313477 317524
rect 313411 317459 313477 317460
rect 312859 314668 312925 314669
rect 312859 314604 312860 314668
rect 312924 314604 312925 314668
rect 312859 314603 312925 314604
rect 312675 314532 312741 314533
rect 312675 314468 312676 314532
rect 312740 314468 312741 314532
rect 312675 314467 312741 314468
rect 313046 302021 313106 317459
rect 313414 307053 313474 317459
rect 313782 311133 313842 320179
rect 313966 319565 314026 320451
rect 314150 320109 314210 390899
rect 317275 390420 317341 390421
rect 317275 390356 317276 390420
rect 317340 390356 317341 390420
rect 317275 390355 317341 390356
rect 316723 389740 316789 389741
rect 316723 389676 316724 389740
rect 316788 389676 316789 389740
rect 316723 389675 316789 389676
rect 314699 377364 314765 377365
rect 314699 377300 314700 377364
rect 314764 377300 314765 377364
rect 314699 377299 314765 377300
rect 314331 371924 314397 371925
rect 314331 371860 314332 371924
rect 314396 371860 314397 371924
rect 314331 371859 314397 371860
rect 314147 320108 314213 320109
rect 314147 320044 314148 320108
rect 314212 320044 314213 320108
rect 314147 320043 314213 320044
rect 313963 319564 314029 319565
rect 313963 319500 313964 319564
rect 314028 319500 314029 319564
rect 313963 319499 314029 319500
rect 314150 311910 314210 320043
rect 314334 318749 314394 371859
rect 314515 321332 314581 321333
rect 314515 321268 314516 321332
rect 314580 321268 314581 321332
rect 314515 321267 314581 321268
rect 314518 320789 314578 321267
rect 314515 320788 314581 320789
rect 314515 320724 314516 320788
rect 314580 320724 314581 320788
rect 314515 320723 314581 320724
rect 314702 320109 314762 377299
rect 315619 369884 315685 369885
rect 315619 369820 315620 369884
rect 315684 369820 315685 369884
rect 315619 369819 315685 369820
rect 315435 369068 315501 369069
rect 315435 369004 315436 369068
rect 315500 369004 315501 369068
rect 315435 369003 315501 369004
rect 315438 321570 315498 369003
rect 314886 321510 315498 321570
rect 314699 320108 314765 320109
rect 314699 320044 314700 320108
rect 314764 320044 314765 320108
rect 314699 320043 314765 320044
rect 314331 318748 314397 318749
rect 314331 318684 314332 318748
rect 314396 318684 314397 318748
rect 314331 318683 314397 318684
rect 314515 317524 314581 317525
rect 314515 317460 314516 317524
rect 314580 317460 314581 317524
rect 314515 317459 314581 317460
rect 313966 311850 314210 311910
rect 313779 311132 313845 311133
rect 313779 311068 313780 311132
rect 313844 311068 313845 311132
rect 313779 311067 313845 311068
rect 313411 307052 313477 307053
rect 313411 306988 313412 307052
rect 313476 306988 313477 307052
rect 313411 306987 313477 306988
rect 313043 302020 313109 302021
rect 313043 301956 313044 302020
rect 313108 301956 313109 302020
rect 313043 301955 313109 301956
rect 313779 299436 313845 299437
rect 313779 299372 313780 299436
rect 313844 299372 313845 299436
rect 313779 299371 313845 299372
rect 310835 220420 310901 220421
rect 310835 220356 310836 220420
rect 310900 220356 310901 220420
rect 310835 220355 310901 220356
rect 313782 220149 313842 299371
rect 313966 224773 314026 311850
rect 314518 299437 314578 317459
rect 314515 299436 314581 299437
rect 314515 299372 314516 299436
rect 314580 299372 314581 299436
rect 314515 299371 314581 299372
rect 313963 224772 314029 224773
rect 313963 224708 313964 224772
rect 314028 224708 314029 224772
rect 313963 224707 314029 224708
rect 314702 220285 314762 320043
rect 314886 265573 314946 321510
rect 315438 320789 315498 321510
rect 315435 320788 315501 320789
rect 315435 320724 315436 320788
rect 315500 320724 315501 320788
rect 315435 320723 315501 320724
rect 315622 320245 315682 369819
rect 316726 321570 316786 389675
rect 316907 370564 316973 370565
rect 316907 370500 316908 370564
rect 316972 370500 316973 370564
rect 316907 370499 316973 370500
rect 316358 321510 316786 321570
rect 316358 320245 316418 321510
rect 315619 320244 315685 320245
rect 315619 320180 315620 320244
rect 315684 320180 315685 320244
rect 315619 320179 315685 320180
rect 316355 320244 316421 320245
rect 316355 320180 316356 320244
rect 316420 320180 316421 320244
rect 316355 320179 316421 320180
rect 315067 318068 315133 318069
rect 315067 318004 315068 318068
rect 315132 318004 315133 318068
rect 315067 318003 315133 318004
rect 315070 312629 315130 318003
rect 316171 317796 316237 317797
rect 316171 317732 316172 317796
rect 316236 317732 316237 317796
rect 316171 317731 316237 317732
rect 316174 312765 316234 317731
rect 316171 312764 316237 312765
rect 316171 312700 316172 312764
rect 316236 312700 316237 312764
rect 316171 312699 316237 312700
rect 315067 312628 315133 312629
rect 315067 312564 315068 312628
rect 315132 312564 315133 312628
rect 315067 312563 315133 312564
rect 314883 265572 314949 265573
rect 314883 265508 314884 265572
rect 314948 265508 314949 265572
rect 314883 265507 314949 265508
rect 316174 245173 316234 312699
rect 316358 267205 316418 320179
rect 316910 320109 316970 370499
rect 316907 320108 316973 320109
rect 316907 320044 316908 320108
rect 316972 320044 316973 320108
rect 316907 320043 316973 320044
rect 316539 318068 316605 318069
rect 316539 318004 316540 318068
rect 316604 318004 316605 318068
rect 316539 318003 316605 318004
rect 316542 286381 316602 318003
rect 316539 286380 316605 286381
rect 316539 286316 316540 286380
rect 316604 286316 316605 286380
rect 316539 286315 316605 286316
rect 316355 267204 316421 267205
rect 316355 267140 316356 267204
rect 316420 267140 316421 267204
rect 316355 267139 316421 267140
rect 316171 245172 316237 245173
rect 316171 245108 316172 245172
rect 316236 245108 316237 245172
rect 316171 245107 316237 245108
rect 316910 242317 316970 320043
rect 317278 319565 317338 390355
rect 319667 369884 319733 369885
rect 319667 369820 319668 369884
rect 319732 369820 319733 369884
rect 319667 369819 319733 369820
rect 319299 369612 319365 369613
rect 319299 369548 319300 369612
rect 319364 369548 319365 369612
rect 319299 369547 319365 369548
rect 318011 369476 318077 369477
rect 318011 369412 318012 369476
rect 318076 369412 318077 369476
rect 318011 369411 318077 369412
rect 318014 321570 318074 369411
rect 317646 321510 318074 321570
rect 317646 320109 317706 321510
rect 318931 320516 318997 320517
rect 318931 320452 318932 320516
rect 318996 320452 318997 320516
rect 318931 320451 318997 320452
rect 317643 320108 317709 320109
rect 317643 320044 317644 320108
rect 317708 320044 317709 320108
rect 317643 320043 317709 320044
rect 317275 319564 317341 319565
rect 317275 319500 317276 319564
rect 317340 319500 317341 319564
rect 317275 319499 317341 319500
rect 317459 318068 317525 318069
rect 317459 318004 317460 318068
rect 317524 318004 317525 318068
rect 317459 318003 317525 318004
rect 317462 303517 317522 318003
rect 317459 303516 317525 303517
rect 317459 303452 317460 303516
rect 317524 303452 317525 303516
rect 317459 303451 317525 303452
rect 317459 300796 317525 300797
rect 317459 300732 317460 300796
rect 317524 300732 317525 300796
rect 317459 300731 317525 300732
rect 316907 242316 316973 242317
rect 316907 242252 316908 242316
rect 316972 242252 316973 242316
rect 316907 242251 316973 242252
rect 317462 231709 317522 300731
rect 317646 294813 317706 320043
rect 318747 317932 318813 317933
rect 318747 317868 318748 317932
rect 318812 317868 318813 317932
rect 318747 317867 318813 317868
rect 318195 317796 318261 317797
rect 318195 317732 318196 317796
rect 318260 317732 318261 317796
rect 318195 317731 318261 317732
rect 318198 298893 318258 317731
rect 318379 317524 318445 317525
rect 318379 317460 318380 317524
rect 318444 317460 318445 317524
rect 318379 317459 318445 317460
rect 318382 300797 318442 317459
rect 318379 300796 318445 300797
rect 318379 300732 318380 300796
rect 318444 300732 318445 300796
rect 318379 300731 318445 300732
rect 318195 298892 318261 298893
rect 318195 298828 318196 298892
rect 318260 298828 318261 298892
rect 318195 298827 318261 298828
rect 317643 294812 317709 294813
rect 317643 294748 317644 294812
rect 317708 294748 317709 294812
rect 317643 294747 317709 294748
rect 318750 258090 318810 317867
rect 318934 264349 318994 320451
rect 319302 320109 319362 369547
rect 319670 320245 319730 369819
rect 319851 369476 319917 369477
rect 319851 369412 319852 369476
rect 319916 369412 319917 369476
rect 319851 369411 319917 369412
rect 320771 369476 320837 369477
rect 320771 369412 320772 369476
rect 320836 369412 320837 369476
rect 320771 369411 320837 369412
rect 319854 320517 319914 369411
rect 320219 321468 320285 321469
rect 320219 321404 320220 321468
rect 320284 321404 320285 321468
rect 320219 321403 320285 321404
rect 320222 320653 320282 321403
rect 320219 320652 320285 320653
rect 320219 320588 320220 320652
rect 320284 320588 320285 320652
rect 320219 320587 320285 320588
rect 319851 320516 319917 320517
rect 319851 320452 319852 320516
rect 319916 320452 319917 320516
rect 319851 320451 319917 320452
rect 319667 320244 319733 320245
rect 319667 320180 319668 320244
rect 319732 320180 319733 320244
rect 319667 320179 319733 320180
rect 319851 320244 319917 320245
rect 319851 320180 319852 320244
rect 319916 320180 319917 320244
rect 319851 320179 319917 320180
rect 320587 320244 320653 320245
rect 320587 320180 320588 320244
rect 320652 320180 320653 320244
rect 320587 320179 320653 320180
rect 319299 320108 319365 320109
rect 319299 320044 319300 320108
rect 319364 320044 319365 320108
rect 319299 320043 319365 320044
rect 319483 320108 319549 320109
rect 319483 320044 319484 320108
rect 319548 320044 319549 320108
rect 319483 320043 319549 320044
rect 319486 319021 319546 320043
rect 319483 319020 319549 319021
rect 319483 318956 319484 319020
rect 319548 318956 319549 319020
rect 319483 318955 319549 318956
rect 319670 308685 319730 320179
rect 319854 319021 319914 320179
rect 320035 320108 320101 320109
rect 320035 320044 320036 320108
rect 320100 320044 320101 320108
rect 320035 320043 320101 320044
rect 319851 319020 319917 319021
rect 319851 318956 319852 319020
rect 319916 318956 319917 319020
rect 319851 318955 319917 318956
rect 320038 318885 320098 320043
rect 320590 319565 320650 320179
rect 320587 319564 320653 319565
rect 320587 319500 320588 319564
rect 320652 319500 320653 319564
rect 320587 319499 320653 319500
rect 320035 318884 320101 318885
rect 320035 318820 320036 318884
rect 320100 318820 320101 318884
rect 320035 318819 320101 318820
rect 320774 317933 320834 369411
rect 321139 367708 321205 367709
rect 321139 367644 321140 367708
rect 321204 367644 321205 367708
rect 321139 367643 321205 367644
rect 321142 321570 321202 367643
rect 320958 321510 321202 321570
rect 320958 320109 321018 321510
rect 321326 320109 321386 394163
rect 323163 371380 323229 371381
rect 323163 371316 323164 371380
rect 323228 371316 323229 371380
rect 323163 371315 323229 371316
rect 322059 369476 322125 369477
rect 322059 369412 322060 369476
rect 322124 369412 322125 369476
rect 322059 369411 322125 369412
rect 321691 322012 321757 322013
rect 321691 321948 321692 322012
rect 321756 321948 321757 322012
rect 321691 321947 321757 321948
rect 321507 321740 321573 321741
rect 321507 321676 321508 321740
rect 321572 321676 321573 321740
rect 321507 321675 321573 321676
rect 321510 320925 321570 321675
rect 321507 320924 321573 320925
rect 321507 320860 321508 320924
rect 321572 320860 321573 320924
rect 321507 320859 321573 320860
rect 321694 320789 321754 321947
rect 322062 320789 322122 369411
rect 323166 366349 323226 371315
rect 323163 366348 323229 366349
rect 323163 366284 323164 366348
rect 323228 366284 323229 366348
rect 323163 366283 323229 366284
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325371 345676 325437 345677
rect 325371 345612 325372 345676
rect 325436 345612 325437 345676
rect 325371 345611 325437 345612
rect 324267 342956 324333 342957
rect 324267 342892 324268 342956
rect 324332 342892 324333 342956
rect 324267 342891 324333 342892
rect 323347 325820 323413 325821
rect 323347 325756 323348 325820
rect 323412 325756 323413 325820
rect 323347 325755 323413 325756
rect 321691 320788 321757 320789
rect 321691 320724 321692 320788
rect 321756 320724 321757 320788
rect 321691 320723 321757 320724
rect 322059 320788 322125 320789
rect 322059 320724 322060 320788
rect 322124 320724 322125 320788
rect 322059 320723 322125 320724
rect 320955 320108 321021 320109
rect 320955 320044 320956 320108
rect 321020 320044 321021 320108
rect 320955 320043 321021 320044
rect 321323 320108 321389 320109
rect 321323 320044 321324 320108
rect 321388 320044 321389 320108
rect 321323 320043 321389 320044
rect 320771 317932 320837 317933
rect 320771 317868 320772 317932
rect 320836 317868 320837 317932
rect 320771 317867 320837 317868
rect 320587 317524 320653 317525
rect 320587 317460 320588 317524
rect 320652 317460 320653 317524
rect 320587 317459 320653 317460
rect 319667 308684 319733 308685
rect 319667 308620 319668 308684
rect 319732 308620 319733 308684
rect 319667 308619 319733 308620
rect 320590 305013 320650 317459
rect 320774 313173 320834 317867
rect 320771 313172 320837 313173
rect 320771 313108 320772 313172
rect 320836 313108 320837 313172
rect 320771 313107 320837 313108
rect 320587 305012 320653 305013
rect 320587 304948 320588 305012
rect 320652 304948 320653 305012
rect 320587 304947 320653 304948
rect 318931 264348 318997 264349
rect 318931 264284 318932 264348
rect 318996 264284 318997 264348
rect 318931 264283 318997 264284
rect 318750 258030 318994 258090
rect 317459 231708 317525 231709
rect 317459 231644 317460 231708
rect 317524 231644 317525 231708
rect 317459 231643 317525 231644
rect 314699 220284 314765 220285
rect 314699 220220 314700 220284
rect 314764 220220 314765 220284
rect 314699 220219 314765 220220
rect 313779 220148 313845 220149
rect 313779 220084 313780 220148
rect 313844 220084 313845 220148
rect 313779 220083 313845 220084
rect 302923 219196 302989 219197
rect 302923 219132 302924 219196
rect 302988 219132 302989 219196
rect 302923 219131 302989 219132
rect 302739 219060 302805 219061
rect 302739 218996 302740 219060
rect 302804 218996 302805 219060
rect 302739 218995 302805 218996
rect 299611 218788 299677 218789
rect 299611 218724 299612 218788
rect 299676 218724 299677 218788
rect 299611 218723 299677 218724
rect 318934 216613 318994 258030
rect 320958 243677 321018 320043
rect 321326 318341 321386 320043
rect 321323 318340 321389 318341
rect 321323 318276 321324 318340
rect 321388 318276 321389 318340
rect 321323 318275 321389 318276
rect 322062 311910 322122 320723
rect 323163 320516 323229 320517
rect 323163 320452 323164 320516
rect 323228 320452 323229 320516
rect 323163 320451 323229 320452
rect 322979 320380 323045 320381
rect 322979 320316 322980 320380
rect 323044 320316 323045 320380
rect 322979 320315 323045 320316
rect 322795 320108 322861 320109
rect 322795 320044 322796 320108
rect 322860 320044 322861 320108
rect 322795 320043 322861 320044
rect 322798 317933 322858 320043
rect 322795 317932 322861 317933
rect 322795 317868 322796 317932
rect 322860 317868 322861 317932
rect 322795 317867 322861 317868
rect 322795 317660 322861 317661
rect 322795 317596 322796 317660
rect 322860 317596 322861 317660
rect 322795 317595 322861 317596
rect 322611 317524 322677 317525
rect 322611 317460 322612 317524
rect 322676 317460 322677 317524
rect 322611 317459 322677 317460
rect 321326 311850 322122 311910
rect 321326 302250 321386 311850
rect 322614 311133 322674 317459
rect 322611 311132 322677 311133
rect 322611 311068 322612 311132
rect 322676 311068 322677 311132
rect 322611 311067 322677 311068
rect 322798 307597 322858 317595
rect 322795 307596 322861 307597
rect 322795 307532 322796 307596
rect 322860 307532 322861 307596
rect 322795 307531 322861 307532
rect 321326 302190 321570 302250
rect 320955 243676 321021 243677
rect 320955 243612 320956 243676
rect 321020 243612 321021 243676
rect 320955 243611 321021 243612
rect 321510 223141 321570 302190
rect 322982 243813 323042 320315
rect 323166 313173 323226 320451
rect 323350 318613 323410 325755
rect 323531 325004 323597 325005
rect 323531 324940 323532 325004
rect 323596 324940 323597 325004
rect 323531 324939 323597 324940
rect 323534 320381 323594 324939
rect 323715 322964 323781 322965
rect 323715 322900 323716 322964
rect 323780 322900 323781 322964
rect 323715 322899 323781 322900
rect 323531 320380 323597 320381
rect 323531 320316 323532 320380
rect 323596 320316 323597 320380
rect 323531 320315 323597 320316
rect 323531 320108 323597 320109
rect 323531 320044 323532 320108
rect 323596 320044 323597 320108
rect 323531 320043 323597 320044
rect 323534 319565 323594 320043
rect 323718 319565 323778 322899
rect 324083 321876 324149 321877
rect 324083 321812 324084 321876
rect 324148 321812 324149 321876
rect 324083 321811 324149 321812
rect 324086 320789 324146 321811
rect 324083 320788 324149 320789
rect 324083 320724 324084 320788
rect 324148 320724 324149 320788
rect 324083 320723 324149 320724
rect 324270 320381 324330 342891
rect 325187 322012 325253 322013
rect 325187 321948 325188 322012
rect 325252 321948 325253 322012
rect 325187 321947 325253 321948
rect 325190 320789 325250 321947
rect 325187 320788 325253 320789
rect 325187 320724 325188 320788
rect 325252 320724 325253 320788
rect 325187 320723 325253 320724
rect 324819 320652 324885 320653
rect 324819 320588 324820 320652
rect 324884 320588 324885 320652
rect 324819 320587 324885 320588
rect 324635 320516 324701 320517
rect 324635 320452 324636 320516
rect 324700 320452 324701 320516
rect 324635 320451 324701 320452
rect 324267 320380 324333 320381
rect 324267 320316 324268 320380
rect 324332 320316 324333 320380
rect 324267 320315 324333 320316
rect 324451 320108 324517 320109
rect 324451 320044 324452 320108
rect 324516 320044 324517 320108
rect 324451 320043 324517 320044
rect 323531 319564 323597 319565
rect 323531 319500 323532 319564
rect 323596 319500 323597 319564
rect 323531 319499 323597 319500
rect 323715 319564 323781 319565
rect 323715 319500 323716 319564
rect 323780 319500 323781 319564
rect 323715 319499 323781 319500
rect 324454 319021 324514 320043
rect 324451 319020 324517 319021
rect 324451 318956 324452 319020
rect 324516 318956 324517 319020
rect 324451 318955 324517 318956
rect 324638 318885 324698 320451
rect 324822 318885 324882 320587
rect 325187 320380 325253 320381
rect 325187 320316 325188 320380
rect 325252 320316 325253 320380
rect 325187 320315 325253 320316
rect 325003 319972 325069 319973
rect 325003 319908 325004 319972
rect 325068 319908 325069 319972
rect 325003 319907 325069 319908
rect 325006 319021 325066 319907
rect 325003 319020 325069 319021
rect 325003 318956 325004 319020
rect 325068 318956 325069 319020
rect 325003 318955 325069 318956
rect 325190 318885 325250 320315
rect 325374 320109 325434 345611
rect 325794 327454 326414 362898
rect 329514 705798 330134 705830
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 343955 451620 344021 451621
rect 343955 451556 343956 451620
rect 344020 451556 344021 451620
rect 343955 451555 344021 451556
rect 343771 449444 343837 449445
rect 343771 449380 343772 449444
rect 343836 449380 343837 449444
rect 343771 449379 343837 449380
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 343774 408510 343834 449379
rect 343958 443597 344018 451555
rect 355179 451348 355245 451349
rect 355179 451284 355180 451348
rect 355244 451284 355245 451348
rect 355179 451283 355245 451284
rect 345795 449444 345861 449445
rect 345795 449380 345796 449444
rect 345860 449380 345861 449444
rect 345795 449379 345861 449380
rect 347451 449444 347517 449445
rect 347451 449380 347452 449444
rect 347516 449380 347517 449444
rect 347451 449379 347517 449380
rect 345798 447813 345858 449379
rect 347454 447949 347514 449379
rect 347635 449308 347701 449309
rect 347635 449244 347636 449308
rect 347700 449244 347701 449308
rect 347635 449243 347701 449244
rect 347638 448629 347698 449243
rect 347635 448628 347701 448629
rect 347635 448564 347636 448628
rect 347700 448564 347701 448628
rect 347635 448563 347701 448564
rect 347451 447948 347517 447949
rect 347451 447884 347452 447948
rect 347516 447884 347517 447948
rect 347451 447883 347517 447884
rect 345795 447812 345861 447813
rect 345795 447748 345796 447812
rect 345860 447748 345861 447812
rect 345795 447747 345861 447748
rect 343955 443596 344021 443597
rect 343955 443532 343956 443596
rect 344020 443532 344021 443596
rect 343955 443531 344021 443532
rect 343774 408450 344018 408510
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 343958 402253 344018 408450
rect 343955 402252 344021 402253
rect 343955 402188 343956 402252
rect 344020 402188 344021 402252
rect 343955 402187 344021 402188
rect 343035 402116 343101 402117
rect 343035 402052 343036 402116
rect 343100 402052 343101 402116
rect 343035 402051 343101 402052
rect 343038 399941 343098 402051
rect 343771 400484 343837 400485
rect 343771 400420 343772 400484
rect 343836 400420 343837 400484
rect 343771 400419 343837 400420
rect 343774 399941 343834 400419
rect 343035 399940 343101 399941
rect 343035 399876 343036 399940
rect 343100 399876 343101 399940
rect 343035 399875 343101 399876
rect 343771 399940 343837 399941
rect 343771 399876 343772 399940
rect 343836 399876 343837 399940
rect 343771 399875 343837 399876
rect 342299 399804 342365 399805
rect 342299 399740 342300 399804
rect 342364 399740 342365 399804
rect 342299 399739 342365 399740
rect 343219 399804 343285 399805
rect 343219 399740 343220 399804
rect 343284 399740 343285 399804
rect 343219 399739 343285 399740
rect 342302 395589 342362 399739
rect 343222 398173 343282 399739
rect 343958 399397 344018 402187
rect 347635 401708 347701 401709
rect 347635 401644 347636 401708
rect 347700 401644 347701 401708
rect 347635 401643 347701 401644
rect 345795 400348 345861 400349
rect 345795 400284 345796 400348
rect 345860 400284 345861 400348
rect 345795 400283 345861 400284
rect 345798 399941 345858 400283
rect 347638 399941 347698 401643
rect 355182 401301 355242 451283
rect 360331 449988 360397 449989
rect 360331 449924 360332 449988
rect 360396 449924 360397 449988
rect 360331 449923 360397 449924
rect 360147 447540 360213 447541
rect 360147 447476 360148 447540
rect 360212 447476 360213 447540
rect 360147 447475 360213 447476
rect 360150 401981 360210 447475
rect 360334 414030 360394 449923
rect 360515 449852 360581 449853
rect 360515 449788 360516 449852
rect 360580 449788 360581 449852
rect 360515 449787 360581 449788
rect 360518 447541 360578 449787
rect 360515 447540 360581 447541
rect 360515 447476 360516 447540
rect 360580 447476 360581 447540
rect 360515 447475 360581 447476
rect 361794 435454 362414 470898
rect 365514 705798 366134 705830
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 362907 451348 362973 451349
rect 362907 451284 362908 451348
rect 362972 451284 362973 451348
rect 362907 451283 362973 451284
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 360334 413970 360578 414030
rect 360518 412650 360578 413970
rect 360518 412590 360946 412650
rect 360886 411270 360946 412590
rect 360334 411210 360946 411270
rect 360147 401980 360213 401981
rect 360147 401916 360148 401980
rect 360212 401916 360213 401980
rect 360147 401915 360213 401916
rect 355179 401300 355245 401301
rect 355179 401236 355180 401300
rect 355244 401236 355245 401300
rect 355179 401235 355245 401236
rect 360334 401029 360394 411210
rect 360515 401980 360581 401981
rect 360515 401916 360516 401980
rect 360580 401916 360581 401980
rect 360515 401915 360581 401916
rect 360331 401028 360397 401029
rect 360331 400964 360332 401028
rect 360396 400964 360397 401028
rect 360331 400963 360397 400964
rect 352419 400756 352485 400757
rect 352419 400692 352420 400756
rect 352484 400692 352485 400756
rect 352419 400691 352485 400692
rect 344691 399940 344757 399941
rect 344691 399876 344692 399940
rect 344756 399876 344757 399940
rect 344691 399875 344757 399876
rect 345059 399940 345125 399941
rect 345059 399876 345060 399940
rect 345124 399876 345125 399940
rect 345059 399875 345125 399876
rect 345427 399940 345493 399941
rect 345427 399876 345428 399940
rect 345492 399876 345493 399940
rect 345427 399875 345493 399876
rect 345795 399940 345861 399941
rect 345795 399876 345796 399940
rect 345860 399876 345861 399940
rect 345795 399875 345861 399876
rect 347267 399940 347333 399941
rect 347267 399876 347268 399940
rect 347332 399876 347333 399940
rect 347267 399875 347333 399876
rect 347635 399940 347701 399941
rect 347635 399876 347636 399940
rect 347700 399876 347701 399940
rect 347635 399875 347701 399876
rect 348003 399940 348069 399941
rect 348003 399876 348004 399940
rect 348068 399876 348069 399940
rect 348003 399875 348069 399876
rect 348371 399940 348437 399941
rect 348371 399876 348372 399940
rect 348436 399876 348437 399940
rect 348371 399875 348437 399876
rect 348555 399940 348621 399941
rect 348555 399876 348556 399940
rect 348620 399876 348621 399940
rect 348555 399875 348621 399876
rect 350395 399940 350461 399941
rect 350395 399876 350396 399940
rect 350460 399876 350461 399940
rect 350395 399875 350461 399876
rect 350579 399940 350645 399941
rect 350579 399876 350580 399940
rect 350644 399876 350645 399940
rect 350579 399875 350645 399876
rect 352235 399940 352301 399941
rect 352235 399876 352236 399940
rect 352300 399876 352301 399940
rect 352235 399875 352301 399876
rect 343955 399396 344021 399397
rect 343955 399332 343956 399396
rect 344020 399332 344021 399396
rect 343955 399331 344021 399332
rect 343219 398172 343285 398173
rect 343219 398108 343220 398172
rect 343284 398108 343285 398172
rect 343219 398107 343285 398108
rect 342299 395588 342365 395589
rect 342299 395524 342300 395588
rect 342364 395524 342365 395588
rect 342299 395523 342365 395524
rect 344694 393413 344754 399875
rect 344691 393412 344757 393413
rect 344691 393348 344692 393412
rect 344756 393348 344757 393412
rect 344691 393347 344757 393348
rect 341011 392052 341077 392053
rect 341011 391988 341012 392052
rect 341076 391988 341077 392052
rect 341011 391987 341077 391988
rect 341014 389190 341074 391987
rect 345062 390010 345122 399875
rect 345243 399804 345309 399805
rect 345243 399740 345244 399804
rect 345308 399740 345309 399804
rect 345243 399739 345309 399740
rect 340830 389130 341074 389190
rect 344878 389950 345122 390010
rect 331811 370020 331877 370021
rect 331811 369956 331812 370020
rect 331876 369956 331877 370020
rect 331811 369955 331877 369956
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 326843 328540 326909 328541
rect 326843 328476 326844 328540
rect 326908 328476 326909 328540
rect 326843 328475 326909 328476
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325555 320924 325621 320925
rect 325555 320860 325556 320924
rect 325620 320860 325621 320924
rect 325555 320859 325621 320860
rect 325371 320108 325437 320109
rect 325371 320044 325372 320108
rect 325436 320044 325437 320108
rect 325371 320043 325437 320044
rect 325371 319972 325437 319973
rect 325371 319908 325372 319972
rect 325436 319908 325437 319972
rect 325371 319907 325437 319908
rect 325374 319565 325434 319907
rect 325371 319564 325437 319565
rect 325371 319500 325372 319564
rect 325436 319500 325437 319564
rect 325371 319499 325437 319500
rect 324635 318884 324701 318885
rect 324635 318820 324636 318884
rect 324700 318820 324701 318884
rect 324635 318819 324701 318820
rect 324819 318884 324885 318885
rect 324819 318820 324820 318884
rect 324884 318820 324885 318884
rect 324819 318819 324885 318820
rect 325187 318884 325253 318885
rect 325187 318820 325188 318884
rect 325252 318820 325253 318884
rect 325187 318819 325253 318820
rect 325558 318749 325618 320859
rect 325555 318748 325621 318749
rect 325555 318684 325556 318748
rect 325620 318684 325621 318748
rect 325555 318683 325621 318684
rect 323347 318612 323413 318613
rect 323347 318548 323348 318612
rect 323412 318548 323413 318612
rect 323347 318547 323413 318548
rect 324451 317932 324517 317933
rect 324451 317868 324452 317932
rect 324516 317868 324517 317932
rect 324451 317867 324517 317868
rect 323163 313172 323229 313173
rect 323163 313108 323164 313172
rect 323228 313108 323229 313172
rect 323163 313107 323229 313108
rect 322979 243812 323045 243813
rect 322979 243748 322980 243812
rect 323044 243748 323045 243812
rect 322979 243747 323045 243748
rect 324454 243541 324514 317867
rect 325555 317796 325621 317797
rect 325555 317732 325556 317796
rect 325620 317732 325621 317796
rect 325555 317731 325621 317732
rect 325558 316845 325618 317731
rect 325555 316844 325621 316845
rect 325555 316780 325556 316844
rect 325620 316780 325621 316844
rect 325555 316779 325621 316780
rect 325794 291454 326414 326898
rect 326659 321604 326725 321605
rect 326659 321540 326660 321604
rect 326724 321540 326725 321604
rect 326659 321539 326725 321540
rect 326662 320789 326722 321539
rect 326659 320788 326725 320789
rect 326659 320724 326660 320788
rect 326724 320724 326725 320788
rect 326659 320723 326725 320724
rect 326846 320517 326906 328475
rect 327579 326364 327645 326365
rect 327579 326300 327580 326364
rect 327644 326300 327645 326364
rect 327579 326299 327645 326300
rect 327395 320788 327461 320789
rect 327395 320724 327396 320788
rect 327460 320724 327461 320788
rect 327395 320723 327461 320724
rect 326843 320516 326909 320517
rect 326843 320452 326844 320516
rect 326908 320452 326909 320516
rect 326843 320451 326909 320452
rect 327211 320108 327277 320109
rect 327211 320044 327212 320108
rect 327276 320044 327277 320108
rect 327211 320043 327277 320044
rect 326659 319972 326725 319973
rect 326659 319908 326660 319972
rect 326724 319908 326725 319972
rect 326659 319907 326725 319908
rect 326662 319565 326722 319907
rect 327214 319565 327274 320043
rect 327398 319565 327458 320723
rect 327582 320653 327642 326299
rect 327763 324460 327829 324461
rect 327763 324396 327764 324460
rect 327828 324396 327829 324460
rect 327763 324395 327829 324396
rect 327579 320652 327645 320653
rect 327579 320588 327580 320652
rect 327644 320588 327645 320652
rect 327579 320587 327645 320588
rect 327582 319973 327642 320587
rect 327766 320517 327826 324395
rect 327763 320516 327829 320517
rect 327763 320452 327764 320516
rect 327828 320452 327829 320516
rect 327763 320451 327829 320452
rect 327579 319972 327645 319973
rect 327579 319908 327580 319972
rect 327644 319908 327645 319972
rect 327579 319907 327645 319908
rect 326659 319564 326725 319565
rect 326659 319500 326660 319564
rect 326724 319500 326725 319564
rect 326659 319499 326725 319500
rect 327211 319564 327277 319565
rect 327211 319500 327212 319564
rect 327276 319500 327277 319564
rect 327211 319499 327277 319500
rect 327395 319564 327461 319565
rect 327395 319500 327396 319564
rect 327460 319500 327461 319564
rect 327395 319499 327461 319500
rect 328499 318884 328565 318885
rect 328499 318820 328500 318884
rect 328564 318820 328565 318884
rect 328499 318819 328565 318820
rect 326659 318068 326725 318069
rect 326659 318004 326660 318068
rect 326724 318004 326725 318068
rect 326659 318003 326725 318004
rect 326662 316981 326722 318003
rect 327579 317932 327645 317933
rect 327579 317868 327580 317932
rect 327644 317868 327645 317932
rect 327579 317867 327645 317868
rect 327027 317796 327093 317797
rect 327027 317732 327028 317796
rect 327092 317732 327093 317796
rect 327027 317731 327093 317732
rect 326843 317524 326909 317525
rect 326843 317460 326844 317524
rect 326908 317460 326909 317524
rect 326843 317459 326909 317460
rect 326659 316980 326725 316981
rect 326659 316916 326660 316980
rect 326724 316916 326725 316980
rect 326659 316915 326725 316916
rect 326846 310453 326906 317459
rect 326843 310452 326909 310453
rect 326843 310388 326844 310452
rect 326908 310388 326909 310452
rect 326843 310387 326909 310388
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 324451 243540 324517 243541
rect 324451 243476 324452 243540
rect 324516 243476 324517 243540
rect 324451 243475 324517 243476
rect 321507 223140 321573 223141
rect 321507 223076 321508 223140
rect 321572 223076 321573 223140
rect 321507 223075 321573 223076
rect 325794 219454 326414 254898
rect 327030 249253 327090 317731
rect 327582 306509 327642 317867
rect 327579 306508 327645 306509
rect 327579 306444 327580 306508
rect 327644 306444 327645 306508
rect 327579 306443 327645 306444
rect 327027 249252 327093 249253
rect 327027 249188 327028 249252
rect 327092 249188 327093 249252
rect 327027 249187 327093 249188
rect 327582 231301 327642 306443
rect 328502 240821 328562 318819
rect 328683 317932 328749 317933
rect 328683 317868 328684 317932
rect 328748 317868 328749 317932
rect 328683 317867 328749 317868
rect 328686 309501 328746 317867
rect 328683 309500 328749 309501
rect 328683 309436 328684 309500
rect 328748 309436 328749 309500
rect 328683 309435 328749 309436
rect 329514 295174 330134 330618
rect 330339 325140 330405 325141
rect 330339 325076 330340 325140
rect 330404 325076 330405 325140
rect 330339 325075 330405 325076
rect 330342 324461 330402 325075
rect 330339 324460 330405 324461
rect 330339 324396 330340 324460
rect 330404 324396 330405 324460
rect 330339 324395 330405 324396
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 328499 240820 328565 240821
rect 328499 240756 328500 240820
rect 328564 240756 328565 240820
rect 328499 240755 328565 240756
rect 327579 231300 327645 231301
rect 327579 231236 327580 231300
rect 327644 231236 327645 231300
rect 327579 231235 327645 231236
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 318931 216612 318997 216613
rect 318931 216548 318932 216612
rect 318996 216548 318997 216612
rect 318931 216547 318997 216548
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -1894 294134 -1862
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 223174 330134 258618
rect 330342 228853 330402 324395
rect 330707 321876 330773 321877
rect 330707 321812 330708 321876
rect 330772 321812 330773 321876
rect 330707 321811 330773 321812
rect 330523 321604 330589 321605
rect 330523 321540 330524 321604
rect 330588 321540 330589 321604
rect 330523 321539 330589 321540
rect 330339 228852 330405 228853
rect 330339 228788 330340 228852
rect 330404 228788 330405 228852
rect 330339 228787 330405 228788
rect 330526 227493 330586 321539
rect 330710 300253 330770 321811
rect 330707 300252 330773 300253
rect 330707 300188 330708 300252
rect 330772 300188 330773 300252
rect 330707 300187 330773 300188
rect 330523 227492 330589 227493
rect 330523 227428 330524 227492
rect 330588 227428 330589 227492
rect 330523 227427 330589 227428
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 331814 111893 331874 369955
rect 335859 369884 335925 369885
rect 335859 369820 335860 369884
rect 335924 369820 335925 369884
rect 335859 369819 335925 369820
rect 331811 111892 331877 111893
rect 331811 111828 331812 111892
rect 331876 111828 331877 111892
rect 331811 111827 331877 111828
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 335862 59397 335922 369819
rect 338251 329084 338317 329085
rect 338251 329020 338252 329084
rect 338316 329020 338317 329084
rect 338251 329019 338317 329020
rect 338254 228989 338314 329019
rect 340830 316709 340890 389130
rect 344878 388517 344938 389950
rect 345059 389876 345125 389877
rect 345059 389812 345060 389876
rect 345124 389812 345125 389876
rect 345059 389811 345125 389812
rect 344875 388516 344941 388517
rect 344875 388452 344876 388516
rect 344940 388452 344941 388516
rect 344875 388451 344941 388452
rect 340827 316708 340893 316709
rect 340827 316644 340828 316708
rect 340892 316644 340893 316708
rect 340827 316643 340893 316644
rect 345062 307053 345122 389811
rect 345246 388381 345306 399739
rect 345430 394773 345490 399875
rect 346347 399804 346413 399805
rect 346347 399740 346348 399804
rect 346412 399740 346413 399804
rect 346347 399739 346413 399740
rect 345427 394772 345493 394773
rect 345427 394708 345428 394772
rect 345492 394708 345493 394772
rect 345427 394707 345493 394708
rect 345243 388380 345309 388381
rect 345243 388316 345244 388380
rect 345308 388316 345309 388380
rect 345243 388315 345309 388316
rect 345059 307052 345125 307053
rect 345059 306988 345060 307052
rect 345124 306988 345125 307052
rect 345059 306987 345125 306988
rect 346350 296989 346410 399739
rect 347270 387021 347330 399875
rect 348006 398173 348066 399875
rect 348003 398172 348069 398173
rect 348003 398108 348004 398172
rect 348068 398108 348069 398172
rect 348003 398107 348069 398108
rect 347819 393412 347885 393413
rect 347819 393348 347820 393412
rect 347884 393348 347885 393412
rect 347819 393347 347885 393348
rect 347267 387020 347333 387021
rect 347267 386956 347268 387020
rect 347332 386956 347333 387020
rect 347267 386955 347333 386956
rect 346347 296988 346413 296989
rect 346347 296924 346348 296988
rect 346412 296924 346413 296988
rect 346347 296923 346413 296924
rect 347822 294677 347882 393347
rect 348374 388789 348434 399875
rect 348371 388788 348437 388789
rect 348371 388724 348372 388788
rect 348436 388724 348437 388788
rect 348371 388723 348437 388724
rect 348558 388653 348618 399875
rect 350027 399804 350093 399805
rect 350027 399740 350028 399804
rect 350092 399740 350093 399804
rect 350027 399739 350093 399740
rect 349107 399260 349173 399261
rect 349107 399196 349108 399260
rect 349172 399196 349173 399260
rect 349107 399195 349173 399196
rect 348555 388652 348621 388653
rect 348555 388588 348556 388652
rect 348620 388588 348621 388652
rect 348555 388587 348621 388588
rect 349110 298757 349170 399195
rect 350030 393549 350090 399739
rect 350398 397493 350458 399875
rect 350395 397492 350461 397493
rect 350395 397428 350396 397492
rect 350460 397428 350461 397492
rect 350395 397427 350461 397428
rect 350027 393548 350093 393549
rect 350027 393484 350028 393548
rect 350092 393484 350093 393548
rect 350027 393483 350093 393484
rect 349291 393412 349357 393413
rect 349291 393348 349292 393412
rect 349356 393348 349357 393412
rect 349291 393347 349357 393348
rect 349294 299165 349354 393347
rect 350582 299301 350642 399875
rect 351683 399804 351749 399805
rect 351683 399740 351684 399804
rect 351748 399740 351749 399804
rect 351683 399739 351749 399740
rect 350763 398580 350829 398581
rect 350763 398516 350764 398580
rect 350828 398516 350829 398580
rect 350763 398515 350829 398516
rect 350766 321333 350826 398515
rect 351686 393330 351746 399739
rect 351686 393270 352114 393330
rect 350763 321332 350829 321333
rect 350763 321268 350764 321332
rect 350828 321268 350829 321332
rect 350763 321267 350829 321268
rect 350579 299300 350645 299301
rect 350579 299236 350580 299300
rect 350644 299236 350645 299300
rect 350579 299235 350645 299236
rect 349291 299164 349357 299165
rect 349291 299100 349292 299164
rect 349356 299100 349357 299164
rect 349291 299099 349357 299100
rect 349107 298756 349173 298757
rect 349107 298692 349108 298756
rect 349172 298692 349173 298756
rect 349107 298691 349173 298692
rect 352054 295085 352114 393270
rect 352238 392597 352298 399875
rect 352422 399805 352482 400691
rect 355363 400620 355429 400621
rect 355363 400556 355364 400620
rect 355428 400556 355429 400620
rect 355363 400555 355429 400556
rect 354075 400348 354141 400349
rect 354075 400284 354076 400348
rect 354140 400284 354141 400348
rect 354075 400283 354141 400284
rect 353707 399940 353773 399941
rect 353707 399876 353708 399940
rect 353772 399876 353773 399940
rect 353707 399875 353773 399876
rect 352419 399804 352485 399805
rect 352419 399740 352420 399804
rect 352484 399740 352485 399804
rect 352419 399739 352485 399740
rect 353155 399804 353221 399805
rect 353155 399740 353156 399804
rect 353220 399740 353221 399804
rect 353155 399739 353221 399740
rect 352419 398308 352485 398309
rect 352419 398244 352420 398308
rect 352484 398244 352485 398308
rect 352419 398243 352485 398244
rect 352235 392596 352301 392597
rect 352235 392532 352236 392596
rect 352300 392532 352301 392596
rect 352235 392531 352301 392532
rect 352422 315485 352482 398243
rect 353158 397493 353218 399739
rect 353339 399260 353405 399261
rect 353339 399196 353340 399260
rect 353404 399196 353405 399260
rect 353339 399195 353405 399196
rect 353155 397492 353221 397493
rect 353155 397428 353156 397492
rect 353220 397428 353221 397492
rect 353155 397427 353221 397428
rect 353342 377909 353402 399195
rect 353710 391645 353770 399875
rect 354078 399805 354138 400283
rect 354262 400150 354690 400210
rect 354075 399804 354141 399805
rect 354075 399740 354076 399804
rect 354140 399740 354141 399804
rect 354075 399739 354141 399740
rect 354262 396269 354322 400150
rect 354630 400077 354690 400150
rect 354443 400076 354509 400077
rect 354443 400012 354444 400076
rect 354508 400012 354509 400076
rect 354443 400011 354509 400012
rect 354627 400076 354693 400077
rect 354627 400012 354628 400076
rect 354692 400012 354693 400076
rect 354627 400011 354693 400012
rect 355179 400076 355245 400077
rect 355179 400012 355180 400076
rect 355244 400012 355245 400076
rect 355179 400011 355245 400012
rect 354259 396268 354325 396269
rect 354259 396204 354260 396268
rect 354324 396204 354325 396268
rect 354259 396203 354325 396204
rect 353707 391644 353773 391645
rect 353707 391580 353708 391644
rect 353772 391580 353773 391644
rect 353707 391579 353773 391580
rect 353339 377908 353405 377909
rect 353339 377844 353340 377908
rect 353404 377844 353405 377908
rect 353339 377843 353405 377844
rect 352419 315484 352485 315485
rect 352419 315420 352420 315484
rect 352484 315420 352485 315484
rect 352419 315419 352485 315420
rect 354446 295221 354506 400011
rect 354627 399940 354693 399941
rect 354627 399876 354628 399940
rect 354692 399876 354693 399940
rect 354627 399875 354693 399876
rect 354630 395317 354690 399875
rect 355182 399669 355242 400011
rect 355366 399669 355426 400555
rect 355547 400212 355613 400213
rect 355547 400148 355548 400212
rect 355612 400148 355613 400212
rect 355547 400147 355613 400148
rect 357387 400212 357453 400213
rect 357387 400148 357388 400212
rect 357452 400148 357453 400212
rect 357387 400147 357453 400148
rect 355550 399941 355610 400147
rect 355547 399940 355613 399941
rect 355547 399876 355548 399940
rect 355612 399876 355613 399940
rect 355547 399875 355613 399876
rect 355179 399668 355245 399669
rect 355179 399604 355180 399668
rect 355244 399604 355245 399668
rect 355179 399603 355245 399604
rect 355363 399668 355429 399669
rect 355363 399604 355364 399668
rect 355428 399604 355429 399668
rect 355363 399603 355429 399604
rect 355547 399668 355613 399669
rect 355547 399604 355548 399668
rect 355612 399604 355613 399668
rect 355547 399603 355613 399604
rect 355179 398036 355245 398037
rect 355179 397972 355180 398036
rect 355244 397972 355245 398036
rect 355179 397971 355245 397972
rect 355182 396541 355242 397971
rect 355550 397085 355610 399603
rect 357390 399397 357450 400147
rect 360518 399805 360578 401915
rect 360515 399804 360581 399805
rect 360515 399740 360516 399804
rect 360580 399740 360581 399804
rect 360515 399739 360581 399740
rect 360883 399804 360949 399805
rect 360883 399740 360884 399804
rect 360948 399740 360949 399804
rect 360883 399739 360949 399740
rect 358675 399668 358741 399669
rect 358675 399604 358676 399668
rect 358740 399604 358741 399668
rect 358675 399603 358741 399604
rect 360699 399668 360765 399669
rect 360699 399604 360700 399668
rect 360764 399604 360765 399668
rect 360699 399603 360765 399604
rect 357387 399396 357453 399397
rect 357387 399332 357388 399396
rect 357452 399332 357453 399396
rect 357387 399331 357453 399332
rect 358123 399260 358189 399261
rect 358123 399196 358124 399260
rect 358188 399196 358189 399260
rect 358123 399195 358189 399196
rect 357571 398172 357637 398173
rect 357571 398108 357572 398172
rect 357636 398108 357637 398172
rect 357571 398107 357637 398108
rect 357387 397900 357453 397901
rect 357387 397836 357388 397900
rect 357452 397836 357453 397900
rect 357387 397835 357453 397836
rect 356467 397492 356533 397493
rect 356467 397428 356468 397492
rect 356532 397428 356533 397492
rect 356467 397427 356533 397428
rect 355547 397084 355613 397085
rect 355547 397020 355548 397084
rect 355612 397020 355613 397084
rect 355547 397019 355613 397020
rect 355179 396540 355245 396541
rect 355179 396476 355180 396540
rect 355244 396476 355245 396540
rect 355179 396475 355245 396476
rect 354811 395996 354877 395997
rect 354811 395932 354812 395996
rect 354876 395932 354877 395996
rect 354811 395931 354877 395932
rect 354627 395316 354693 395317
rect 354627 395252 354628 395316
rect 354692 395252 354693 395316
rect 354627 395251 354693 395252
rect 354814 378045 354874 395931
rect 354811 378044 354877 378045
rect 354811 377980 354812 378044
rect 354876 377980 354877 378044
rect 354811 377979 354877 377980
rect 356470 308413 356530 397427
rect 357019 397084 357085 397085
rect 357019 397020 357020 397084
rect 357084 397020 357085 397084
rect 357019 397019 357085 397020
rect 356651 396812 356717 396813
rect 356651 396748 356652 396812
rect 356716 396748 356717 396812
rect 356651 396747 356717 396748
rect 356467 308412 356533 308413
rect 356467 308348 356468 308412
rect 356532 308348 356533 308412
rect 356467 308347 356533 308348
rect 356654 305829 356714 396747
rect 356835 395316 356901 395317
rect 356835 395252 356836 395316
rect 356900 395252 356901 395316
rect 356835 395251 356901 395252
rect 356838 313989 356898 395251
rect 357022 387157 357082 397019
rect 357390 396677 357450 397835
rect 357387 396676 357453 396677
rect 357387 396612 357388 396676
rect 357452 396612 357453 396676
rect 357387 396611 357453 396612
rect 357574 394501 357634 398107
rect 358126 397493 358186 399195
rect 358123 397492 358189 397493
rect 358123 397428 358124 397492
rect 358188 397428 358189 397492
rect 358123 397427 358189 397428
rect 358123 397220 358189 397221
rect 358123 397156 358124 397220
rect 358188 397156 358189 397220
rect 358123 397155 358189 397156
rect 357571 394500 357637 394501
rect 357571 394436 357572 394500
rect 357636 394436 357637 394500
rect 357571 394435 357637 394436
rect 357939 393548 358005 393549
rect 357939 393484 357940 393548
rect 358004 393484 358005 393548
rect 357939 393483 358005 393484
rect 357019 387156 357085 387157
rect 357019 387092 357020 387156
rect 357084 387092 357085 387156
rect 357019 387091 357085 387092
rect 356835 313988 356901 313989
rect 356835 313924 356836 313988
rect 356900 313924 356901 313988
rect 356835 313923 356901 313924
rect 357942 305965 358002 393483
rect 358126 306101 358186 397155
rect 358307 396676 358373 396677
rect 358307 396612 358308 396676
rect 358372 396612 358373 396676
rect 358307 396611 358373 396612
rect 358310 308821 358370 396611
rect 358678 392597 358738 399603
rect 360331 397764 360397 397765
rect 360331 397700 360332 397764
rect 360396 397700 360397 397764
rect 360331 397699 360397 397700
rect 359411 397492 359477 397493
rect 359411 397428 359412 397492
rect 359476 397428 359477 397492
rect 359411 397427 359477 397428
rect 358859 396948 358925 396949
rect 358859 396884 358860 396948
rect 358924 396884 358925 396948
rect 358859 396883 358925 396884
rect 358675 392596 358741 392597
rect 358675 392532 358676 392596
rect 358740 392532 358741 392596
rect 358675 392531 358741 392532
rect 358307 308820 358373 308821
rect 358307 308756 358308 308820
rect 358372 308756 358373 308820
rect 358307 308755 358373 308756
rect 358123 306100 358189 306101
rect 358123 306036 358124 306100
rect 358188 306036 358189 306100
rect 358123 306035 358189 306036
rect 357939 305964 358005 305965
rect 357939 305900 357940 305964
rect 358004 305900 358005 305964
rect 357939 305899 358005 305900
rect 356651 305828 356717 305829
rect 356651 305764 356652 305828
rect 356716 305764 356717 305828
rect 356651 305763 356717 305764
rect 358862 302157 358922 396883
rect 359414 307325 359474 397427
rect 360334 385661 360394 397699
rect 360331 385660 360397 385661
rect 360331 385596 360332 385660
rect 360396 385596 360397 385660
rect 360331 385595 360397 385596
rect 359411 307324 359477 307325
rect 359411 307260 359412 307324
rect 359476 307260 359477 307324
rect 359411 307259 359477 307260
rect 360702 304877 360762 399603
rect 360886 393277 360946 399739
rect 361794 399454 362414 434898
rect 362910 401165 362970 451283
rect 363275 449988 363341 449989
rect 363275 449924 363276 449988
rect 363340 449924 363341 449988
rect 363275 449923 363341 449924
rect 364379 449988 364445 449989
rect 364379 449924 364380 449988
rect 364444 449924 364445 449988
rect 364379 449923 364445 449924
rect 362907 401164 362973 401165
rect 362907 401100 362908 401164
rect 362972 401100 362973 401164
rect 362907 401099 362973 401100
rect 362539 399804 362605 399805
rect 362539 399740 362540 399804
rect 362604 399802 362605 399804
rect 363091 399804 363157 399805
rect 362604 399742 362786 399802
rect 362604 399740 362605 399742
rect 362539 399739 362605 399740
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 360883 393276 360949 393277
rect 360883 393212 360884 393276
rect 360948 393212 360949 393276
rect 360883 393211 360949 393212
rect 361794 363454 362414 398898
rect 362539 393412 362605 393413
rect 362539 393348 362540 393412
rect 362604 393348 362605 393412
rect 362539 393347 362605 393348
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 360699 304876 360765 304877
rect 360699 304812 360700 304876
rect 360764 304812 360765 304876
rect 360699 304811 360765 304812
rect 358859 302156 358925 302157
rect 358859 302092 358860 302156
rect 358924 302092 358925 302156
rect 358859 302091 358925 302092
rect 354443 295220 354509 295221
rect 354443 295156 354444 295220
rect 354508 295156 354509 295220
rect 354443 295155 354509 295156
rect 352051 295084 352117 295085
rect 352051 295020 352052 295084
rect 352116 295020 352117 295084
rect 352051 295019 352117 295020
rect 347819 294676 347885 294677
rect 347819 294612 347820 294676
rect 347884 294612 347885 294676
rect 347819 294611 347885 294612
rect 361794 291454 362414 326898
rect 362542 297669 362602 393347
rect 362726 307733 362786 399742
rect 363091 399740 363092 399804
rect 363156 399740 363157 399804
rect 363091 399739 363157 399740
rect 362907 396948 362973 396949
rect 362907 396884 362908 396948
rect 362972 396884 362973 396948
rect 362907 396883 362973 396884
rect 362723 307732 362789 307733
rect 362723 307668 362724 307732
rect 362788 307668 362789 307732
rect 362723 307667 362789 307668
rect 362910 297805 362970 396883
rect 363094 297941 363154 399739
rect 363278 384301 363338 449923
rect 364382 400077 364442 449923
rect 365514 439174 366134 474618
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 374131 452572 374197 452573
rect 374131 452508 374132 452572
rect 374196 452508 374197 452572
rect 374131 452507 374197 452508
rect 368243 451348 368309 451349
rect 368243 451284 368244 451348
rect 368308 451284 368309 451348
rect 368243 451283 368309 451284
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 364379 400076 364445 400077
rect 364379 400012 364380 400076
rect 364444 400012 364445 400076
rect 364379 400011 364445 400012
rect 364195 399804 364261 399805
rect 364195 399740 364196 399804
rect 364260 399740 364261 399804
rect 364195 399739 364261 399740
rect 363459 396540 363525 396541
rect 363459 396476 363460 396540
rect 363524 396476 363525 396540
rect 363459 396475 363525 396476
rect 363275 384300 363341 384301
rect 363275 384236 363276 384300
rect 363340 384236 363341 384300
rect 363275 384235 363341 384236
rect 363462 306237 363522 396475
rect 364198 393141 364258 399739
rect 365115 398716 365181 398717
rect 365115 398652 365116 398716
rect 365180 398652 365181 398716
rect 365115 398651 365181 398652
rect 364379 397356 364445 397357
rect 364379 397292 364380 397356
rect 364444 397292 364445 397356
rect 364379 397291 364445 397292
rect 364195 393140 364261 393141
rect 364195 393076 364196 393140
rect 364260 393076 364261 393140
rect 364195 393075 364261 393076
rect 364382 381989 364442 397291
rect 364931 393276 364997 393277
rect 364931 393212 364932 393276
rect 364996 393212 364997 393276
rect 364931 393211 364997 393212
rect 364379 381988 364445 381989
rect 364379 381924 364380 381988
rect 364444 381924 364445 381988
rect 364379 381923 364445 381924
rect 364934 306373 364994 393211
rect 365118 315621 365178 398651
rect 365514 367174 366134 402618
rect 366587 399940 366653 399941
rect 366587 399938 366588 399940
rect 366406 399878 366588 399938
rect 366219 399668 366285 399669
rect 366219 399604 366220 399668
rect 366284 399604 366285 399668
rect 366219 399603 366285 399604
rect 366222 393005 366282 399603
rect 366219 393004 366285 393005
rect 366219 392940 366220 393004
rect 366284 392940 366285 393004
rect 366219 392939 366285 392940
rect 366406 382125 366466 399878
rect 366587 399876 366588 399878
rect 366652 399876 366653 399940
rect 366587 399875 366653 399876
rect 366771 399940 366837 399941
rect 366771 399876 366772 399940
rect 366836 399876 366837 399940
rect 366771 399875 366837 399876
rect 368059 399940 368125 399941
rect 368059 399876 368060 399940
rect 368124 399876 368125 399940
rect 368059 399875 368125 399876
rect 366587 399804 366653 399805
rect 366587 399740 366588 399804
rect 366652 399740 366653 399804
rect 366587 399739 366653 399740
rect 366590 387701 366650 399739
rect 366774 393141 366834 399875
rect 367507 399804 367573 399805
rect 367507 399740 367508 399804
rect 367572 399740 367573 399804
rect 367507 399739 367573 399740
rect 366771 393140 366837 393141
rect 366771 393076 366772 393140
rect 366836 393076 366837 393140
rect 366771 393075 366837 393076
rect 367510 390570 367570 399739
rect 367875 397356 367941 397357
rect 367875 397292 367876 397356
rect 367940 397292 367941 397356
rect 367875 397291 367941 397292
rect 367878 393277 367938 397291
rect 367875 393276 367941 393277
rect 367875 393212 367876 393276
rect 367940 393212 367941 393276
rect 367875 393211 367941 393212
rect 367691 393140 367757 393141
rect 367691 393076 367692 393140
rect 367756 393076 367757 393140
rect 367691 393075 367757 393076
rect 367326 390510 367570 390570
rect 366587 387700 366653 387701
rect 366587 387636 366588 387700
rect 366652 387636 366653 387700
rect 366587 387635 366653 387636
rect 366403 382124 366469 382125
rect 366403 382060 366404 382124
rect 366468 382060 366469 382124
rect 366403 382059 366469 382060
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365115 315620 365181 315621
rect 365115 315556 365116 315620
rect 365180 315556 365181 315620
rect 365115 315555 365181 315556
rect 364931 306372 364997 306373
rect 364931 306308 364932 306372
rect 364996 306308 364997 306372
rect 364931 306307 364997 306308
rect 363459 306236 363525 306237
rect 363459 306172 363460 306236
rect 363524 306172 363525 306236
rect 363459 306171 363525 306172
rect 363091 297940 363157 297941
rect 363091 297876 363092 297940
rect 363156 297876 363157 297940
rect 363091 297875 363157 297876
rect 362907 297804 362973 297805
rect 362907 297740 362908 297804
rect 362972 297740 362973 297804
rect 362907 297739 362973 297740
rect 362539 297668 362605 297669
rect 362539 297604 362540 297668
rect 362604 297604 362605 297668
rect 362539 297603 362605 297604
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 338251 228988 338317 228989
rect 338251 228924 338252 228988
rect 338316 228924 338317 228988
rect 338251 228923 338317 228924
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 335859 59396 335925 59397
rect 335859 59332 335860 59396
rect 335924 59332 335925 59396
rect 335859 59331 335925 59332
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -1894 330134 -1862
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 295174 366134 330618
rect 367326 303381 367386 390510
rect 367694 318205 367754 393075
rect 368062 392869 368122 399875
rect 368246 399669 368306 451283
rect 374134 449581 374194 452507
rect 376891 451348 376957 451349
rect 376891 451284 376892 451348
rect 376956 451284 376957 451348
rect 376891 451283 376957 451284
rect 374131 449580 374197 449581
rect 374131 449516 374132 449580
rect 374196 449516 374197 449580
rect 374131 449515 374197 449516
rect 370451 449444 370517 449445
rect 370451 449380 370452 449444
rect 370516 449380 370517 449444
rect 370451 449379 370517 449380
rect 373211 449444 373277 449445
rect 373211 449380 373212 449444
rect 373276 449380 373277 449444
rect 373211 449379 373277 449380
rect 370454 400213 370514 449379
rect 371187 449308 371253 449309
rect 371187 449244 371188 449308
rect 371252 449244 371253 449308
rect 371187 449243 371253 449244
rect 371190 401573 371250 449243
rect 371187 401572 371253 401573
rect 371187 401508 371188 401572
rect 371252 401508 371253 401572
rect 371187 401507 371253 401508
rect 370451 400212 370517 400213
rect 370451 400148 370452 400212
rect 370516 400148 370517 400212
rect 370451 400147 370517 400148
rect 368427 399940 368493 399941
rect 368427 399876 368428 399940
rect 368492 399876 368493 399940
rect 368427 399875 368493 399876
rect 369715 399940 369781 399941
rect 369715 399876 369716 399940
rect 369780 399876 369781 399940
rect 369715 399875 369781 399876
rect 371003 399940 371069 399941
rect 371003 399876 371004 399940
rect 371068 399876 371069 399940
rect 371003 399875 371069 399876
rect 371187 399940 371253 399941
rect 371187 399876 371188 399940
rect 371252 399876 371253 399940
rect 371187 399875 371253 399876
rect 371739 399940 371805 399941
rect 371739 399876 371740 399940
rect 371804 399876 371805 399940
rect 371739 399875 371805 399876
rect 368243 399668 368309 399669
rect 368243 399604 368244 399668
rect 368308 399604 368309 399668
rect 368243 399603 368309 399604
rect 368430 399125 368490 399875
rect 368427 399124 368493 399125
rect 368427 399060 368428 399124
rect 368492 399060 368493 399124
rect 368427 399059 368493 399060
rect 368979 398036 369045 398037
rect 368979 397972 368980 398036
rect 369044 397972 369045 398036
rect 368979 397971 369045 397972
rect 368611 395588 368677 395589
rect 368611 395524 368612 395588
rect 368676 395524 368677 395588
rect 368611 395523 368677 395524
rect 368427 395180 368493 395181
rect 368427 395116 368428 395180
rect 368492 395116 368493 395180
rect 368427 395115 368493 395116
rect 368059 392868 368125 392869
rect 368059 392804 368060 392868
rect 368124 392804 368125 392868
rect 368059 392803 368125 392804
rect 368430 329357 368490 395115
rect 368614 381717 368674 395523
rect 368611 381716 368677 381717
rect 368611 381652 368612 381716
rect 368676 381652 368677 381716
rect 368611 381651 368677 381652
rect 368427 329356 368493 329357
rect 368427 329292 368428 329356
rect 368492 329292 368493 329356
rect 368427 329291 368493 329292
rect 367691 318204 367757 318205
rect 367691 318140 367692 318204
rect 367756 318140 367757 318204
rect 367691 318139 367757 318140
rect 367323 303380 367389 303381
rect 367323 303316 367324 303380
rect 367388 303316 367389 303380
rect 367323 303315 367389 303316
rect 368982 297533 369042 397971
rect 369163 397356 369229 397357
rect 369163 397292 369164 397356
rect 369228 397292 369229 397356
rect 369163 397291 369229 397292
rect 369166 307461 369226 397291
rect 369718 393413 369778 399875
rect 369899 399804 369965 399805
rect 369899 399740 369900 399804
rect 369964 399740 369965 399804
rect 369899 399739 369965 399740
rect 369715 393412 369781 393413
rect 369715 393348 369716 393412
rect 369780 393348 369781 393412
rect 369715 393347 369781 393348
rect 369902 318069 369962 399739
rect 370451 399532 370517 399533
rect 370451 399468 370452 399532
rect 370516 399468 370517 399532
rect 370451 399467 370517 399468
rect 369899 318068 369965 318069
rect 369899 318004 369900 318068
rect 369964 318004 369965 318068
rect 369899 318003 369965 318004
rect 369163 307460 369229 307461
rect 369163 307396 369164 307460
rect 369228 307396 369229 307460
rect 369163 307395 369229 307396
rect 370454 299029 370514 399467
rect 371006 398717 371066 399875
rect 371003 398716 371069 398717
rect 371003 398652 371004 398716
rect 371068 398652 371069 398716
rect 371003 398651 371069 398652
rect 371190 391781 371250 399875
rect 371555 399804 371621 399805
rect 371555 399740 371556 399804
rect 371620 399740 371621 399804
rect 371555 399739 371621 399740
rect 371187 391780 371253 391781
rect 371187 391716 371188 391780
rect 371252 391716 371253 391780
rect 371187 391715 371253 391716
rect 371558 390570 371618 399739
rect 371742 399125 371802 399875
rect 372843 399804 372909 399805
rect 372843 399740 372844 399804
rect 372908 399740 372909 399804
rect 372843 399739 372909 399740
rect 372291 399668 372357 399669
rect 372291 399604 372292 399668
rect 372356 399604 372357 399668
rect 372291 399603 372357 399604
rect 371739 399124 371805 399125
rect 371739 399060 371740 399124
rect 371804 399060 371805 399124
rect 371739 399059 371805 399060
rect 371739 398988 371805 398989
rect 371739 398924 371740 398988
rect 371804 398924 371805 398988
rect 371739 398923 371805 398924
rect 371374 390510 371618 390570
rect 371374 325413 371434 390510
rect 371742 381853 371802 398923
rect 372294 397629 372354 399603
rect 372291 397628 372357 397629
rect 372291 397564 372292 397628
rect 372356 397564 372357 397628
rect 372291 397563 372357 397564
rect 372846 397493 372906 399739
rect 373214 399261 373274 449379
rect 374134 400077 374194 449515
rect 374315 449444 374381 449445
rect 374315 449380 374316 449444
rect 374380 449380 374381 449444
rect 374315 449379 374381 449380
rect 374318 400893 374378 449379
rect 374315 400892 374381 400893
rect 374315 400828 374316 400892
rect 374380 400828 374381 400892
rect 374315 400827 374381 400828
rect 374131 400076 374197 400077
rect 374131 400012 374132 400076
rect 374196 400012 374197 400076
rect 374131 400011 374197 400012
rect 374315 399940 374381 399941
rect 374315 399876 374316 399940
rect 374380 399876 374381 399940
rect 374315 399875 374381 399876
rect 373211 399260 373277 399261
rect 373211 399196 373212 399260
rect 373276 399196 373277 399260
rect 373211 399195 373277 399196
rect 373947 399260 374013 399261
rect 373947 399196 373948 399260
rect 374012 399196 374013 399260
rect 373947 399195 374013 399196
rect 372843 397492 372909 397493
rect 372843 397428 372844 397492
rect 372908 397428 372909 397492
rect 372843 397427 372909 397428
rect 372291 397220 372357 397221
rect 372291 397156 372292 397220
rect 372356 397156 372357 397220
rect 372291 397155 372357 397156
rect 372294 394637 372354 397155
rect 373763 395452 373829 395453
rect 373763 395388 373764 395452
rect 373828 395388 373829 395452
rect 373763 395387 373829 395388
rect 372291 394636 372357 394637
rect 372291 394572 372292 394636
rect 372356 394572 372357 394636
rect 372291 394571 372357 394572
rect 372659 393956 372725 393957
rect 372659 393892 372660 393956
rect 372724 393892 372725 393956
rect 372659 393891 372725 393892
rect 371739 381852 371805 381853
rect 371739 381788 371740 381852
rect 371804 381788 371805 381852
rect 371739 381787 371805 381788
rect 372662 371925 372722 393891
rect 372659 371924 372725 371925
rect 372659 371860 372660 371924
rect 372724 371860 372725 371924
rect 372659 371859 372725 371860
rect 371371 325412 371437 325413
rect 371371 325348 371372 325412
rect 371436 325348 371437 325412
rect 371371 325347 371437 325348
rect 373766 324461 373826 395387
rect 373950 389197 374010 399195
rect 374318 397085 374378 399875
rect 374867 399804 374933 399805
rect 374867 399740 374868 399804
rect 374932 399740 374933 399804
rect 374867 399739 374933 399740
rect 374315 397084 374381 397085
rect 374315 397020 374316 397084
rect 374380 397020 374381 397084
rect 374315 397019 374381 397020
rect 374131 395452 374197 395453
rect 374131 395388 374132 395452
rect 374196 395388 374197 395452
rect 374131 395387 374197 395388
rect 373947 389196 374013 389197
rect 373947 389132 373948 389196
rect 374012 389132 374013 389196
rect 373947 389131 374013 389132
rect 373947 383892 374013 383893
rect 373947 383828 373948 383892
rect 374012 383828 374013 383892
rect 373947 383827 374013 383828
rect 373950 383485 374010 383827
rect 373947 383484 374013 383485
rect 373947 383420 373948 383484
rect 374012 383420 374013 383484
rect 373947 383419 374013 383420
rect 373947 374100 374013 374101
rect 373947 374036 373948 374100
rect 374012 374036 374013 374100
rect 373947 374035 374013 374036
rect 373950 373829 374010 374035
rect 373947 373828 374013 373829
rect 373947 373764 373948 373828
rect 374012 373764 374013 373828
rect 373947 373763 374013 373764
rect 373947 364444 374013 364445
rect 373947 364380 373948 364444
rect 374012 364380 374013 364444
rect 373947 364379 374013 364380
rect 373950 364173 374010 364379
rect 373947 364172 374013 364173
rect 373947 364108 373948 364172
rect 374012 364108 374013 364172
rect 373947 364107 374013 364108
rect 373947 354788 374013 354789
rect 373947 354724 373948 354788
rect 374012 354724 374013 354788
rect 373947 354723 374013 354724
rect 373950 354517 374010 354723
rect 373947 354516 374013 354517
rect 373947 354452 373948 354516
rect 374012 354452 374013 354516
rect 373947 354451 374013 354452
rect 373947 345132 374013 345133
rect 373947 345068 373948 345132
rect 374012 345068 374013 345132
rect 373947 345067 374013 345068
rect 373950 344997 374010 345067
rect 373947 344996 374013 344997
rect 373947 344932 373948 344996
rect 374012 344932 374013 344996
rect 373947 344931 374013 344932
rect 373947 340780 374013 340781
rect 373947 340716 373948 340780
rect 374012 340716 374013 340780
rect 373947 340715 374013 340716
rect 373950 331261 374010 340715
rect 373947 331260 374013 331261
rect 373947 331196 373948 331260
rect 374012 331196 374013 331260
rect 373947 331195 374013 331196
rect 374134 326501 374194 395387
rect 374870 390570 374930 399739
rect 375971 397900 376037 397901
rect 375971 397836 375972 397900
rect 376036 397836 376037 397900
rect 375971 397835 376037 397836
rect 375419 397356 375485 397357
rect 375419 397292 375420 397356
rect 375484 397292 375485 397356
rect 375419 397291 375485 397292
rect 374870 390510 375298 390570
rect 375238 328541 375298 390510
rect 375235 328540 375301 328541
rect 375235 328476 375236 328540
rect 375300 328476 375301 328540
rect 375235 328475 375301 328476
rect 375238 327725 375298 328475
rect 375235 327724 375301 327725
rect 375235 327660 375236 327724
rect 375300 327660 375301 327724
rect 375235 327659 375301 327660
rect 374131 326500 374197 326501
rect 374131 326436 374132 326500
rect 374196 326436 374197 326500
rect 374131 326435 374197 326436
rect 373947 325956 374013 325957
rect 373947 325892 373948 325956
rect 374012 325892 374013 325956
rect 373947 325891 374013 325892
rect 373950 325710 374010 325891
rect 373950 325650 374194 325710
rect 374134 325277 374194 325650
rect 374131 325276 374197 325277
rect 374131 325212 374132 325276
rect 374196 325212 374197 325276
rect 374131 325211 374197 325212
rect 373763 324460 373829 324461
rect 373763 324396 373764 324460
rect 373828 324396 373829 324460
rect 373763 324395 373829 324396
rect 375422 299437 375482 397291
rect 375974 310045 376034 397835
rect 376894 385797 376954 451283
rect 384987 449444 385053 449445
rect 384987 449380 384988 449444
rect 385052 449380 385053 449444
rect 384987 449379 385053 449380
rect 382227 449308 382293 449309
rect 382227 449244 382228 449308
rect 382292 449244 382293 449308
rect 382227 449243 382293 449244
rect 383699 449308 383765 449309
rect 383699 449244 383700 449308
rect 383764 449244 383765 449308
rect 383699 449243 383765 449244
rect 378363 400212 378429 400213
rect 378363 400148 378364 400212
rect 378428 400148 378429 400212
rect 378363 400147 378429 400148
rect 377627 399940 377693 399941
rect 377627 399876 377628 399940
rect 377692 399876 377693 399940
rect 377627 399875 377693 399876
rect 377259 397764 377325 397765
rect 377259 397700 377260 397764
rect 377324 397700 377325 397764
rect 377259 397699 377325 397700
rect 376891 385796 376957 385797
rect 376891 385732 376892 385796
rect 376956 385732 376957 385796
rect 376891 385731 376957 385732
rect 375971 310044 376037 310045
rect 375971 309980 375972 310044
rect 376036 309980 376037 310044
rect 375971 309979 376037 309980
rect 377262 304605 377322 397699
rect 377630 396541 377690 399875
rect 378179 399804 378245 399805
rect 378179 399740 378180 399804
rect 378244 399740 378245 399804
rect 378179 399739 378245 399740
rect 378182 396813 378242 399739
rect 378179 396812 378245 396813
rect 378179 396748 378180 396812
rect 378244 396748 378245 396812
rect 378179 396747 378245 396748
rect 378179 396676 378245 396677
rect 378179 396612 378180 396676
rect 378244 396612 378245 396676
rect 378179 396611 378245 396612
rect 377627 396540 377693 396541
rect 377627 396476 377628 396540
rect 377692 396476 377693 396540
rect 377627 396475 377693 396476
rect 378182 326637 378242 396611
rect 378366 393549 378426 400147
rect 379283 400076 379349 400077
rect 379283 400012 379284 400076
rect 379348 400012 379349 400076
rect 379283 400011 379349 400012
rect 381675 400076 381741 400077
rect 381675 400012 381676 400076
rect 381740 400012 381741 400076
rect 381675 400011 381741 400012
rect 379099 399940 379165 399941
rect 379099 399876 379100 399940
rect 379164 399876 379165 399940
rect 379099 399875 379165 399876
rect 378547 399532 378613 399533
rect 378547 399468 378548 399532
rect 378612 399468 378613 399532
rect 378547 399467 378613 399468
rect 378363 393548 378429 393549
rect 378363 393484 378364 393548
rect 378428 393484 378429 393548
rect 378363 393483 378429 393484
rect 378550 389333 378610 399467
rect 379102 395181 379162 399875
rect 379099 395180 379165 395181
rect 379099 395116 379100 395180
rect 379164 395116 379165 395180
rect 379099 395115 379165 395116
rect 378547 389332 378613 389333
rect 378547 389268 378548 389332
rect 378612 389268 378613 389332
rect 378547 389267 378613 389268
rect 379286 389190 379346 400011
rect 379835 399804 379901 399805
rect 379835 399740 379836 399804
rect 379900 399740 379901 399804
rect 379835 399739 379901 399740
rect 379838 396677 379898 399739
rect 380939 397628 381005 397629
rect 380939 397564 380940 397628
rect 381004 397564 381005 397628
rect 380939 397563 381005 397564
rect 379835 396676 379901 396677
rect 379835 396612 379836 396676
rect 379900 396612 379901 396676
rect 379835 396611 379901 396612
rect 379651 395316 379717 395317
rect 379651 395252 379652 395316
rect 379716 395252 379717 395316
rect 379651 395251 379717 395252
rect 379286 389130 379530 389190
rect 379470 340890 379530 389130
rect 379654 367709 379714 395251
rect 379651 367708 379717 367709
rect 379651 367644 379652 367708
rect 379716 367644 379717 367708
rect 379651 367643 379717 367644
rect 379286 340830 379530 340890
rect 379286 337381 379346 340830
rect 379283 337380 379349 337381
rect 379283 337316 379284 337380
rect 379348 337316 379349 337380
rect 379283 337315 379349 337316
rect 378179 326636 378245 326637
rect 378179 326572 378180 326636
rect 378244 326572 378245 326636
rect 378179 326571 378245 326572
rect 380942 307597 381002 397563
rect 381678 345677 381738 400011
rect 382230 399397 382290 449243
rect 382411 399940 382477 399941
rect 382411 399876 382412 399940
rect 382476 399876 382477 399940
rect 382411 399875 382477 399876
rect 382227 399396 382293 399397
rect 382227 399332 382228 399396
rect 382292 399332 382293 399396
rect 382227 399331 382293 399332
rect 382227 397628 382293 397629
rect 382227 397564 382228 397628
rect 382292 397564 382293 397628
rect 382227 397563 382293 397564
rect 382043 397492 382109 397493
rect 382043 397428 382044 397492
rect 382108 397428 382109 397492
rect 382043 397427 382109 397428
rect 381675 345676 381741 345677
rect 381675 345612 381676 345676
rect 381740 345612 381741 345676
rect 381675 345611 381741 345612
rect 382046 329901 382106 397427
rect 382043 329900 382109 329901
rect 382043 329836 382044 329900
rect 382108 329836 382109 329900
rect 382043 329835 382109 329836
rect 382230 325005 382290 397563
rect 382414 397357 382474 399875
rect 382411 397356 382477 397357
rect 382411 397292 382412 397356
rect 382476 397292 382477 397356
rect 382411 397291 382477 397292
rect 382779 397356 382845 397357
rect 382779 397292 382780 397356
rect 382844 397292 382845 397356
rect 382779 397291 382845 397292
rect 382782 342957 382842 397291
rect 383702 388517 383762 449243
rect 383699 388516 383765 388517
rect 383699 388452 383700 388516
rect 383764 388452 383765 388516
rect 383699 388451 383765 388452
rect 384990 388381 385050 449379
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 384987 388380 385053 388381
rect 384987 388316 384988 388380
rect 385052 388316 385053 388380
rect 384987 388315 385053 388316
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 382779 342956 382845 342957
rect 382779 342892 382780 342956
rect 382844 342892 382845 342956
rect 382779 342891 382845 342892
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 382227 325004 382293 325005
rect 382227 324940 382228 325004
rect 382292 324940 382293 325004
rect 382227 324939 382293 324940
rect 380939 307596 381005 307597
rect 380939 307532 380940 307596
rect 381004 307532 381005 307596
rect 380939 307531 381005 307532
rect 377259 304604 377325 304605
rect 377259 304540 377260 304604
rect 377324 304540 377325 304604
rect 377259 304539 377325 304540
rect 375419 299436 375485 299437
rect 375419 299372 375420 299436
rect 375484 299372 375485 299436
rect 375419 299371 375485 299372
rect 370451 299028 370517 299029
rect 370451 298964 370452 299028
rect 370516 298964 370517 299028
rect 370451 298963 370517 298964
rect 368979 297532 369045 297533
rect 368979 297468 368980 297532
rect 369044 297468 369045 297532
rect 368979 297467 369045 297468
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -1894 366134 -1862
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 705798 402134 705830
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -1894 402134 -1862
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 705798 438134 705830
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -1894 438134 -1862
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 705798 474134 705830
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -1894 474134 -1862
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 705798 510134 705830
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -1894 510134 -1862
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 705798 546134 705830
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -1894 546134 -1862
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 705798 582134 705830
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -1894 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 164250 183218 164486 183454
rect 164250 182898 164486 183134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 179610 186938 179846 187174
rect 179610 186618 179846 186854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 194970 183218 195206 183454
rect 194970 182898 195206 183134
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 691174 586890 691206
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect -2966 690854 586890 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect -2966 690586 586890 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 655174 586890 655206
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect -2966 654854 586890 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect -2966 654586 586890 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 619174 586890 619206
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect -2966 618854 586890 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect -2966 618586 586890 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -2966 583174 586890 583206
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect -2966 582854 586890 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect -2966 582586 586890 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 547174 586890 547206
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect -2966 546854 586890 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect -2966 546586 586890 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 511174 586890 511206
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect -2966 510854 586890 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect -2966 510586 586890 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -2966 475174 586890 475206
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect -2966 474854 586890 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect -2966 474586 586890 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -2966 439174 586890 439206
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect -2966 438854 586890 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect -2966 438586 586890 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -2966 403174 586890 403206
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect -2966 402854 586890 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect -2966 402586 586890 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -2966 367174 586890 367206
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect -2966 366854 586890 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect -2966 366586 586890 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -2966 331174 586890 331206
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect -2966 330854 586890 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect -2966 330586 586890 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 295174 586890 295206
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect -2966 294854 586890 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect -2966 294586 586890 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -2966 259174 586890 259206
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect -2966 258854 586890 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect -2966 258586 586890 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 223174 586890 223206
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect -2966 222854 586890 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect -2966 222586 586890 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 187174 586890 187206
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 179610 187174
rect 179846 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect -2966 186854 586890 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 179610 186854
rect 179846 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect -2966 186586 586890 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 164250 183454
rect 164486 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 194970 183454
rect 195206 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 164250 183134
rect 164486 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 194970 183134
rect 195206 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -2966 151174 586890 151206
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect -2966 150854 586890 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect -2966 150586 586890 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 115174 586890 115206
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect -2966 114854 586890 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect -2966 114586 586890 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 79174 586890 79206
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect -2966 78854 586890 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect -2966 78586 586890 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -2966 43174 586890 43206
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect -2966 42854 586890 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect -2966 42586 586890 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 7174 586890 7206
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect -2966 6854 586890 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect -2966 6586 586890 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use macro_2to3  u_macro_2to3
timestamp 0
transform 1 0 280000 0 1 320000
box 1066 0 48890 50000
use macro_2xdrive  u_macro_2xdrive
timestamp 0
transform 1 0 220000 0 1 240000
box 1066 0 48890 50000
use macro_and_inv  u_macro_and_inv
timestamp 0
transform 1 0 340000 0 1 400000
box 1066 0 48890 50000
use macro_golden  u_macro_golden
timestamp 0
transform 1 0 160000 0 1 160000
box 1066 0 48890 50000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -1894 2414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -1894 38414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -1894 74414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -1894 110414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -1894 146414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -1894 182414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -1894 218414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -1894 254414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -1894 290414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -1894 326414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -1894 362414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -1894 398414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -1894 434414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -1894 470414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -1894 506414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -1894 542414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -1894 578414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 2866 586890 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 38866 586890 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 74866 586890 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 110866 586890 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 146866 586890 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 182866 586890 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 218866 586890 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 254866 586890 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 290866 586890 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 326866 586890 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 362866 586890 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 398866 586890 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 434866 586890 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 470866 586890 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 506866 586890 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 542866 586890 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 578866 586890 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 614866 586890 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 650866 586890 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 686866 586890 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 5514 -1894 6134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 41514 -1894 42134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 77514 -1894 78134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 113514 -1894 114134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 149514 -1894 150134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 185514 -1894 186134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 221514 -1894 222134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 257514 -1894 258134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 293514 -1894 294134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 329514 -1894 330134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 365514 -1894 366134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 401514 -1894 402134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 437514 -1894 438134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 473514 -1894 474134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 509514 -1894 510134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 545514 -1894 546134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 581514 -1894 582134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 6586 586890 7206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 42586 586890 43206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 78586 586890 79206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 114586 586890 115206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 150586 586890 151206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 186586 586890 187206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 222586 586890 223206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 258586 586890 259206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 294586 586890 295206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 330586 586890 331206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 366586 586890 367206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 402586 586890 403206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 438586 586890 439206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 474586 586890 475206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 510586 586890 511206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 546586 586890 547206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 582586 586890 583206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 618586 586890 619206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 654586 586890 655206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 690586 586890 691206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 533 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 534 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 535 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 536 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 537 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 538 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 539 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 540 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 541 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 542 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 543 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 544 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 545 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 546 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 547 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 548 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 549 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 550 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 551 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 552 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 553 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 554 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 555 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 556 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 557 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 558 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 559 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 560 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 561 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 562 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 563 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 564 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 565 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 566 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 567 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 568 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 569 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 570 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 571 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 572 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 573 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 574 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 575 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 576 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 577 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 578 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 579 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 580 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 581 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 582 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 583 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 584 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 585 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 586 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 587 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 588 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 589 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 590 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 591 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 592 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 593 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 594 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 595 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 596 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 597 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 598 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 599 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 600 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 601 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 602 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 603 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 604 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 605 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 606 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 607 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 608 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 609 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 610 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 611 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 612 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 613 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 614 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 615 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 616 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 617 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 618 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 619 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 620 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 621 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 622 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 623 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 624 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 625 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 626 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 627 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 628 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 629 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 630 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 631 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 632 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 633 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 634 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 635 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 636 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 637 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 638 nsew signal input
rlabel via4 195088 183336 195088 183336 0 vccd1
rlabel via4 185984 187056 185984 187056 0 vssd1
rlabel metal3 581954 6596 581954 6596 0 io_in[0]
rlabel metal2 175398 210926 175398 210926 0 io_in[10]
rlabel metal2 176502 211062 176502 211062 0 io_in[11]
rlabel metal2 177606 211198 177606 211198 0 io_in[12]
rlabel metal2 178565 209916 178565 209916 0 io_in[13]
rlabel metal2 179814 211096 179814 211096 0 io_in[14]
rlabel metal2 558946 580625 558946 580625 0 io_in[15]
rlabel metal2 214682 254388 214682 254388 0 io_in[16]
rlabel metal2 214774 255306 214774 255306 0 io_in[17]
rlabel metal2 365010 701124 365010 701124 0 io_in[18]
rlabel metal2 185281 209916 185281 209916 0 io_in[19]
rlabel metal3 581908 46308 581908 46308 0 io_in[1]
rlabel metal2 234830 703596 234830 703596 0 io_in[20]
rlabel metal2 215050 255714 215050 255714 0 io_in[21]
rlabel metal2 273286 465392 273286 465392 0 io_in[22]
rlabel metal2 40204 703596 40204 703596 0 io_in[23]
rlabel metal2 190755 209916 190755 209916 0 io_in[24]
rlabel metal2 191905 209916 191905 209916 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1648 527884 1648 527884 0 io_in[27]
rlabel metal2 195125 209916 195125 209916 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal3 581908 86156 581908 86156 0 io_in[2]
rlabel metal3 1786 371348 1786 371348 0 io_in[30]
rlabel metal3 1878 319260 1878 319260 0 io_in[31]
rlabel metal3 1694 267172 1694 267172 0 io_in[32]
rlabel metal3 1740 214948 1740 214948 0 io_in[33]
rlabel metal2 191774 210868 191774 210868 0 io_in[34]
rlabel metal3 1832 110636 1832 110636 0 io_in[35]
rlabel metal2 383978 449956 383978 449956 0 io_in[36]
rlabel metal2 385128 449956 385128 449956 0 io_in[37]
rlabel metal3 582046 126004 582046 126004 0 io_in[3]
rlabel metal2 218546 209372 218546 209372 0 io_in[4]
rlabel metal2 229862 291166 229862 291166 0 io_in[5]
rlabel metal2 230867 289884 230867 289884 0 io_in[6]
rlabel metal2 172086 210960 172086 210960 0 io_in[7]
rlabel metal2 173045 209916 173045 209916 0 io_in[8]
rlabel metal2 174294 210314 174294 210314 0 io_in[9]
rlabel via2 580198 33099 580198 33099 0 io_oeb[0]
rlabel metal2 175766 211028 175766 211028 0 io_oeb[10]
rlabel metal2 176771 209916 176771 209916 0 io_oeb[11]
rlabel metal2 177829 209916 177829 209916 0 io_oeb[12]
rlabel metal2 178933 209916 178933 209916 0 io_oeb[13]
rlabel metal2 180037 209916 180037 209916 0 io_oeb[14]
rlabel metal2 527206 586714 527206 586714 0 io_oeb[15]
rlabel metal2 462346 579812 462346 579812 0 io_oeb[16]
rlabel metal2 183349 209916 183349 209916 0 io_oeb[17]
rlabel metal2 332534 701940 332534 701940 0 io_oeb[18]
rlabel metal2 185557 209916 185557 209916 0 io_oeb[19]
rlabel metal3 583556 72352 583556 72352 0 io_oeb[1]
rlabel metal2 306406 415140 306406 415140 0 io_oeb[20]
rlabel metal2 137172 703596 137172 703596 0 io_oeb[21]
rlabel metal3 233956 289408 233956 289408 0 io_oeb[22]
rlabel metal2 370040 449956 370040 449956 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal2 192181 209916 192181 209916 0 io_oeb[25]
rlabel metal2 193430 213000 193430 213000 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1740 449548 1740 449548 0 io_oeb[28]
rlabel metal2 256726 290826 256726 290826 0 io_oeb[29]
rlabel metal4 331844 240924 331844 240924 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 1832 241060 1832 241060 0 io_oeb[32]
rlabel metal3 1832 188836 1832 188836 0 io_oeb[33]
rlabel metal3 1694 136748 1694 136748 0 io_oeb[34]
rlabel metal3 1924 84660 1924 84660 0 io_oeb[35]
rlabel metal3 1924 45492 1924 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 276046 368577 276046 368577 0 io_oeb[3]
rlabel metal2 229126 292050 229126 292050 0 io_oeb[4]
rlabel metal2 230230 292152 230230 292152 0 io_oeb[5]
rlabel metal2 171297 209916 171297 209916 0 io_oeb[6]
rlabel metal2 172309 209916 172309 209916 0 io_oeb[7]
rlabel metal2 173413 209916 173413 209916 0 io_oeb[8]
rlabel metal2 174662 210994 174662 210994 0 io_oeb[9]
rlabel metal1 334282 369002 334282 369002 0 io_out[0]
rlabel metal2 175989 209916 175989 209916 0 io_out[10]
rlabel metal2 177238 211674 177238 211674 0 io_out[11]
rlabel metal2 178243 209916 178243 209916 0 io_out[12]
rlabel metal2 179446 253562 179446 253562 0 io_out[13]
rlabel metal2 180550 210960 180550 210960 0 io_out[14]
rlabel metal2 542386 583379 542386 583379 0 io_out[15]
rlabel metal2 182613 209916 182613 209916 0 io_out[16]
rlabel metal3 333477 384268 333477 384268 0 io_out[17]
rlabel metal2 348818 701974 348818 701974 0 io_out[18]
rlabel metal2 186070 212082 186070 212082 0 io_out[19]
rlabel metal2 166053 209916 166053 209916 0 io_out[1]
rlabel metal2 219006 701634 219006 701634 0 io_out[20]
rlabel metal2 153226 538193 153226 538193 0 io_out[21]
rlabel metal2 189283 209916 189283 209916 0 io_out[22]
rlabel metal2 190539 209916 190539 209916 0 io_out[23]
rlabel metal2 191445 209916 191445 209916 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal2 254787 289884 254787 289884 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 2200 410516 2200 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal3 1740 358428 1740 358428 0 io_out[30]
rlabel metal3 2200 306204 2200 306204 0 io_out[31]
rlabel metal3 1878 254116 1878 254116 0 io_out[32]
rlabel metal3 1832 201892 1832 201892 0 io_out[33]
rlabel metal1 272228 291686 272228 291686 0 io_out[34]
rlabel metal3 1970 97580 1970 97580 0 io_out[35]
rlabel metal3 1694 58548 1694 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel metal3 581908 139332 581908 139332 0 io_out[3]
rlabel metal2 229494 290843 229494 290843 0 io_out[4]
rlabel metal1 230920 296174 230920 296174 0 io_out[5]
rlabel metal2 171573 209916 171573 209916 0 io_out[6]
rlabel metal2 172723 209916 172723 209916 0 io_out[7]
rlabel metal2 233811 289884 233811 289884 0 io_out[8]
rlabel metal2 174885 209916 174885 209916 0 io_out[9]
rlabel metal2 291134 307462 291134 307462 0 la_data_in[0]
rlabel metal2 270434 129370 270434 129370 0 la_data_in[100]
rlabel metal1 269606 154122 269606 154122 0 la_data_in[101]
rlabel metal2 487409 340 487409 340 0 la_data_in[102]
rlabel metal2 274114 126582 274114 126582 0 la_data_in[103]
rlabel metal2 270250 157080 270250 157080 0 la_data_in[104]
rlabel metal2 365654 398191 365654 398191 0 la_data_in[105]
rlabel metal2 501577 340 501577 340 0 la_data_in[106]
rlabel metal2 331338 279021 331338 279021 0 la_data_in[107]
rlabel metal1 287822 154122 287822 154122 0 la_data_in[108]
rlabel metal2 269054 152796 269054 152796 0 la_data_in[109]
rlabel metal1 160724 11798 160724 11798 0 la_data_in[10]
rlabel metal3 294584 236028 294584 236028 0 la_data_in[110]
rlabel metal2 269790 155020 269790 155020 0 la_data_in[111]
rlabel metal2 271814 155516 271814 155516 0 la_data_in[112]
rlabel metal2 526417 340 526417 340 0 la_data_in[113]
rlabel metal2 330418 309808 330418 309808 0 la_data_in[114]
rlabel metal2 270342 144432 270342 144432 0 la_data_in[115]
rlabel metal2 333178 274941 333178 274941 0 la_data_in[116]
rlabel metal2 273838 152830 273838 152830 0 la_data_in[117]
rlabel metal2 331522 277066 331522 277066 0 la_data_in[118]
rlabel metal2 547906 1911 547906 1911 0 la_data_in[119]
rlabel metal2 164910 1928 164910 1928 0 la_data_in[11]
rlabel metal2 269054 141644 269054 141644 0 la_data_in[120]
rlabel metal1 238970 137870 238970 137870 0 la_data_in[121]
rlabel metal2 288282 309315 288282 309315 0 la_data_in[122]
rlabel metal2 295366 147288 295366 147288 0 la_data_in[123]
rlabel metal2 565425 340 565425 340 0 la_data_in[124]
rlabel metal2 272274 135932 272274 135932 0 la_data_in[125]
rlabel metal2 271814 134878 271814 134878 0 la_data_in[126]
rlabel metal2 331430 277236 331430 277236 0 la_data_in[127]
rlabel metal2 175398 155992 175398 155992 0 la_data_in[12]
rlabel metal2 171994 1911 171994 1911 0 la_data_in[13]
rlabel metal2 175444 16560 175444 16560 0 la_data_in[14]
rlabel metal2 179078 1792 179078 1792 0 la_data_in[15]
rlabel metal2 182383 340 182383 340 0 la_data_in[16]
rlabel metal2 185978 16560 185978 16560 0 la_data_in[17]
rlabel metal2 177146 158892 177146 158892 0 la_data_in[18]
rlabel metal1 180090 3536 180090 3536 0 la_data_in[19]
rlabel metal2 129161 340 129161 340 0 la_data_in[1]
rlabel metal2 196834 1996 196834 1996 0 la_data_in[20]
rlabel metal2 200330 2200 200330 2200 0 la_data_in[21]
rlabel metal3 178779 157964 178779 157964 0 la_data_in[22]
rlabel metal1 186645 3366 186645 3366 0 la_data_in[23]
rlabel metal2 211002 2234 211002 2234 0 la_data_in[24]
rlabel metal2 213900 157012 213900 157012 0 la_data_in[25]
rlabel metal2 218086 1894 218086 1894 0 la_data_in[26]
rlabel metal2 211830 80138 211830 80138 0 la_data_in[27]
rlabel metal1 212842 155074 212842 155074 0 la_data_in[28]
rlabel metal2 228758 1962 228758 1962 0 la_data_in[29]
rlabel metal2 132756 16560 132756 16560 0 la_data_in[2]
rlabel metal2 232254 1724 232254 1724 0 la_data_in[30]
rlabel metal1 180642 157930 180642 157930 0 la_data_in[31]
rlabel metal1 217580 152694 217580 152694 0 la_data_in[32]
rlabel metal2 242926 1996 242926 1996 0 la_data_in[33]
rlabel metal2 287822 270708 287822 270708 0 la_data_in[34]
rlabel metal2 250010 2166 250010 2166 0 la_data_in[35]
rlabel metal2 253506 1962 253506 1962 0 la_data_in[36]
rlabel metal2 257094 2132 257094 2132 0 la_data_in[37]
rlabel metal2 250470 77214 250470 77214 0 la_data_in[38]
rlabel metal2 253414 16560 253414 16560 0 la_data_in[39]
rlabel metal2 136482 1894 136482 1894 0 la_data_in[3]
rlabel metal2 267766 2132 267766 2132 0 la_data_in[40]
rlabel metal2 271262 2098 271262 2098 0 la_data_in[41]
rlabel metal2 274850 1860 274850 1860 0 la_data_in[42]
rlabel metal2 271814 233716 271814 233716 0 la_data_in[43]
rlabel metal2 281934 1860 281934 1860 0 la_data_in[44]
rlabel metal2 285430 1758 285430 1758 0 la_data_in[45]
rlabel metal2 289018 1928 289018 1928 0 la_data_in[46]
rlabel metal2 292606 1962 292606 1962 0 la_data_in[47]
rlabel metal1 276506 229738 276506 229738 0 la_data_in[48]
rlabel metal2 296010 77316 296010 77316 0 la_data_in[49]
rlabel metal2 139833 340 139833 340 0 la_data_in[4]
rlabel metal2 303186 2030 303186 2030 0 la_data_in[50]
rlabel metal2 306774 2132 306774 2132 0 la_data_in[51]
rlabel metal2 310270 1758 310270 1758 0 la_data_in[52]
rlabel metal2 313858 1860 313858 1860 0 la_data_in[53]
rlabel metal2 314042 72080 314042 72080 0 la_data_in[54]
rlabel metal2 307326 273751 307326 273751 0 la_data_in[55]
rlabel metal2 287730 67728 287730 67728 0 la_data_in[56]
rlabel metal1 272734 233818 272734 233818 0 la_data_in[57]
rlabel metal2 276230 232118 276230 232118 0 la_data_in[58]
rlabel metal2 335110 1758 335110 1758 0 la_data_in[59]
rlabel metal2 143566 78700 143566 78700 0 la_data_in[5]
rlabel metal1 308430 305014 308430 305014 0 la_data_in[60]
rlabel metal2 296286 269433 296286 269433 0 la_data_in[61]
rlabel metal2 345545 340 345545 340 0 la_data_in[62]
rlabel metal1 275080 229738 275080 229738 0 la_data_in[63]
rlabel metal2 293250 270198 293250 270198 0 la_data_in[64]
rlabel metal2 251114 145894 251114 145894 0 la_data_in[65]
rlabel metal2 309764 303076 309764 303076 0 la_data_in[66]
rlabel metal2 215970 76568 215970 76568 0 la_data_in[67]
rlabel metal2 367034 2132 367034 2132 0 la_data_in[68]
rlabel metal2 370385 340 370385 340 0 la_data_in[69]
rlabel metal2 292974 307734 292974 307734 0 la_data_in[6]
rlabel metal2 249734 134912 249734 134912 0 la_data_in[70]
rlabel metal1 311098 307666 311098 307666 0 la_data_in[71]
rlabel metal2 273286 143106 273286 143106 0 la_data_in[72]
rlabel metal2 384553 340 384553 340 0 la_data_in[73]
rlabel metal2 388049 340 388049 340 0 la_data_in[74]
rlabel metal2 252494 133552 252494 133552 0 la_data_in[75]
rlabel metal2 304566 270215 304566 270215 0 la_data_in[76]
rlabel metal1 351348 326366 351348 326366 0 la_data_in[77]
rlabel metal2 272366 155618 272366 155618 0 la_data_in[78]
rlabel metal2 288558 190536 288558 190536 0 la_data_in[79]
rlabel metal2 150558 16560 150558 16560 0 la_data_in[7]
rlabel metal2 409393 340 409393 340 0 la_data_in[80]
rlabel metal2 412889 340 412889 340 0 la_data_in[81]
rlabel metal2 416714 1928 416714 1928 0 la_data_in[82]
rlabel metal1 327382 309230 327382 309230 0 la_data_in[83]
rlabel metal2 423798 1928 423798 1928 0 la_data_in[84]
rlabel metal2 427057 340 427057 340 0 la_data_in[85]
rlabel metal2 430744 16560 430744 16560 0 la_data_in[86]
rlabel metal2 291134 156944 291134 156944 0 la_data_in[87]
rlabel metal2 289754 144568 289754 144568 0 la_data_in[88]
rlabel metal2 255898 136204 255898 136204 0 la_data_in[89]
rlabel metal2 154001 340 154001 340 0 la_data_in[8]
rlabel metal1 291778 231438 291778 231438 0 la_data_in[90]
rlabel metal2 448638 1928 448638 1928 0 la_data_in[91]
rlabel metal1 291640 231778 291640 231778 0 la_data_in[92]
rlabel metal1 287684 226338 287684 226338 0 la_data_in[93]
rlabel metal1 229494 140658 229494 140658 0 la_data_in[94]
rlabel metal2 462569 340 462569 340 0 la_data_in[95]
rlabel metal2 466111 340 466111 340 0 la_data_in[96]
rlabel metal2 469890 1928 469890 1928 0 la_data_in[97]
rlabel metal2 292606 125120 292606 125120 0 la_data_in[98]
rlabel metal2 476737 340 476737 340 0 la_data_in[99]
rlabel metal2 293986 307496 293986 307496 0 la_data_in[9]
rlabel metal2 127006 1826 127006 1826 0 la_data_out[0]
rlabel metal2 481758 3627 481758 3627 0 la_data_out[100]
rlabel metal2 485017 340 485017 340 0 la_data_out[101]
rlabel metal2 488704 16560 488704 16560 0 la_data_out[102]
rlabel metal1 406364 251226 406364 251226 0 la_data_out[103]
rlabel metal2 390678 351016 390678 351016 0 la_data_out[104]
rlabel metal2 268732 277380 268732 277380 0 la_data_out[105]
rlabel metal2 502688 16560 502688 16560 0 la_data_out[106]
rlabel metal2 506506 119602 506506 119602 0 la_data_out[107]
rlabel metal2 349922 347004 349922 347004 0 la_data_out[108]
rlabel metal1 334696 307666 334696 307666 0 la_data_out[109]
rlabel metal2 174846 130043 174846 130043 0 la_data_out[10]
rlabel metal1 322828 276046 322828 276046 0 la_data_out[110]
rlabel metal2 520529 340 520529 340 0 la_data_out[111]
rlabel metal2 524025 340 524025 340 0 la_data_out[112]
rlabel metal2 527850 3627 527850 3627 0 la_data_out[113]
rlabel metal2 327290 253164 327290 253164 0 la_data_out[114]
rlabel metal2 323058 249424 323058 249424 0 la_data_out[115]
rlabel metal2 538331 340 538331 340 0 la_data_out[116]
rlabel metal2 296378 232964 296378 232964 0 la_data_out[117]
rlabel metal2 545514 1724 545514 1724 0 la_data_out[118]
rlabel metal1 385480 327046 385480 327046 0 la_data_out[119]
rlabel metal2 292054 265761 292054 265761 0 la_data_out[11]
rlabel metal2 527896 16560 527896 16560 0 la_data_out[120]
rlabel metal1 222870 156910 222870 156910 0 la_data_out[121]
rlabel metal2 559537 340 559537 340 0 la_data_out[122]
rlabel metal2 563171 340 563171 340 0 la_data_out[123]
rlabel metal2 566858 1894 566858 1894 0 la_data_out[124]
rlabel metal2 386998 329443 386998 329443 0 la_data_out[125]
rlabel metal1 238050 177310 238050 177310 0 la_data_out[126]
rlabel metal2 577438 2234 577438 2234 0 la_data_out[127]
rlabel metal1 235198 227766 235198 227766 0 la_data_out[12]
rlabel metal2 172953 340 172953 340 0 la_data_out[13]
rlabel metal1 176318 23494 176318 23494 0 la_data_out[14]
rlabel metal2 180274 1911 180274 1911 0 la_data_out[15]
rlabel metal2 295366 303042 295366 303042 0 la_data_out[16]
rlabel metal3 177399 157828 177399 157828 0 la_data_out[17]
rlabel metal3 178825 136612 178825 136612 0 la_data_out[18]
rlabel metal2 194442 2030 194442 2030 0 la_data_out[19]
rlabel metal1 289846 305014 289846 305014 0 la_data_out[1]
rlabel metal3 177721 157420 177721 157420 0 la_data_out[20]
rlabel metal1 351164 387158 351164 387158 0 la_data_out[21]
rlabel metal3 178733 157420 178733 157420 0 la_data_out[22]
rlabel metal1 208932 153782 208932 153782 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215694 1826 215694 1826 0 la_data_out[25]
rlabel metal2 219282 1758 219282 1758 0 la_data_out[26]
rlabel metal2 289202 269382 289202 269382 0 la_data_out[27]
rlabel via3 180021 157420 180021 157420 0 la_data_out[28]
rlabel metal2 229625 340 229625 340 0 la_data_out[29]
rlabel metal2 134037 340 134037 340 0 la_data_out[2]
rlabel metal2 180550 159130 180550 159130 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal2 236716 151800 236716 151800 0 la_data_out[32]
rlabel metal2 345966 344692 345966 344692 0 la_data_out[33]
rlabel metal2 348542 346154 348542 346154 0 la_data_out[34]
rlabel metal2 251206 2200 251206 2200 0 la_data_out[35]
rlabel metal2 254702 2234 254702 2234 0 la_data_out[36]
rlabel metal2 182482 159300 182482 159300 0 la_data_out[37]
rlabel metal2 346242 348092 346242 348092 0 la_data_out[38]
rlabel metal2 183080 159732 183080 159732 0 la_data_out[39]
rlabel metal2 137441 340 137441 340 0 la_data_out[3]
rlabel metal2 268870 2030 268870 2030 0 la_data_out[40]
rlabel metal2 272182 16560 272182 16560 0 la_data_out[41]
rlabel metal2 276046 1996 276046 1996 0 la_data_out[42]
rlabel metal2 279305 340 279305 340 0 la_data_out[43]
rlabel metal2 268410 76330 268410 76330 0 la_data_out[44]
rlabel metal2 285706 234940 285706 234940 0 la_data_out[45]
rlabel metal2 290214 1928 290214 1928 0 la_data_out[46]
rlabel metal2 293710 1656 293710 1656 0 la_data_out[47]
rlabel metal1 301208 310386 301208 310386 0 la_data_out[48]
rlabel metal2 185794 158892 185794 158892 0 la_data_out[49]
rlabel metal2 141036 16560 141036 16560 0 la_data_out[4]
rlabel metal2 345874 342346 345874 342346 0 la_data_out[50]
rlabel metal2 307970 1911 307970 1911 0 la_data_out[51]
rlabel metal2 311466 1962 311466 1962 0 la_data_out[52]
rlabel metal2 315054 1690 315054 1690 0 la_data_out[53]
rlabel metal2 314042 3536 314042 3536 0 la_data_out[54]
rlabel metal2 307694 303433 307694 303433 0 la_data_out[55]
rlabel metal2 325634 2166 325634 2166 0 la_data_out[56]
rlabel metal1 307326 216546 307326 216546 0 la_data_out[57]
rlabel metal2 332718 551 332718 551 0 la_data_out[58]
rlabel metal1 292652 213214 292652 213214 0 la_data_out[59]
rlabel metal3 173213 147220 173213 147220 0 la_data_out[5]
rlabel metal2 237038 175950 237038 175950 0 la_data_out[60]
rlabel metal2 235842 173162 235842 173162 0 la_data_out[61]
rlabel metal1 311880 3298 311880 3298 0 la_data_out[62]
rlabel metal2 350474 1962 350474 1962 0 la_data_out[63]
rlabel metal2 353825 340 353825 340 0 la_data_out[64]
rlabel metal1 309856 291890 309856 291890 0 la_data_out[65]
rlabel metal2 309994 241995 309994 241995 0 la_data_out[66]
rlabel metal2 311558 245888 311558 245888 0 la_data_out[67]
rlabel metal2 367993 340 367993 340 0 la_data_out[68]
rlabel metal1 311098 311134 311098 311134 0 la_data_out[69]
rlabel metal2 148113 340 148113 340 0 la_data_out[6]
rlabel metal1 251850 223550 251850 223550 0 la_data_out[70]
rlabel metal1 311098 309026 311098 309026 0 la_data_out[71]
rlabel metal2 312892 248400 312892 248400 0 la_data_out[72]
rlabel metal1 251712 222122 251712 222122 0 la_data_out[73]
rlabel metal2 312478 250750 312478 250750 0 la_data_out[74]
rlabel metal2 392833 340 392833 340 0 la_data_out[75]
rlabel via3 253483 222156 253483 222156 0 la_data_out[76]
rlabel metal1 253138 222054 253138 222054 0 la_data_out[77]
rlabel metal2 372646 292162 372646 292162 0 la_data_out[78]
rlabel metal1 314410 249730 314410 249730 0 la_data_out[79]
rlabel metal2 151846 3627 151846 3627 0 la_data_out[7]
rlabel metal1 254610 221986 254610 221986 0 la_data_out[80]
rlabel metal2 255070 221646 255070 221646 0 la_data_out[81]
rlabel metal1 254610 222122 254610 222122 0 la_data_out[82]
rlabel metal1 254472 218926 254472 218926 0 la_data_out[83]
rlabel metal1 315836 251294 315836 251294 0 la_data_out[84]
rlabel metal2 251850 183243 251850 183243 0 la_data_out[85]
rlabel metal3 285913 257380 285913 257380 0 la_data_out[86]
rlabel metal1 256266 223346 256266 223346 0 la_data_out[87]
rlabel metal2 439024 16560 439024 16560 0 la_data_out[88]
rlabel metal2 442152 16560 442152 16560 0 la_data_out[89]
rlabel metal3 156446 153068 156446 153068 0 la_data_out[8]
rlabel metal2 446009 340 446009 340 0 la_data_out[90]
rlabel metal2 449834 1996 449834 1996 0 la_data_out[91]
rlabel metal2 257462 186728 257462 186728 0 la_data_out[92]
rlabel metal2 257370 184518 257370 184518 0 la_data_out[93]
rlabel metal2 460177 340 460177 340 0 la_data_out[94]
rlabel metal2 464002 1962 464002 1962 0 la_data_out[95]
rlabel metal2 466992 16560 466992 16560 0 la_data_out[96]
rlabel metal2 470849 340 470849 340 0 la_data_out[97]
rlabel metal2 474582 1962 474582 1962 0 la_data_out[98]
rlabel metal3 383640 314024 383640 314024 0 la_data_out[99]
rlabel metal2 293986 308584 293986 308584 0 la_data_out[9]
rlabel metal4 171764 138584 171764 138584 0 la_oenb[0]
rlabel metal2 482625 340 482625 340 0 la_oenb[100]
rlabel metal2 486128 16560 486128 16560 0 la_oenb[101]
rlabel metal2 489946 1843 489946 1843 0 la_oenb[102]
rlabel metal2 493297 340 493297 340 0 la_oenb[103]
rlabel metal3 231288 143276 231288 143276 0 la_oenb[104]
rlabel metal2 500112 16560 500112 16560 0 la_oenb[105]
rlabel metal2 503969 340 503969 340 0 la_oenb[106]
rlabel metal2 507465 340 507465 340 0 la_oenb[107]
rlabel metal3 322529 307564 322529 307564 0 la_oenb[108]
rlabel metal3 358685 101388 358685 101388 0 la_oenb[109]
rlabel metal2 163714 1792 163714 1792 0 la_oenb[10]
rlabel metal2 328486 267172 328486 267172 0 la_oenb[110]
rlabel metal2 521870 1928 521870 1928 0 la_oenb[111]
rlabel metal2 524952 16560 524952 16560 0 la_oenb[112]
rlabel metal2 528809 340 528809 340 0 la_oenb[113]
rlabel metal2 331246 323255 331246 323255 0 la_oenb[114]
rlabel metal2 330418 322371 330418 322371 0 la_oenb[115]
rlabel metal2 539626 3627 539626 3627 0 la_oenb[116]
rlabel metal2 542977 340 542977 340 0 la_oenb[117]
rlabel metal2 546611 340 546611 340 0 la_oenb[118]
rlabel metal1 385572 330514 385572 330514 0 la_oenb[119]
rlabel metal2 171442 3536 171442 3536 0 la_oenb[11]
rlabel metal3 353556 342924 353556 342924 0 la_oenb[120]
rlabel metal2 205804 155958 205804 155958 0 la_oenb[121]
rlabel metal2 560641 340 560641 340 0 la_oenb[122]
rlabel metal2 564466 42575 564466 42575 0 la_oenb[123]
rlabel metal2 567817 340 567817 340 0 la_oenb[124]
rlabel metal3 326669 310420 326669 310420 0 la_oenb[125]
rlabel metal3 237130 174556 237130 174556 0 la_oenb[126]
rlabel metal2 578450 16560 578450 16560 0 la_oenb[127]
rlabel metal3 174501 143412 174501 143412 0 la_oenb[12]
rlabel metal2 174103 340 174103 340 0 la_oenb[13]
rlabel metal1 177238 8262 177238 8262 0 la_oenb[14]
rlabel metal2 181233 340 181233 340 0 la_oenb[15]
rlabel metal2 184966 2064 184966 2064 0 la_oenb[16]
rlabel metal2 188140 16560 188140 16560 0 la_oenb[17]
rlabel metal2 192050 1928 192050 1928 0 la_oenb[18]
rlabel metal2 195401 340 195401 340 0 la_oenb[19]
rlabel metal2 131553 340 131553 340 0 la_oenb[1]
rlabel metal3 177583 157692 177583 157692 0 la_oenb[20]
rlabel metal3 178549 159868 178549 159868 0 la_oenb[21]
rlabel metal2 178434 158977 178434 158977 0 la_oenb[22]
rlabel metal3 178641 159732 178641 159732 0 la_oenb[23]
rlabel metal2 178986 158909 178986 158909 0 la_oenb[24]
rlabel metal2 179262 159385 179262 159385 0 la_oenb[25]
rlabel metal2 179538 158909 179538 158909 0 la_oenb[26]
rlabel metal2 179814 159385 179814 159385 0 la_oenb[27]
rlabel metal2 180090 159997 180090 159997 0 la_oenb[28]
rlabel metal3 180481 157420 180481 157420 0 la_oenb[29]
rlabel metal2 135286 1826 135286 1826 0 la_oenb[2]
rlabel metal2 180642 158977 180642 158977 0 la_oenb[30]
rlabel metal2 237905 340 237905 340 0 la_oenb[31]
rlabel metal3 181355 159868 181355 159868 0 la_oenb[32]
rlabel metal2 210910 275604 210910 275604 0 la_oenb[33]
rlabel metal2 248814 1724 248814 1724 0 la_oenb[34]
rlabel metal2 251850 16560 251850 16560 0 la_oenb[35]
rlabel metal2 255622 16560 255622 16560 0 la_oenb[36]
rlabel metal2 211094 234124 211094 234124 0 la_oenb[37]
rlabel metal2 262745 340 262745 340 0 la_oenb[38]
rlabel metal2 183126 159980 183126 159980 0 la_oenb[39]
rlabel metal2 138460 16560 138460 16560 0 la_oenb[3]
rlabel metal2 269606 16560 269606 16560 0 la_oenb[40]
rlabel metal1 211692 234158 211692 234158 0 la_oenb[41]
rlabel metal2 277150 1843 277150 1843 0 la_oenb[42]
rlabel metal2 184230 159929 184230 159929 0 la_oenb[43]
rlabel metal2 184506 159997 184506 159997 0 la_oenb[44]
rlabel metal2 287585 340 287585 340 0 la_oenb[45]
rlabel metal2 195454 140012 195454 140012 0 la_oenb[46]
rlabel metal2 294906 3475 294906 3475 0 la_oenb[47]
rlabel metal2 298303 340 298303 340 0 la_oenb[48]
rlabel metal2 185886 159436 185886 159436 0 la_oenb[49]
rlabel metal4 292652 268812 292652 268812 0 la_oenb[4]
rlabel metal1 246744 218110 246744 218110 0 la_oenb[50]
rlabel metal3 195316 140352 195316 140352 0 la_oenb[51]
rlabel metal2 312662 1928 312662 1928 0 la_oenb[52]
rlabel metal2 315422 13430 315422 13430 0 la_oenb[53]
rlabel metal3 306912 302260 306912 302260 0 la_oenb[54]
rlabel metal2 238050 182903 238050 182903 0 la_oenb[55]
rlabel metal2 326830 2200 326830 2200 0 la_oenb[56]
rlabel metal2 330418 2574 330418 2574 0 la_oenb[57]
rlabel metal2 333914 1860 333914 1860 0 la_oenb[58]
rlabel metal4 249780 222088 249780 222088 0 la_oenb[59]
rlabel metal2 145721 340 145721 340 0 la_oenb[5]
rlabel via2 309074 297653 309074 297653 0 la_oenb[60]
rlabel metal3 249228 220864 249228 220864 0 la_oenb[61]
rlabel metal2 347944 16560 347944 16560 0 la_oenb[62]
rlabel metal2 351433 340 351433 340 0 la_oenb[63]
rlabel metal4 309212 252964 309212 252964 0 la_oenb[64]
rlabel metal3 206747 141236 206747 141236 0 la_oenb[65]
rlabel metal2 230230 166226 230230 166226 0 la_oenb[66]
rlabel metal2 365838 3407 365838 3407 0 la_oenb[67]
rlabel metal2 369426 3322 369426 3322 0 la_oenb[68]
rlabel metal3 191383 140828 191383 140828 0 la_oenb[69]
rlabel metal2 153870 75582 153870 75582 0 la_oenb[6]
rlabel metal2 235382 180948 235382 180948 0 la_oenb[70]
rlabel metal4 251804 178492 251804 178492 0 la_oenb[71]
rlabel metal1 312846 300730 312846 300730 0 la_oenb[72]
rlabel metal2 387182 4835 387182 4835 0 la_oenb[73]
rlabel metal2 390678 3271 390678 3271 0 la_oenb[74]
rlabel metal3 221444 137428 221444 137428 0 la_oenb[75]
rlabel metal2 253690 160205 253690 160205 0 la_oenb[76]
rlabel metal3 194143 209508 194143 209508 0 la_oenb[77]
rlabel metal2 404609 340 404609 340 0 la_oenb[78]
rlabel metal2 408434 1860 408434 1860 0 la_oenb[79]
rlabel metal2 153042 4988 153042 4988 0 la_oenb[7]
rlabel metal3 314180 299404 314180 299404 0 la_oenb[80]
rlabel metal2 373934 349860 373934 349860 0 la_oenb[81]
rlabel metal1 274942 219130 274942 219130 0 la_oenb[82]
rlabel metal3 195707 209508 195707 209508 0 la_oenb[83]
rlabel metal1 256404 173978 256404 173978 0 la_oenb[84]
rlabel metal2 429449 340 429449 340 0 la_oenb[85]
rlabel metal2 256174 162061 256174 162061 0 la_oenb[86]
rlabel metal2 436770 1707 436770 1707 0 la_oenb[87]
rlabel metal3 318757 11628 318757 11628 0 la_oenb[88]
rlabel metal2 443617 340 443617 340 0 la_oenb[89]
rlabel metal2 156393 340 156393 340 0 la_oenb[8]
rlabel metal2 257646 159239 257646 159239 0 la_oenb[90]
rlabel metal2 450432 16560 450432 16560 0 la_oenb[91]
rlabel metal2 257554 216104 257554 216104 0 la_oenb[92]
rlabel metal2 458114 1928 458114 1928 0 la_oenb[93]
rlabel metal2 198674 140165 198674 140165 0 la_oenb[94]
rlabel metal2 465198 6722 465198 6722 0 la_oenb[95]
rlabel metal2 468457 340 468457 340 0 la_oenb[96]
rlabel metal2 319194 386895 319194 386895 0 la_oenb[97]
rlabel metal2 346334 326196 346334 326196 0 la_oenb[98]
rlabel metal2 479129 340 479129 340 0 la_oenb[99]
rlabel metal2 160126 3627 160126 3627 0 la_oenb[9]
rlabel metal2 1702 1962 1702 1962 0 wb_rst_i
rlabel metal2 2898 1894 2898 1894 0 wbs_ack_o
rlabel metal2 155434 190383 155434 190383 0 wbs_adr_i[0]
rlabel metal2 155802 194582 155802 194582 0 wbs_adr_i[10]
rlabel metal2 156722 154700 156722 154700 0 wbs_adr_i[11]
rlabel metal1 109756 97342 109756 97342 0 wbs_adr_i[12]
rlabel metal2 58236 16560 58236 16560 0 wbs_adr_i[13]
rlabel metal2 61863 340 61863 340 0 wbs_adr_i[14]
rlabel metal2 155526 187000 155526 187000 0 wbs_adr_i[15]
rlabel metal2 156952 166260 156952 166260 0 wbs_adr_i[16]
rlabel metal2 270434 308822 270434 308822 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 152950 156264 152950 156264 0 wbs_adr_i[1]
rlabel metal2 152904 159766 152904 159766 0 wbs_adr_i[20]
rlabel metal2 154514 193528 154514 193528 0 wbs_adr_i[21]
rlabel metal2 153134 190859 153134 190859 0 wbs_adr_i[22]
rlabel metal2 93932 16560 93932 16560 0 wbs_adr_i[23]
rlabel metal2 153042 159460 153042 159460 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal1 156952 166158 156952 166158 0 wbs_adr_i[26]
rlabel metal3 293020 299132 293020 299132 0 wbs_adr_i[27]
rlabel metal2 111642 1962 111642 1962 0 wbs_adr_i[28]
rlabel metal2 115230 1622 115230 1622 0 wbs_adr_i[29]
rlabel metal2 16836 16560 16836 16560 0 wbs_adr_i[2]
rlabel metal2 118818 2030 118818 2030 0 wbs_adr_i[30]
rlabel metal2 172454 141100 172454 141100 0 wbs_adr_i[31]
rlabel metal2 21298 16560 21298 16560 0 wbs_adr_i[3]
rlabel metal2 269882 353617 269882 353617 0 wbs_adr_i[4]
rlabel metal2 212198 278052 212198 278052 0 wbs_adr_i[5]
rlabel metal2 157274 199427 157274 199427 0 wbs_adr_i[6]
rlabel metal2 37023 340 37023 340 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 44298 2098 44298 2098 0 wbs_adr_i[9]
rlabel metal2 4094 1928 4094 1928 0 wbs_cyc_i
rlabel metal1 86020 133178 86020 133178 0 wbs_dat_i[0]
rlabel metal2 212474 277712 212474 277712 0 wbs_dat_i[10]
rlabel via3 166221 137564 166221 137564 0 wbs_dat_i[11]
rlabel metal2 55660 16560 55660 16560 0 wbs_dat_i[12]
rlabel metal2 59517 340 59517 340 0 wbs_dat_i[13]
rlabel metal2 62698 16560 62698 16560 0 wbs_dat_i[14]
rlabel metal1 287730 301546 287730 301546 0 wbs_dat_i[15]
rlabel metal3 292675 299268 292675 299268 0 wbs_dat_i[16]
rlabel metal2 75210 21012 75210 21012 0 wbs_dat_i[17]
rlabel metal2 77418 1826 77418 1826 0 wbs_dat_i[18]
rlabel metal2 231334 294508 231334 294508 0 wbs_dat_i[19]
rlabel metal2 13570 1962 13570 1962 0 wbs_dat_i[1]
rlabel metal2 288650 295069 288650 295069 0 wbs_dat_i[20]
rlabel metal2 87761 340 87761 340 0 wbs_dat_i[21]
rlabel metal2 91356 16560 91356 16560 0 wbs_dat_i[22]
rlabel metal2 95174 1962 95174 1962 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102258 3627 102258 3627 0 wbs_dat_i[25]
rlabel metal2 105340 16560 105340 16560 0 wbs_dat_i[26]
rlabel metal2 109342 1860 109342 1860 0 wbs_dat_i[27]
rlabel metal2 112601 340 112601 340 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18262 1826 18262 1826 0 wbs_dat_i[2]
rlabel metal2 119922 1962 119922 1962 0 wbs_dat_i[30]
rlabel metal2 123273 340 123273 340 0 wbs_dat_i[31]
rlabel metal2 22809 340 22809 340 0 wbs_dat_i[3]
rlabel metal2 27738 1792 27738 1792 0 wbs_dat_i[4]
rlabel metal2 153962 186286 153962 186286 0 wbs_dat_i[5]
rlabel metal1 269238 317390 269238 317390 0 wbs_dat_i[6]
rlabel metal2 38410 1928 38410 1928 0 wbs_dat_i[7]
rlabel metal2 41906 1690 41906 1690 0 wbs_dat_i[8]
rlabel metal2 45303 340 45303 340 0 wbs_dat_i[9]
rlabel metal2 9837 340 9837 340 0 wbs_dat_o[0]
rlabel metal2 166198 156876 166198 156876 0 wbs_dat_o[10]
rlabel metal2 53774 1928 53774 1928 0 wbs_dat_o[11]
rlabel metal2 57033 340 57033 340 0 wbs_dat_o[12]
rlabel metal2 288374 296429 288374 296429 0 wbs_dat_o[13]
rlabel metal2 63940 16560 63940 16560 0 wbs_dat_o[14]
rlabel metal2 257186 309944 257186 309944 0 wbs_dat_o[15]
rlabel metal2 71530 1911 71530 1911 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78614 3968 78614 3968 0 wbs_dat_o[18]
rlabel metal2 81873 340 81873 340 0 wbs_dat_o[19]
rlabel metal2 25530 66334 25530 66334 0 wbs_dat_o[1]
rlabel metal1 289018 311270 289018 311270 0 wbs_dat_o[20]
rlabel metal2 89194 1911 89194 1911 0 wbs_dat_o[21]
rlabel metal2 211094 237796 211094 237796 0 wbs_dat_o[22]
rlabel metal2 96278 1996 96278 1996 0 wbs_dat_o[23]
rlabel metal2 290536 311236 290536 311236 0 wbs_dat_o[24]
rlabel metal2 102810 16560 102810 16560 0 wbs_dat_o[25]
rlabel metal2 106713 340 106713 340 0 wbs_dat_o[26]
rlabel metal2 290996 306360 290996 306360 0 wbs_dat_o[27]
rlabel metal2 114034 1962 114034 1962 0 wbs_dat_o[28]
rlabel metal2 117477 340 117477 340 0 wbs_dat_o[29]
rlabel metal2 19458 2574 19458 2574 0 wbs_dat_o[2]
rlabel metal2 120881 340 120881 340 0 wbs_dat_o[30]
rlabel metal2 160770 80342 160770 80342 0 wbs_dat_o[31]
rlabel metal2 23874 16560 23874 16560 0 wbs_dat_o[3]
rlabel metal2 28697 340 28697 340 0 wbs_dat_o[4]
rlabel metal2 32193 340 32193 340 0 wbs_dat_o[5]
rlabel metal2 36018 5328 36018 5328 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 42957 340 42957 340 0 wbs_dat_o[8]
rlabel metal2 335202 337569 335202 337569 0 wbs_dat_o[9]
rlabel metal2 253782 317849 253782 317849 0 wbs_sel_i[0]
rlabel metal2 192510 235433 192510 235433 0 wbs_sel_i[1]
rlabel metal2 20417 340 20417 340 0 wbs_sel_i[2]
rlabel metal2 25346 6722 25346 6722 0 wbs_sel_i[3]
rlabel metal2 191682 235484 191682 235484 0 wbs_stb_i
rlabel metal2 6486 1996 6486 1996 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
