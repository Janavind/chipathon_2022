magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 67 641 203
rect 30 21 641 67
rect 30 -17 64 21
<< scnmos >>
rect 79 93 109 177
rect 281 47 311 177
rect 365 47 395 177
rect 449 47 479 177
rect 533 47 563 177
<< scpmoshvt >>
rect 79 297 109 381
rect 177 297 207 497
rect 273 297 303 497
rect 437 297 467 497
rect 521 297 551 497
<< ndiff >>
rect 27 152 79 177
rect 27 118 35 152
rect 69 118 79 152
rect 27 93 79 118
rect 109 161 174 177
rect 109 127 119 161
rect 153 127 174 161
rect 109 93 174 127
rect 124 59 132 93
rect 166 59 174 93
rect 124 47 174 59
rect 229 161 281 177
rect 229 127 237 161
rect 271 127 281 161
rect 229 93 281 127
rect 229 59 237 93
rect 271 59 281 93
rect 229 47 281 59
rect 311 161 365 177
rect 311 127 321 161
rect 355 127 365 161
rect 311 47 365 127
rect 395 161 449 177
rect 395 127 405 161
rect 439 127 449 161
rect 395 93 449 127
rect 395 59 405 93
rect 439 59 449 93
rect 395 47 449 59
rect 479 89 533 177
rect 479 55 489 89
rect 523 55 533 89
rect 479 47 533 55
rect 563 161 615 177
rect 563 127 573 161
rect 607 127 615 161
rect 563 93 615 127
rect 563 59 573 93
rect 607 59 615 93
rect 563 47 615 59
<< pdiff >>
rect 125 485 177 497
rect 125 451 133 485
rect 167 451 177 485
rect 125 417 177 451
rect 125 383 133 417
rect 167 383 177 417
rect 125 381 177 383
rect 27 356 79 381
rect 27 322 35 356
rect 69 322 79 356
rect 27 297 79 322
rect 109 297 177 381
rect 207 485 273 497
rect 207 451 223 485
rect 257 451 273 485
rect 207 417 273 451
rect 207 383 223 417
rect 257 383 273 417
rect 207 297 273 383
rect 303 485 437 497
rect 303 451 313 485
rect 347 451 381 485
rect 415 451 437 485
rect 303 297 437 451
rect 467 485 521 497
rect 467 451 477 485
rect 511 451 521 485
rect 467 417 521 451
rect 467 383 477 417
rect 511 383 521 417
rect 467 349 521 383
rect 467 315 477 349
rect 511 315 521 349
rect 467 297 521 315
rect 551 485 606 497
rect 551 451 561 485
rect 595 451 606 485
rect 551 417 606 451
rect 551 383 561 417
rect 595 383 606 417
rect 551 349 606 383
rect 551 315 561 349
rect 595 315 606 349
rect 551 297 606 315
<< ndiffc >>
rect 35 118 69 152
rect 119 127 153 161
rect 132 59 166 93
rect 237 127 271 161
rect 237 59 271 93
rect 321 127 355 161
rect 405 127 439 161
rect 405 59 439 93
rect 489 55 523 89
rect 573 127 607 161
rect 573 59 607 93
<< pdiffc >>
rect 133 451 167 485
rect 133 383 167 417
rect 35 322 69 356
rect 223 451 257 485
rect 223 383 257 417
rect 313 451 347 485
rect 381 451 415 485
rect 477 451 511 485
rect 477 383 511 417
rect 477 315 511 349
rect 561 451 595 485
rect 561 383 595 417
rect 561 315 595 349
<< poly >>
rect 177 497 207 523
rect 273 497 303 523
rect 437 497 467 523
rect 521 497 551 523
rect 79 381 109 407
rect 79 265 109 297
rect 79 249 135 265
rect 79 215 91 249
rect 125 215 135 249
rect 79 199 135 215
rect 177 259 207 297
rect 273 259 303 297
rect 437 259 467 297
rect 521 261 551 297
rect 521 259 623 261
rect 177 249 395 259
rect 177 215 222 249
rect 256 215 395 249
rect 177 205 395 215
rect 437 249 623 259
rect 437 215 477 249
rect 511 215 573 249
rect 607 215 623 249
rect 437 205 623 215
rect 79 177 109 199
rect 281 177 311 205
rect 365 177 395 205
rect 449 177 479 205
rect 533 203 623 205
rect 533 177 563 203
rect 79 67 109 93
rect 281 21 311 47
rect 365 21 395 47
rect 449 21 479 47
rect 533 21 563 47
<< polycont >>
rect 91 215 125 249
rect 222 215 256 249
rect 477 215 511 249
rect 573 215 607 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 116 485 167 527
rect 116 451 133 485
rect 116 417 167 451
rect 116 383 133 417
rect 22 356 82 372
rect 116 367 167 383
rect 207 485 273 493
rect 207 451 223 485
rect 257 451 273 485
rect 207 417 273 451
rect 307 485 422 527
rect 307 451 313 485
rect 347 451 381 485
rect 415 451 422 485
rect 307 435 422 451
rect 456 485 527 493
rect 456 451 477 485
rect 511 451 527 485
rect 207 383 223 417
rect 257 401 273 417
rect 456 417 527 451
rect 456 401 477 417
rect 257 383 477 401
rect 511 383 527 417
rect 207 367 527 383
rect 22 322 35 356
rect 69 333 82 356
rect 69 322 272 333
rect 22 299 272 322
rect 22 168 56 299
rect 91 249 160 265
rect 125 215 160 249
rect 206 249 272 299
rect 206 215 222 249
rect 256 215 272 249
rect 91 199 160 215
rect 306 181 362 367
rect 472 349 527 367
rect 398 255 436 331
rect 472 315 477 349
rect 511 315 527 349
rect 472 299 527 315
rect 561 485 627 527
rect 595 451 627 485
rect 561 417 627 451
rect 595 383 627 417
rect 561 349 627 383
rect 595 315 627 349
rect 561 299 627 315
rect 398 249 627 255
rect 398 215 477 249
rect 511 215 573 249
rect 607 215 627 249
rect 22 152 69 168
rect 22 118 35 152
rect 22 102 69 118
rect 103 161 169 165
rect 103 127 119 161
rect 153 127 169 161
rect 103 93 169 127
rect 103 59 132 93
rect 166 59 169 93
rect 103 17 169 59
rect 216 161 271 181
rect 306 161 371 181
rect 216 127 237 161
rect 305 127 321 161
rect 355 127 371 161
rect 405 161 627 181
rect 439 139 573 161
rect 439 127 455 139
rect 216 93 271 127
rect 405 93 455 127
rect 557 127 573 139
rect 607 127 627 161
rect 216 59 237 93
rect 271 59 405 93
rect 439 59 455 93
rect 216 51 455 59
rect 489 89 523 105
rect 489 17 523 55
rect 557 93 627 127
rect 557 59 573 93
rect 607 59 627 93
rect 557 51 627 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 582 221 616 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 311 153 345 187 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 306 289 340 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 306 357 340 391 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand2b_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1811168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1804606
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
