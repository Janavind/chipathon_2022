magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 1 21 355 203
rect 30 -17 64 21
<< locali >>
rect 18 456 234 490
rect 18 299 85 456
rect 119 265 166 401
rect 200 333 234 456
rect 200 299 263 333
rect 18 199 85 265
rect 119 199 195 265
rect 229 165 263 299
rect 18 131 263 165
rect 297 131 351 333
rect 18 77 69 131
rect 203 77 237 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 287 367 350 527
rect 103 17 169 97
rect 271 17 337 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 297 131 351 333 6 A
port 1 nsew signal input
rlabel locali s 119 199 195 265 6 B
port 2 nsew signal input
rlabel locali s 119 265 166 401 6 B
port 2 nsew signal input
rlabel locali s 18 199 85 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 355 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 203 77 237 131 6 Y
port 8 nsew signal output
rlabel locali s 18 77 69 131 6 Y
port 8 nsew signal output
rlabel locali s 18 131 263 165 6 Y
port 8 nsew signal output
rlabel locali s 229 165 263 299 6 Y
port 8 nsew signal output
rlabel locali s 200 299 263 333 6 Y
port 8 nsew signal output
rlabel locali s 200 333 234 456 6 Y
port 8 nsew signal output
rlabel locali s 18 299 85 456 6 Y
port 8 nsew signal output
rlabel locali s 18 456 234 490 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2004092
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1999912
<< end >>
