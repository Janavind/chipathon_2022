magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1195 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 530 47 560 177
rect 614 47 644 177
rect 700 47 730 177
rect 784 47 814 177
rect 983 47 1013 177
rect 1087 47 1117 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 596 297 626 497
rect 686 297 716 497
rect 838 297 868 497
rect 923 297 953 497
rect 1087 297 1117 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 247 177
rect 193 127 203 161
rect 237 127 247 161
rect 193 93 247 127
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 47 331 131
rect 361 93 413 177
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 478 93 530 177
rect 478 59 486 93
rect 520 59 530 93
rect 478 47 530 59
rect 560 165 614 177
rect 560 131 570 165
rect 604 131 614 165
rect 560 47 614 131
rect 644 93 700 177
rect 644 59 656 93
rect 690 59 700 93
rect 644 47 700 59
rect 730 161 784 177
rect 730 127 740 161
rect 774 127 784 161
rect 730 47 784 127
rect 814 93 866 177
rect 814 59 824 93
rect 858 59 866 93
rect 814 47 866 59
rect 920 93 983 177
rect 920 59 928 93
rect 962 59 983 93
rect 920 47 983 59
rect 1013 161 1087 177
rect 1013 127 1028 161
rect 1062 127 1087 161
rect 1013 89 1087 127
rect 1013 55 1028 89
rect 1062 55 1087 89
rect 1013 47 1087 55
rect 1117 161 1169 177
rect 1117 127 1127 161
rect 1161 127 1169 161
rect 1117 93 1169 127
rect 1117 59 1127 93
rect 1161 59 1169 93
rect 1117 47 1169 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 425 163 497
rect 109 391 119 425
rect 153 391 163 425
rect 109 357 163 391
rect 109 323 119 357
rect 153 323 163 357
rect 109 297 163 323
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 409 331 497
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 485 596 497
rect 445 451 470 485
rect 504 451 538 485
rect 572 451 596 485
rect 445 297 596 451
rect 626 477 686 497
rect 626 443 636 477
rect 670 443 686 477
rect 626 409 686 443
rect 626 375 636 409
rect 670 375 686 409
rect 626 297 686 375
rect 716 485 838 497
rect 716 451 726 485
rect 760 451 794 485
rect 828 451 838 485
rect 716 297 838 451
rect 868 477 923 497
rect 868 443 878 477
rect 912 443 923 477
rect 868 409 923 443
rect 868 375 878 409
rect 912 375 923 409
rect 868 297 923 375
rect 953 485 1087 497
rect 953 451 969 485
rect 1003 451 1037 485
rect 1071 451 1087 485
rect 953 297 1087 451
rect 1117 477 1169 497
rect 1117 443 1127 477
rect 1161 443 1169 477
rect 1117 409 1169 443
rect 1117 375 1127 409
rect 1161 375 1169 409
rect 1117 297 1169 375
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 203 127 237 161
rect 203 59 237 93
rect 287 131 321 165
rect 371 59 405 93
rect 486 59 520 93
rect 570 131 604 165
rect 656 59 690 93
rect 740 127 774 161
rect 824 59 858 93
rect 928 59 962 93
rect 1028 127 1062 161
rect 1028 55 1062 89
rect 1127 127 1161 161
rect 1127 59 1161 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 391 153 425
rect 119 323 153 357
rect 203 443 237 477
rect 203 375 237 409
rect 287 375 321 409
rect 371 443 405 477
rect 371 375 405 409
rect 470 451 504 485
rect 538 451 572 485
rect 636 443 670 477
rect 636 375 670 409
rect 726 451 760 485
rect 794 451 828 485
rect 878 443 912 477
rect 878 375 912 409
rect 969 451 1003 485
rect 1037 451 1071 485
rect 1127 443 1161 477
rect 1127 375 1161 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 596 497 626 523
rect 686 497 716 523
rect 838 497 868 523
rect 923 497 953 523
rect 1087 497 1117 523
rect 79 265 109 297
rect 163 265 193 297
rect 31 249 193 265
rect 247 259 277 297
rect 331 259 361 297
rect 31 215 47 249
rect 81 215 115 249
rect 149 215 193 249
rect 31 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 235 249 361 259
rect 235 215 251 249
rect 285 215 361 249
rect 235 195 361 215
rect 415 259 445 297
rect 596 259 626 297
rect 686 259 716 297
rect 838 259 868 297
rect 923 259 953 297
rect 1087 261 1117 297
rect 1087 259 1172 261
rect 415 249 644 259
rect 415 215 526 249
rect 560 215 594 249
rect 628 215 644 249
rect 415 205 644 215
rect 686 249 879 259
rect 686 215 761 249
rect 795 215 829 249
rect 863 215 879 249
rect 686 207 879 215
rect 247 177 277 195
rect 331 177 361 195
rect 530 177 560 205
rect 614 177 644 205
rect 700 205 879 207
rect 923 249 1172 259
rect 923 215 986 249
rect 1020 215 1054 249
rect 1088 215 1122 249
rect 1156 215 1172 249
rect 923 205 1172 215
rect 700 177 730 205
rect 784 177 814 205
rect 983 177 1013 205
rect 1087 203 1172 205
rect 1087 177 1117 203
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 530 21 560 47
rect 614 21 644 47
rect 700 21 730 47
rect 784 21 814 47
rect 983 21 1013 47
rect 1087 21 1117 47
<< polycont >>
rect 47 215 81 249
rect 115 215 149 249
rect 251 215 285 249
rect 526 215 560 249
rect 594 215 628 249
rect 761 215 795 249
rect 829 215 863 249
rect 986 215 1020 249
rect 1054 215 1088 249
rect 1122 215 1156 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 35 477 405 493
rect 69 459 203 477
rect 35 409 69 443
rect 237 459 371 477
rect 103 391 119 425
rect 153 391 169 425
rect 203 409 237 443
rect 454 485 588 527
rect 454 451 470 485
rect 504 451 538 485
rect 572 451 588 485
rect 636 477 670 493
rect 35 359 69 375
rect 119 357 153 391
rect 203 359 237 375
rect 287 409 321 425
rect 29 257 65 325
rect 287 325 321 375
rect 371 417 405 443
rect 710 485 844 527
rect 710 451 726 485
rect 760 451 794 485
rect 828 451 844 485
rect 878 477 912 493
rect 636 417 670 443
rect 953 485 1087 527
rect 953 451 969 485
rect 1003 451 1037 485
rect 1071 451 1087 485
rect 1127 477 1161 493
rect 878 417 912 443
rect 1127 417 1161 443
rect 371 409 1161 417
rect 405 383 636 409
rect 371 359 405 375
rect 670 383 878 409
rect 636 359 670 375
rect 912 383 1127 409
rect 878 359 912 375
rect 1127 359 1161 375
rect 153 323 436 325
rect 119 291 436 323
rect 29 249 165 257
rect 29 215 47 249
rect 81 215 115 249
rect 149 215 165 249
rect 209 249 345 257
rect 209 216 251 249
rect 235 215 251 216
rect 285 216 345 249
rect 285 215 301 216
rect 35 161 237 177
rect 393 165 436 291
rect 483 249 644 325
rect 483 215 526 249
rect 560 215 594 249
rect 628 215 644 249
rect 745 249 896 325
rect 745 215 761 249
rect 795 215 829 249
rect 863 215 896 249
rect 943 249 1172 325
rect 943 215 986 249
rect 1020 215 1054 249
rect 1088 215 1122 249
rect 1156 215 1172 249
rect 69 143 203 161
rect 35 93 69 127
rect 271 131 287 165
rect 321 131 570 165
rect 604 131 620 165
rect 1112 161 1177 177
rect 724 127 740 161
rect 774 127 1028 161
rect 1062 127 1078 161
rect 119 93 153 109
rect 203 93 237 127
rect 19 59 35 93
rect 69 59 85 93
rect 187 59 203 93
rect 237 59 371 93
rect 405 59 423 93
rect 470 59 486 93
rect 520 59 656 93
rect 690 59 824 93
rect 858 59 874 93
rect 911 59 928 93
rect 962 59 978 93
rect 119 17 153 59
rect 911 17 978 59
rect 1012 89 1078 127
rect 1012 55 1028 89
rect 1062 55 1078 89
rect 1112 127 1127 161
rect 1161 127 1177 161
rect 1112 93 1177 127
rect 1112 59 1127 93
rect 1161 59 1177 93
rect 1112 17 1177 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 950 289 984 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1042 289 1076 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1134 221 1168 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1134 289 1168 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 858 289 892 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 766 289 800 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 582 289 616 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 490 289 524 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 398 153 432 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a32oi_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 3504422
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3493188
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
