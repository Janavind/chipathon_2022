magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect 0 1464 978 2596
<< pwell >>
rect 20 606 1032 1386
rect 20 400 110 606
rect 20 83 1090 400
rect 20 10 110 83
<< mvnmos >>
rect 211 1060 311 1360
rect 353 1060 553 1360
rect 609 1060 809 1360
rect 853 1060 953 1360
rect 211 632 311 932
rect 353 632 553 932
rect 609 632 809 932
rect 853 632 953 932
rect 211 290 1011 374
rect 211 109 1011 193
<< mvpmos >>
rect 211 1530 331 2530
rect 387 1530 507 2530
rect 563 1530 683 2530
rect 739 1530 859 2530
<< mvndiff >>
rect 158 1348 211 1360
rect 158 1314 166 1348
rect 200 1314 211 1348
rect 158 1280 211 1314
rect 158 1246 166 1280
rect 200 1246 211 1280
rect 158 1212 211 1246
rect 158 1178 166 1212
rect 200 1178 211 1212
rect 158 1144 211 1178
rect 158 1110 166 1144
rect 200 1110 211 1144
rect 158 1060 211 1110
rect 311 1060 353 1360
rect 553 1348 609 1360
rect 553 1314 564 1348
rect 598 1314 609 1348
rect 553 1280 609 1314
rect 553 1246 564 1280
rect 598 1246 609 1280
rect 553 1212 609 1246
rect 553 1178 564 1212
rect 598 1178 609 1212
rect 553 1144 609 1178
rect 553 1110 564 1144
rect 598 1110 609 1144
rect 553 1060 609 1110
rect 809 1060 853 1360
rect 953 1348 1006 1360
rect 953 1314 964 1348
rect 998 1314 1006 1348
rect 953 1280 1006 1314
rect 953 1246 964 1280
rect 998 1246 1006 1280
rect 953 1212 1006 1246
rect 953 1178 964 1212
rect 998 1178 1006 1212
rect 953 1144 1006 1178
rect 953 1110 964 1144
rect 998 1110 1006 1144
rect 953 1060 1006 1110
rect 158 882 211 932
rect 158 848 166 882
rect 200 848 211 882
rect 158 814 211 848
rect 158 780 166 814
rect 200 780 211 814
rect 158 746 211 780
rect 158 712 166 746
rect 200 712 211 746
rect 158 678 211 712
rect 158 644 166 678
rect 200 644 211 678
rect 158 632 211 644
rect 311 632 353 932
rect 553 882 609 932
rect 553 848 564 882
rect 598 848 609 882
rect 553 814 609 848
rect 553 780 564 814
rect 598 780 609 814
rect 553 746 609 780
rect 553 712 564 746
rect 598 712 609 746
rect 553 678 609 712
rect 553 644 564 678
rect 598 644 609 678
rect 553 632 609 644
rect 809 632 853 932
rect 953 882 1006 932
rect 953 848 964 882
rect 998 848 1006 882
rect 953 814 1006 848
rect 953 780 964 814
rect 998 780 1006 814
rect 953 746 1006 780
rect 953 712 964 746
rect 998 712 1006 746
rect 953 678 1006 712
rect 953 644 964 678
rect 998 644 1006 678
rect 953 632 1006 644
rect 158 336 211 374
rect 158 302 166 336
rect 200 302 211 336
rect 158 290 211 302
rect 1011 336 1064 374
rect 1011 302 1022 336
rect 1056 302 1064 336
rect 1011 290 1064 302
rect 158 181 211 193
rect 158 147 166 181
rect 200 147 211 181
rect 158 109 211 147
rect 1011 181 1064 193
rect 1011 147 1022 181
rect 1056 147 1064 181
rect 1011 109 1064 147
<< mvpdiff >>
rect 158 2460 211 2530
rect 158 2426 166 2460
rect 200 2426 211 2460
rect 158 2392 211 2426
rect 158 2358 166 2392
rect 200 2358 211 2392
rect 158 2324 211 2358
rect 158 2290 166 2324
rect 200 2290 211 2324
rect 158 2256 211 2290
rect 158 2222 166 2256
rect 200 2222 211 2256
rect 158 2188 211 2222
rect 158 2154 166 2188
rect 200 2154 211 2188
rect 158 2120 211 2154
rect 158 2086 166 2120
rect 200 2086 211 2120
rect 158 2052 211 2086
rect 158 2018 166 2052
rect 200 2018 211 2052
rect 158 1984 211 2018
rect 158 1950 166 1984
rect 200 1950 211 1984
rect 158 1916 211 1950
rect 158 1882 166 1916
rect 200 1882 211 1916
rect 158 1848 211 1882
rect 158 1814 166 1848
rect 200 1814 211 1848
rect 158 1780 211 1814
rect 158 1746 166 1780
rect 200 1746 211 1780
rect 158 1712 211 1746
rect 158 1678 166 1712
rect 200 1678 211 1712
rect 158 1644 211 1678
rect 158 1610 166 1644
rect 200 1610 211 1644
rect 158 1576 211 1610
rect 158 1542 166 1576
rect 200 1542 211 1576
rect 158 1530 211 1542
rect 331 2460 387 2530
rect 331 2426 342 2460
rect 376 2426 387 2460
rect 331 2392 387 2426
rect 331 2358 342 2392
rect 376 2358 387 2392
rect 331 2324 387 2358
rect 331 2290 342 2324
rect 376 2290 387 2324
rect 331 2256 387 2290
rect 331 2222 342 2256
rect 376 2222 387 2256
rect 331 2188 387 2222
rect 331 2154 342 2188
rect 376 2154 387 2188
rect 331 2120 387 2154
rect 331 2086 342 2120
rect 376 2086 387 2120
rect 331 2052 387 2086
rect 331 2018 342 2052
rect 376 2018 387 2052
rect 331 1984 387 2018
rect 331 1950 342 1984
rect 376 1950 387 1984
rect 331 1916 387 1950
rect 331 1882 342 1916
rect 376 1882 387 1916
rect 331 1848 387 1882
rect 331 1814 342 1848
rect 376 1814 387 1848
rect 331 1780 387 1814
rect 331 1746 342 1780
rect 376 1746 387 1780
rect 331 1712 387 1746
rect 331 1678 342 1712
rect 376 1678 387 1712
rect 331 1644 387 1678
rect 331 1610 342 1644
rect 376 1610 387 1644
rect 331 1576 387 1610
rect 331 1542 342 1576
rect 376 1542 387 1576
rect 331 1530 387 1542
rect 507 2460 563 2530
rect 507 2426 518 2460
rect 552 2426 563 2460
rect 507 2392 563 2426
rect 507 2358 518 2392
rect 552 2358 563 2392
rect 507 2324 563 2358
rect 507 2290 518 2324
rect 552 2290 563 2324
rect 507 2256 563 2290
rect 507 2222 518 2256
rect 552 2222 563 2256
rect 507 2188 563 2222
rect 507 2154 518 2188
rect 552 2154 563 2188
rect 507 2120 563 2154
rect 507 2086 518 2120
rect 552 2086 563 2120
rect 507 2052 563 2086
rect 507 2018 518 2052
rect 552 2018 563 2052
rect 507 1984 563 2018
rect 507 1950 518 1984
rect 552 1950 563 1984
rect 507 1916 563 1950
rect 507 1882 518 1916
rect 552 1882 563 1916
rect 507 1848 563 1882
rect 507 1814 518 1848
rect 552 1814 563 1848
rect 507 1780 563 1814
rect 507 1746 518 1780
rect 552 1746 563 1780
rect 507 1712 563 1746
rect 507 1678 518 1712
rect 552 1678 563 1712
rect 507 1644 563 1678
rect 507 1610 518 1644
rect 552 1610 563 1644
rect 507 1576 563 1610
rect 507 1542 518 1576
rect 552 1542 563 1576
rect 507 1530 563 1542
rect 683 2460 739 2530
rect 683 2426 694 2460
rect 728 2426 739 2460
rect 683 2392 739 2426
rect 683 2358 694 2392
rect 728 2358 739 2392
rect 683 2324 739 2358
rect 683 2290 694 2324
rect 728 2290 739 2324
rect 683 2256 739 2290
rect 683 2222 694 2256
rect 728 2222 739 2256
rect 683 2188 739 2222
rect 683 2154 694 2188
rect 728 2154 739 2188
rect 683 2120 739 2154
rect 683 2086 694 2120
rect 728 2086 739 2120
rect 683 2052 739 2086
rect 683 2018 694 2052
rect 728 2018 739 2052
rect 683 1984 739 2018
rect 683 1950 694 1984
rect 728 1950 739 1984
rect 683 1916 739 1950
rect 683 1882 694 1916
rect 728 1882 739 1916
rect 683 1848 739 1882
rect 683 1814 694 1848
rect 728 1814 739 1848
rect 683 1780 739 1814
rect 683 1746 694 1780
rect 728 1746 739 1780
rect 683 1712 739 1746
rect 683 1678 694 1712
rect 728 1678 739 1712
rect 683 1644 739 1678
rect 683 1610 694 1644
rect 728 1610 739 1644
rect 683 1576 739 1610
rect 683 1542 694 1576
rect 728 1542 739 1576
rect 683 1530 739 1542
rect 859 2460 912 2530
rect 859 2426 870 2460
rect 904 2426 912 2460
rect 859 2392 912 2426
rect 859 2358 870 2392
rect 904 2358 912 2392
rect 859 2324 912 2358
rect 859 2290 870 2324
rect 904 2290 912 2324
rect 859 2256 912 2290
rect 859 2222 870 2256
rect 904 2222 912 2256
rect 859 2188 912 2222
rect 859 2154 870 2188
rect 904 2154 912 2188
rect 859 2120 912 2154
rect 859 2086 870 2120
rect 904 2086 912 2120
rect 859 2052 912 2086
rect 859 2018 870 2052
rect 904 2018 912 2052
rect 859 1984 912 2018
rect 859 1950 870 1984
rect 904 1950 912 1984
rect 859 1916 912 1950
rect 859 1882 870 1916
rect 904 1882 912 1916
rect 859 1848 912 1882
rect 859 1814 870 1848
rect 904 1814 912 1848
rect 859 1780 912 1814
rect 859 1746 870 1780
rect 904 1746 912 1780
rect 859 1712 912 1746
rect 859 1678 870 1712
rect 904 1678 912 1712
rect 859 1644 912 1678
rect 859 1610 870 1644
rect 904 1610 912 1644
rect 859 1576 912 1610
rect 859 1542 870 1576
rect 904 1542 912 1576
rect 859 1530 912 1542
<< mvndiffc >>
rect 166 1314 200 1348
rect 166 1246 200 1280
rect 166 1178 200 1212
rect 166 1110 200 1144
rect 564 1314 598 1348
rect 564 1246 598 1280
rect 564 1178 598 1212
rect 564 1110 598 1144
rect 964 1314 998 1348
rect 964 1246 998 1280
rect 964 1178 998 1212
rect 964 1110 998 1144
rect 166 848 200 882
rect 166 780 200 814
rect 166 712 200 746
rect 166 644 200 678
rect 564 848 598 882
rect 564 780 598 814
rect 564 712 598 746
rect 564 644 598 678
rect 964 848 998 882
rect 964 780 998 814
rect 964 712 998 746
rect 964 644 998 678
rect 166 302 200 336
rect 1022 302 1056 336
rect 166 147 200 181
rect 1022 147 1056 181
<< mvpdiffc >>
rect 166 2426 200 2460
rect 166 2358 200 2392
rect 166 2290 200 2324
rect 166 2222 200 2256
rect 166 2154 200 2188
rect 166 2086 200 2120
rect 166 2018 200 2052
rect 166 1950 200 1984
rect 166 1882 200 1916
rect 166 1814 200 1848
rect 166 1746 200 1780
rect 166 1678 200 1712
rect 166 1610 200 1644
rect 166 1542 200 1576
rect 342 2426 376 2460
rect 342 2358 376 2392
rect 342 2290 376 2324
rect 342 2222 376 2256
rect 342 2154 376 2188
rect 342 2086 376 2120
rect 342 2018 376 2052
rect 342 1950 376 1984
rect 342 1882 376 1916
rect 342 1814 376 1848
rect 342 1746 376 1780
rect 342 1678 376 1712
rect 342 1610 376 1644
rect 342 1542 376 1576
rect 518 2426 552 2460
rect 518 2358 552 2392
rect 518 2290 552 2324
rect 518 2222 552 2256
rect 518 2154 552 2188
rect 518 2086 552 2120
rect 518 2018 552 2052
rect 518 1950 552 1984
rect 518 1882 552 1916
rect 518 1814 552 1848
rect 518 1746 552 1780
rect 518 1678 552 1712
rect 518 1610 552 1644
rect 518 1542 552 1576
rect 694 2426 728 2460
rect 694 2358 728 2392
rect 694 2290 728 2324
rect 694 2222 728 2256
rect 694 2154 728 2188
rect 694 2086 728 2120
rect 694 2018 728 2052
rect 694 1950 728 1984
rect 694 1882 728 1916
rect 694 1814 728 1848
rect 694 1746 728 1780
rect 694 1678 728 1712
rect 694 1610 728 1644
rect 694 1542 728 1576
rect 870 2426 904 2460
rect 870 2358 904 2392
rect 870 2290 904 2324
rect 870 2222 904 2256
rect 870 2154 904 2188
rect 870 2086 904 2120
rect 870 2018 904 2052
rect 870 1950 904 1984
rect 870 1882 904 1916
rect 870 1814 904 1848
rect 870 1746 904 1780
rect 870 1678 904 1712
rect 870 1610 904 1644
rect 870 1542 904 1576
<< mvpsubdiff >>
rect 46 1323 84 1360
rect 46 1289 48 1323
rect 82 1289 84 1323
rect 46 1255 84 1289
rect 46 1221 48 1255
rect 82 1221 84 1255
rect 46 1187 84 1221
rect 46 1153 48 1187
rect 82 1153 84 1187
rect 46 1119 84 1153
rect 46 1085 48 1119
rect 82 1085 84 1119
rect 46 1051 84 1085
rect 46 1017 48 1051
rect 82 1017 84 1051
rect 46 983 84 1017
rect 46 949 48 983
rect 82 949 84 983
rect 46 915 84 949
rect 46 881 48 915
rect 82 881 84 915
rect 46 847 84 881
rect 46 813 48 847
rect 82 813 84 847
rect 46 779 84 813
rect 46 745 48 779
rect 82 745 84 779
rect 46 711 84 745
rect 46 677 48 711
rect 82 677 84 711
rect 46 643 84 677
rect 46 609 48 643
rect 82 609 84 643
rect 46 575 84 609
rect 46 541 48 575
rect 82 541 84 575
rect 46 507 84 541
rect 46 473 48 507
rect 82 473 84 507
rect 46 439 84 473
rect 46 405 48 439
rect 82 405 84 439
rect 46 371 84 405
rect 46 337 48 371
rect 82 337 84 371
rect 46 303 84 337
rect 46 269 48 303
rect 82 269 84 303
rect 46 235 84 269
rect 46 201 48 235
rect 82 201 84 235
rect 46 167 84 201
rect 46 133 48 167
rect 82 133 84 167
rect 46 99 84 133
rect 46 65 48 99
rect 82 65 84 99
rect 46 36 84 65
<< mvnsubdiff >>
rect 66 2485 104 2530
rect 66 2451 68 2485
rect 102 2451 104 2485
rect 66 2417 104 2451
rect 66 2383 68 2417
rect 102 2383 104 2417
rect 66 2349 104 2383
rect 66 2315 68 2349
rect 102 2315 104 2349
rect 66 2281 104 2315
rect 66 2247 68 2281
rect 102 2247 104 2281
rect 66 2213 104 2247
rect 66 2179 68 2213
rect 102 2179 104 2213
rect 66 2145 104 2179
rect 66 2111 68 2145
rect 102 2111 104 2145
rect 66 2077 104 2111
rect 66 2043 68 2077
rect 102 2043 104 2077
rect 66 2009 104 2043
rect 66 1975 68 2009
rect 102 1975 104 2009
rect 66 1941 104 1975
rect 66 1907 68 1941
rect 102 1907 104 1941
rect 66 1873 104 1907
rect 66 1839 68 1873
rect 102 1839 104 1873
rect 66 1798 104 1839
rect 66 1764 68 1798
rect 102 1764 104 1798
rect 66 1730 104 1764
rect 66 1696 68 1730
rect 102 1696 104 1730
rect 66 1662 104 1696
rect 66 1628 68 1662
rect 102 1628 104 1662
rect 66 1594 104 1628
rect 66 1560 68 1594
rect 102 1560 104 1594
rect 66 1530 104 1560
<< mvpsubdiffcont >>
rect 48 1289 82 1323
rect 48 1221 82 1255
rect 48 1153 82 1187
rect 48 1085 82 1119
rect 48 1017 82 1051
rect 48 949 82 983
rect 48 881 82 915
rect 48 813 82 847
rect 48 745 82 779
rect 48 677 82 711
rect 48 609 82 643
rect 48 541 82 575
rect 48 473 82 507
rect 48 405 82 439
rect 48 337 82 371
rect 48 269 82 303
rect 48 201 82 235
rect 48 133 82 167
rect 48 65 82 99
<< mvnsubdiffcont >>
rect 68 2451 102 2485
rect 68 2383 102 2417
rect 68 2315 102 2349
rect 68 2247 102 2281
rect 68 2179 102 2213
rect 68 2111 102 2145
rect 68 2043 102 2077
rect 68 1975 102 2009
rect 68 1907 102 1941
rect 68 1839 102 1873
rect 68 1764 102 1798
rect 68 1696 102 1730
rect 68 1628 102 1662
rect 68 1560 102 1594
<< poly >>
rect 211 2612 683 2632
rect 211 2578 240 2612
rect 274 2578 308 2612
rect 342 2578 376 2612
rect 410 2578 444 2612
rect 478 2578 512 2612
rect 546 2578 580 2612
rect 614 2578 683 2612
rect 211 2556 683 2578
rect 211 2530 331 2556
rect 387 2530 507 2556
rect 563 2530 683 2556
rect 739 2612 881 2632
rect 739 2578 759 2612
rect 793 2578 827 2612
rect 861 2578 881 2612
rect 739 2556 881 2578
rect 739 2530 859 2556
rect 1008 2536 1074 2552
rect 1008 2502 1024 2536
rect 1058 2502 1074 2536
rect 1008 2468 1074 2502
rect 1008 2434 1024 2468
rect 1058 2434 1074 2468
rect 1008 1600 1024 1634
rect 1058 1600 1074 1634
rect 1008 1566 1074 1600
rect 1008 1532 1024 1566
rect 1058 1532 1074 1566
rect 211 1504 331 1530
rect 387 1504 507 1530
rect 563 1504 683 1530
rect 739 1504 859 1530
rect 1008 1516 1074 1532
rect 1170 2536 1236 2552
rect 1170 2502 1186 2536
rect 1220 2502 1236 2536
rect 1170 2468 1236 2502
rect 1170 2434 1186 2468
rect 1220 2434 1236 2468
rect 211 1360 311 1504
rect 353 1442 555 1462
rect 353 1408 369 1442
rect 403 1408 437 1442
rect 471 1408 505 1442
rect 539 1408 555 1442
rect 353 1386 555 1408
rect 609 1442 811 1462
rect 609 1408 625 1442
rect 659 1408 693 1442
rect 727 1408 761 1442
rect 795 1408 811 1442
rect 609 1386 811 1408
rect 353 1360 553 1386
rect 609 1360 809 1386
rect 853 1360 953 1386
rect 211 1029 311 1060
rect 353 1034 553 1060
rect 609 1034 809 1060
rect 853 1034 953 1060
rect 177 1013 311 1029
rect 177 979 193 1013
rect 227 979 261 1013
rect 295 979 311 1013
rect 177 963 311 979
rect 211 932 311 963
rect 853 1013 995 1034
rect 853 979 869 1013
rect 903 979 937 1013
rect 971 979 995 1013
rect 853 958 995 979
rect 353 932 553 958
rect 609 932 809 958
rect 853 932 953 958
rect 211 476 311 632
rect 353 606 553 632
rect 609 606 809 632
rect 353 584 555 606
rect 353 550 369 584
rect 403 550 437 584
rect 471 550 505 584
rect 539 550 555 584
rect 353 530 555 550
rect 609 584 811 606
rect 609 550 625 584
rect 659 550 693 584
rect 727 550 761 584
rect 795 550 811 584
rect 609 530 811 550
rect 853 476 953 632
rect 211 456 1011 476
rect 211 422 231 456
rect 265 422 299 456
rect 333 422 367 456
rect 401 422 435 456
rect 469 422 503 456
rect 537 422 571 456
rect 605 422 639 456
rect 673 422 707 456
rect 741 422 775 456
rect 809 422 843 456
rect 877 422 911 456
rect 945 422 1011 456
rect 211 374 1011 422
rect 211 264 1011 290
rect 211 193 1011 219
rect 1170 200 1186 234
rect 1220 200 1236 234
rect 1170 166 1236 200
rect 1170 132 1186 166
rect 1220 132 1236 166
rect 1170 116 1236 132
rect 211 61 1011 109
rect 211 27 320 61
rect 354 27 388 61
rect 422 27 456 61
rect 490 27 524 61
rect 558 27 592 61
rect 626 27 660 61
rect 694 27 728 61
rect 762 27 796 61
rect 830 27 864 61
rect 898 27 932 61
rect 966 27 1011 61
rect 211 7 1011 27
<< polycont >>
rect 240 2578 274 2612
rect 308 2578 342 2612
rect 376 2578 410 2612
rect 444 2578 478 2612
rect 512 2578 546 2612
rect 580 2578 614 2612
rect 759 2578 793 2612
rect 827 2578 861 2612
rect 1024 2502 1058 2536
rect 1024 2434 1058 2468
rect 1024 1600 1058 1634
rect 1024 1532 1058 1566
rect 1186 2502 1220 2536
rect 1186 2434 1220 2468
rect 369 1408 403 1442
rect 437 1408 471 1442
rect 505 1408 539 1442
rect 625 1408 659 1442
rect 693 1408 727 1442
rect 761 1408 795 1442
rect 193 979 227 1013
rect 261 979 295 1013
rect 869 979 903 1013
rect 937 979 971 1013
rect 369 550 403 584
rect 437 550 471 584
rect 505 550 539 584
rect 625 550 659 584
rect 693 550 727 584
rect 761 550 795 584
rect 231 422 265 456
rect 299 422 333 456
rect 367 422 401 456
rect 435 422 469 456
rect 503 422 537 456
rect 571 422 605 456
rect 639 422 673 456
rect 707 422 741 456
rect 775 422 809 456
rect 843 422 877 456
rect 911 422 945 456
rect 1186 200 1220 234
rect 1186 132 1220 166
rect 320 27 354 61
rect 388 27 422 61
rect 456 27 490 61
rect 524 27 558 61
rect 592 27 626 61
rect 660 27 694 61
rect 728 27 762 61
rect 796 27 830 61
rect 864 27 898 61
rect 932 27 966 61
<< npolyres >>
rect 1008 1634 1074 2434
rect 1170 234 1236 2434
<< locali >>
rect 224 2578 240 2612
rect 274 2578 308 2612
rect 346 2578 376 2612
rect 410 2578 444 2612
rect 478 2578 512 2612
rect 546 2578 580 2612
rect 614 2578 630 2612
rect 743 2578 759 2612
rect 803 2578 827 2612
rect 875 2578 877 2612
rect 1008 2502 1024 2536
rect 1058 2502 1186 2536
rect 1220 2502 1240 2536
rect 68 2485 102 2501
rect 68 2417 102 2451
rect 68 2349 102 2383
rect 68 2281 102 2315
rect 68 2213 102 2247
rect 68 2145 102 2179
rect 68 2077 102 2111
rect 68 2009 102 2043
rect 68 1941 102 1975
rect 68 1873 102 1907
rect 68 1798 102 1839
rect 68 1754 102 1764
rect 68 1682 102 1696
rect 68 1610 102 1628
rect 68 1538 102 1560
rect 166 2460 200 2476
rect 166 2392 200 2426
rect 166 2324 200 2358
rect 166 2256 200 2290
rect 166 2188 200 2222
rect 166 2120 200 2154
rect 166 2052 200 2086
rect 166 1984 200 2018
rect 166 1916 200 1950
rect 166 1848 200 1882
rect 342 2460 376 2476
rect 342 2392 376 2426
rect 342 2324 376 2358
rect 342 2256 376 2290
rect 342 2188 376 2222
rect 342 2120 376 2154
rect 342 2052 376 2086
rect 342 1984 376 2018
rect 342 1916 376 1950
rect 342 1848 376 1882
rect 200 1806 238 1840
rect 518 2460 552 2476
rect 518 2392 552 2426
rect 518 2324 552 2358
rect 518 2256 552 2290
rect 518 2188 552 2222
rect 518 2120 552 2154
rect 518 2052 552 2086
rect 518 1984 552 2018
rect 518 1916 552 1950
rect 518 1848 552 1882
rect 166 1780 200 1806
rect 166 1712 200 1746
rect 166 1644 200 1678
rect 166 1576 200 1610
rect 166 1526 200 1542
rect 342 1780 376 1814
rect 694 2460 728 2476
rect 694 2392 728 2426
rect 694 2324 728 2358
rect 694 2256 728 2290
rect 694 2188 728 2222
rect 694 2120 728 2154
rect 694 2052 728 2086
rect 694 1984 728 2018
rect 694 1916 728 1950
rect 694 1848 728 1882
rect 552 1814 556 1840
rect 518 1806 556 1814
rect 870 2460 904 2476
rect 1008 2468 1240 2502
rect 1008 2434 1024 2468
rect 1058 2434 1186 2468
rect 1220 2434 1240 2468
rect 870 2392 904 2426
rect 870 2324 904 2358
rect 870 2256 904 2290
rect 870 2188 904 2222
rect 870 2120 904 2154
rect 870 2052 904 2086
rect 870 1984 904 2018
rect 870 1916 904 1950
rect 870 1848 904 1882
rect 1170 1840 1236 1914
rect 342 1712 376 1726
rect 342 1644 376 1654
rect 342 1576 376 1582
rect 342 1526 376 1542
rect 518 1780 552 1806
rect 518 1712 552 1746
rect 518 1644 552 1678
rect 518 1576 552 1610
rect 518 1526 552 1542
rect 694 1780 728 1814
rect 828 1806 866 1840
rect 900 1806 904 1814
rect 1024 1806 1062 1840
rect 1096 1806 1236 1840
rect 694 1712 728 1726
rect 694 1644 728 1654
rect 694 1576 728 1582
rect 694 1526 728 1542
rect 870 1780 904 1806
rect 870 1712 904 1746
rect 870 1644 904 1678
rect 870 1576 904 1610
rect 870 1526 904 1542
rect 1008 1634 1074 1806
rect 1008 1600 1024 1634
rect 1058 1600 1074 1634
rect 1008 1566 1074 1600
rect 1008 1532 1024 1566
rect 1058 1532 1074 1566
rect 353 1408 369 1442
rect 403 1408 437 1442
rect 471 1408 505 1442
rect 539 1408 555 1442
rect 609 1408 625 1442
rect 659 1408 693 1442
rect 727 1408 761 1442
rect 795 1408 811 1442
rect 48 1323 82 1352
rect 48 1255 82 1289
rect 48 1187 82 1206
rect 48 1119 82 1134
rect 48 1051 82 1062
rect 48 983 82 1017
rect 48 915 82 949
rect 48 847 82 881
rect 48 779 82 813
rect 48 711 82 716
rect 48 643 82 644
rect 116 1348 200 1364
rect 116 1314 166 1348
rect 116 1280 200 1314
rect 116 1246 166 1280
rect 116 1212 200 1246
rect 116 1178 166 1212
rect 116 1144 200 1178
rect 116 1110 166 1144
rect 116 1094 200 1110
rect 564 1348 598 1364
rect 564 1280 598 1314
rect 564 1234 598 1246
rect 564 1162 598 1178
rect 116 898 150 1094
rect 564 1090 598 1110
rect 964 1348 1059 1364
rect 998 1314 1059 1348
rect 964 1280 1059 1314
rect 998 1246 1059 1280
rect 964 1212 1059 1246
rect 998 1178 1059 1212
rect 964 1144 1059 1178
rect 998 1110 1059 1144
rect 964 1094 1059 1110
rect 193 1013 295 1029
rect 227 1006 261 1013
rect 869 1013 971 1029
rect 234 979 261 1006
rect 193 972 200 979
rect 234 972 272 979
rect 903 979 937 1013
rect 193 963 295 972
rect 901 970 939 979
rect 869 963 971 970
rect 1025 898 1059 1094
rect 1170 972 1236 1806
rect 1152 938 1190 972
rect 1224 938 1236 972
rect 116 882 200 898
rect 116 848 166 882
rect 116 830 200 848
rect 564 882 598 898
rect 116 814 178 830
rect 116 780 166 814
rect 212 796 250 830
rect 564 814 598 848
rect 964 882 1059 898
rect 998 848 1059 882
rect 964 830 1059 848
rect 1170 830 1236 836
rect 116 746 200 780
rect 116 712 166 746
rect 116 678 200 712
rect 116 644 166 678
rect 116 628 200 644
rect 912 796 950 830
rect 984 814 1059 830
rect 564 750 598 780
rect 564 678 598 712
rect 564 628 598 644
rect 998 780 1059 814
rect 1152 796 1190 830
rect 1224 796 1236 830
rect 964 746 1059 780
rect 998 712 1059 746
rect 964 678 1059 712
rect 998 644 1059 678
rect 964 628 1059 644
rect 48 575 82 609
rect 353 550 369 584
rect 403 550 437 584
rect 471 550 505 584
rect 539 550 555 584
rect 609 550 625 584
rect 659 550 693 584
rect 727 550 761 584
rect 795 550 811 584
rect 48 507 82 541
rect 48 439 82 473
rect 215 422 223 456
rect 265 422 295 456
rect 333 422 367 456
rect 401 422 435 456
rect 469 422 503 456
rect 537 422 571 456
rect 605 422 639 456
rect 673 422 707 456
rect 741 422 775 456
rect 809 422 843 456
rect 877 422 911 456
rect 945 422 961 456
rect 48 371 82 405
rect 48 303 82 337
rect 48 235 82 269
rect 48 167 82 201
rect 48 99 82 100
rect 166 336 200 352
rect 166 181 200 302
rect 1022 340 1056 352
rect 1022 268 1056 302
rect 1170 234 1236 796
rect 166 98 200 147
rect 901 180 939 214
rect 1170 200 1186 234
rect 1220 200 1236 234
rect 48 62 82 65
rect 867 61 973 180
rect 1022 181 1056 197
rect 1022 134 1056 147
rect 1170 166 1236 200
rect 1170 132 1186 166
rect 1220 132 1236 166
rect 1022 62 1056 100
rect 304 27 320 61
rect 354 27 388 61
rect 422 27 456 61
rect 490 27 524 61
rect 558 27 592 61
rect 626 27 660 61
rect 694 27 728 61
rect 762 27 796 61
rect 830 27 864 61
rect 898 27 932 61
rect 966 27 982 61
<< viali >>
rect 240 2578 274 2612
rect 312 2578 342 2612
rect 342 2578 346 2612
rect 769 2578 793 2612
rect 793 2578 803 2612
rect 841 2578 861 2612
rect 861 2578 875 2612
rect 68 1730 102 1754
rect 68 1720 102 1730
rect 68 1662 102 1682
rect 68 1648 102 1662
rect 68 1594 102 1610
rect 68 1576 102 1594
rect 166 1814 200 1840
rect 166 1806 200 1814
rect 238 1806 272 1840
rect 484 1806 518 1840
rect 556 1806 590 1840
rect 342 1746 376 1760
rect 342 1726 376 1746
rect 342 1678 376 1688
rect 342 1654 376 1678
rect 342 1610 376 1616
rect 342 1582 376 1610
rect 794 1806 828 1840
rect 866 1814 870 1840
rect 870 1814 900 1840
rect 866 1806 900 1814
rect 990 1806 1024 1840
rect 1062 1806 1096 1840
rect 694 1746 728 1760
rect 694 1726 728 1746
rect 694 1678 728 1688
rect 694 1654 728 1678
rect 694 1610 728 1616
rect 694 1582 728 1610
rect 48 1221 82 1240
rect 48 1206 82 1221
rect 48 1153 82 1168
rect 48 1134 82 1153
rect 48 1085 82 1096
rect 48 1062 82 1085
rect 48 745 82 750
rect 48 716 82 745
rect 48 677 82 678
rect 48 644 82 677
rect 564 1212 598 1234
rect 564 1200 598 1212
rect 564 1144 598 1162
rect 564 1128 598 1144
rect 564 1056 598 1090
rect 200 979 227 1006
rect 227 979 234 1006
rect 272 979 295 1006
rect 295 979 306 1006
rect 200 972 234 979
rect 272 972 306 979
rect 867 979 869 1004
rect 869 979 901 1004
rect 939 979 971 1004
rect 971 979 973 1004
rect 867 970 901 979
rect 939 970 973 979
rect 1118 938 1152 972
rect 1190 938 1224 972
rect 178 814 212 830
rect 178 796 200 814
rect 200 796 212 814
rect 250 796 284 830
rect 878 796 912 830
rect 950 814 984 830
rect 950 796 964 814
rect 964 796 984 814
rect 564 746 598 750
rect 564 716 598 746
rect 564 644 598 678
rect 1118 796 1152 830
rect 1190 796 1224 830
rect 223 422 231 456
rect 231 422 257 456
rect 295 422 299 456
rect 299 422 329 456
rect 48 133 82 134
rect 48 100 82 133
rect 1022 336 1056 340
rect 1022 306 1056 336
rect 1022 234 1056 268
rect 867 180 901 214
rect 939 180 973 214
rect 48 28 82 62
rect 1022 100 1056 134
rect 1022 28 1056 62
<< metal1 >>
rect 211 2616 391 2622
rect 263 2612 275 2616
rect 327 2612 339 2616
rect 274 2578 275 2612
rect 263 2564 275 2578
rect 327 2564 339 2578
rect 211 2558 391 2564
rect 757 2616 933 2622
rect 757 2612 817 2616
rect 869 2612 881 2616
rect 757 2578 769 2612
rect 803 2578 817 2612
rect 875 2578 881 2612
rect 757 2564 817 2578
rect 869 2564 881 2578
rect 757 2558 933 2564
rect 1013 1922 1065 1928
tri 985 1846 1013 1874 se
rect 1013 1858 1065 1870
rect 0 1840 1013 1846
tri 1065 1846 1093 1874 sw
rect 1065 1840 1236 1846
rect 0 1806 166 1840
rect 200 1806 238 1840
rect 272 1806 484 1840
rect 518 1806 556 1840
rect 590 1806 794 1840
rect 828 1806 866 1840
rect 900 1806 990 1840
rect 1096 1806 1236 1840
rect 0 1800 1236 1806
rect 0 1760 1284 1772
rect 0 1754 342 1760
rect 0 1720 68 1754
rect 102 1726 342 1754
rect 376 1726 694 1760
rect 728 1726 1284 1760
rect 102 1720 1284 1726
rect 0 1688 1284 1720
rect 0 1682 342 1688
rect 0 1648 68 1682
rect 102 1654 342 1682
rect 376 1654 694 1688
rect 728 1654 1284 1688
rect 102 1648 1284 1654
rect 0 1616 1284 1648
rect 0 1610 342 1616
rect 0 1576 68 1610
rect 102 1582 342 1610
rect 376 1582 694 1616
rect 728 1582 1284 1616
rect 102 1576 1284 1582
rect 0 1570 1284 1576
rect 0 1240 1284 1246
rect 0 1206 48 1240
rect 82 1234 1284 1240
rect 82 1206 564 1234
rect 0 1200 564 1206
rect 598 1200 1111 1234
rect 0 1182 1111 1200
rect 1163 1182 1284 1234
rect 0 1170 1284 1182
rect 0 1168 1111 1170
rect 0 1134 48 1168
rect 82 1162 1111 1168
rect 82 1134 564 1162
rect 0 1128 564 1134
rect 598 1128 1111 1162
rect 0 1118 1111 1128
rect 1163 1118 1284 1170
rect 0 1106 1284 1118
rect 0 1096 1111 1106
rect 0 1062 48 1096
rect 82 1090 1111 1096
rect 82 1062 564 1090
rect 0 1056 564 1062
rect 598 1056 1111 1090
rect 0 1054 1111 1056
rect 1163 1054 1284 1106
rect 0 1044 1284 1054
rect 188 1006 217 1016
rect 269 1006 281 1016
rect 188 972 200 1006
rect 269 972 272 1006
rect 333 1004 985 1016
rect 188 964 217 972
rect 269 964 281 972
rect 333 970 867 1004
rect 901 970 939 1004
rect 973 970 985 1004
rect 333 964 985 970
rect 1106 972 1236 978
rect 1106 938 1118 972
rect 1152 938 1190 972
rect 1224 938 1236 972
rect 1106 932 1236 938
tri 1156 904 1184 932 ne
rect 1184 904 1236 932
rect 1185 902 1235 903
rect 1184 866 1236 902
rect 1185 865 1235 866
tri 1156 836 1184 864 se
rect 1184 836 1236 864
rect 166 830 1236 836
rect 166 796 178 830
rect 212 796 250 830
rect 284 796 878 830
rect 912 796 950 830
rect 984 796 1118 830
rect 1152 796 1190 830
rect 1224 796 1236 830
rect 166 790 1236 796
rect 0 754 1284 762
rect 0 750 1111 754
rect 0 716 48 750
rect 82 716 564 750
rect 598 716 1111 750
rect 0 702 1111 716
rect 1163 702 1284 754
rect 0 690 1284 702
rect 0 678 1111 690
rect 0 644 48 678
rect 82 644 564 678
rect 598 644 1111 678
rect 0 638 1111 644
rect 1163 638 1284 690
rect 0 632 1284 638
rect 211 418 217 470
rect 269 418 281 470
rect 333 418 341 470
rect 211 416 341 418
rect 1013 340 1065 352
rect 933 296 985 302
tri 919 234 933 248 se
rect 933 234 985 244
tri 905 220 919 234 se
rect 919 232 985 234
rect 919 220 933 232
rect 855 214 933 220
rect 1013 276 1065 288
rect 1013 218 1065 224
rect 855 180 867 214
rect 901 180 933 214
rect 855 174 985 180
rect 42 140 1169 146
rect 42 134 1111 140
rect 42 100 48 134
rect 82 100 1022 134
rect 1056 100 1111 134
rect 42 88 1111 100
rect 1163 88 1169 140
rect 42 76 1169 88
rect 42 62 1111 76
rect 42 28 48 62
rect 82 28 1022 62
rect 1056 28 1111 62
rect 42 24 1111 28
rect 1163 24 1169 76
rect 42 16 1169 24
<< rmetal1 >>
rect 1184 903 1236 904
rect 1184 902 1185 903
rect 1235 902 1236 903
rect 1184 865 1185 866
rect 1235 865 1236 866
rect 1184 864 1236 865
<< via1 >>
rect 211 2612 263 2616
rect 275 2612 327 2616
rect 339 2612 391 2616
rect 211 2578 240 2612
rect 240 2578 263 2612
rect 275 2578 312 2612
rect 312 2578 327 2612
rect 339 2578 346 2612
rect 346 2578 391 2612
rect 211 2564 263 2578
rect 275 2564 327 2578
rect 339 2564 391 2578
rect 817 2612 869 2616
rect 817 2578 841 2612
rect 841 2578 869 2612
rect 817 2564 869 2578
rect 881 2564 933 2616
rect 1013 1870 1065 1922
rect 1013 1840 1065 1858
rect 1013 1806 1024 1840
rect 1024 1806 1062 1840
rect 1062 1806 1065 1840
rect 1111 1182 1163 1234
rect 1111 1118 1163 1170
rect 1111 1054 1163 1106
rect 217 1006 269 1016
rect 281 1006 333 1016
rect 217 972 234 1006
rect 234 972 269 1006
rect 281 972 306 1006
rect 306 972 333 1006
rect 217 964 269 972
rect 281 964 333 972
rect 1111 702 1163 754
rect 1111 638 1163 690
rect 217 456 269 470
rect 217 422 223 456
rect 223 422 257 456
rect 257 422 269 456
rect 217 418 269 422
rect 281 456 333 470
rect 281 422 295 456
rect 295 422 329 456
rect 329 422 333 456
rect 281 418 333 422
rect 1013 306 1022 340
rect 1022 306 1056 340
rect 1056 306 1065 340
rect 933 244 985 296
rect 933 214 985 232
rect 1013 288 1065 306
rect 1013 268 1065 276
rect 1013 234 1022 268
rect 1022 234 1056 268
rect 1056 234 1065 268
rect 1013 224 1065 234
rect 933 180 939 214
rect 939 180 973 214
rect 973 180 985 214
rect 1111 88 1163 140
rect 1111 24 1163 76
<< metal2 >>
rect 211 2616 391 2622
rect 263 2564 275 2616
rect 327 2564 339 2616
rect 211 2558 391 2564
rect 817 2616 985 2622
rect 869 2564 881 2616
rect 933 2564 985 2616
rect 817 2558 985 2564
rect 211 1016 263 2558
tri 263 2530 291 2558 nw
tri 905 2530 933 2558 ne
tri 263 1016 291 1044 sw
rect 211 964 217 1016
rect 269 964 281 1016
rect 333 964 339 1016
rect 211 470 263 964
tri 263 936 291 964 nw
tri 263 470 291 498 sw
rect 211 418 217 470
rect 269 418 281 470
rect 333 418 339 470
rect 933 296 985 2558
rect 933 232 985 244
rect 1013 1922 1065 1928
rect 1013 1858 1065 1870
rect 1013 340 1065 1806
rect 1013 276 1065 288
rect 1013 218 1065 224
rect 1105 1234 1169 1246
rect 1105 1182 1111 1234
rect 1163 1182 1169 1234
rect 1105 1170 1169 1182
rect 1105 1118 1111 1170
rect 1163 1118 1169 1170
rect 1105 1106 1169 1118
rect 1105 1054 1111 1106
rect 1163 1054 1169 1106
rect 1105 754 1169 1054
rect 1105 702 1111 754
rect 1163 702 1169 754
rect 1105 690 1169 702
rect 1105 638 1111 690
rect 1163 638 1169 690
rect 933 174 985 180
rect 1105 140 1169 638
rect 1105 88 1111 140
rect 1163 88 1169 140
rect 1105 76 1169 88
rect 1105 24 1111 76
rect 1163 24 1169 76
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1666199351
transform 0 1 1184 1 0 812
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808281  sky130_fd_pr__nfet_01v8__example_55959141808281_0
timestamp 1666199351
transform 1 0 211 0 1 290
box -1 0 801 1
use sky130_fd_pr__nfet_01v8__example_55959141808282  sky130_fd_pr__nfet_01v8__example_55959141808282_0
timestamp 1666199351
transform 1 0 211 0 1 632
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808282  sky130_fd_pr__nfet_01v8__example_55959141808282_1
timestamp 1666199351
transform -1 0 953 0 1 632
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808282  sky130_fd_pr__nfet_01v8__example_55959141808282_2
timestamp 1666199351
transform -1 0 953 0 -1 1360
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808282  sky130_fd_pr__nfet_01v8__example_55959141808282_3
timestamp 1666199351
transform 1 0 211 0 -1 1360
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808287  sky130_fd_pr__nfet_01v8__example_55959141808287_0
timestamp 1666199351
transform -1 0 553 0 1 632
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808287  sky130_fd_pr__nfet_01v8__example_55959141808287_1
timestamp 1666199351
transform 1 0 609 0 1 632
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808287  sky130_fd_pr__nfet_01v8__example_55959141808287_2
timestamp 1666199351
transform 1 0 609 0 -1 1360
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808287  sky130_fd_pr__nfet_01v8__example_55959141808287_3
timestamp 1666199351
transform -1 0 553 0 -1 1360
box -1 0 0 1
use sky130_fd_pr__nfet_01v8__example_55959141808644  sky130_fd_pr__nfet_01v8__example_55959141808644_0
timestamp 1666199351
transform -1 0 1011 0 -1 193
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808283  sky130_fd_pr__pfet_01v8__example_55959141808283_0
timestamp 1666199351
transform -1 0 683 0 1 1530
box -1 0 473 1
use sky130_fd_pr__pfet_01v8__example_55959141808284  sky130_fd_pr__pfet_01v8__example_55959141808284_0
timestamp 1666199351
transform 1 0 739 0 1 1530
box -1 0 121 1
use sky130_fd_pr__res_generic_po__example_55959141808285  sky130_fd_pr__res_generic_po__example_55959141808285_0
timestamp 1666199351
transform 0 -1 1074 -1 0 2434
box 15 0 785 1
use sky130_fd_pr__res_generic_po__example_55959141808286  sky130_fd_pr__res_generic_po__example_55959141808286_0
timestamp 1666199351
transform 0 -1 1236 -1 0 2434
box 15 0 2185 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1666199351
transform -1 0 973 0 -1 214
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1666199351
transform 0 1 48 1 0 28
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1666199351
transform 1 0 1118 0 -1 972
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1666199351
transform 0 1 1022 1 0 234
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1666199351
transform 1 0 990 0 -1 1840
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1666199351
transform 0 1 564 1 0 644
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1666199351
transform -1 0 284 0 1 796
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1666199351
transform 1 0 1118 0 -1 830
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1666199351
transform -1 0 984 0 1 796
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1666199351
transform 1 0 200 0 1 972
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1666199351
transform 1 0 794 0 1 1806
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1666199351
transform 1 0 484 0 1 1806
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1666199351
transform 1 0 166 0 1 1806
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1666199351
transform 1 0 867 0 1 970
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1666199351
transform 0 -1 1056 1 0 28
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1666199351
transform -1 0 875 0 -1 2612
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1666199351
transform 0 1 48 1 0 644
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1666199351
transform 1 0 240 0 1 2578
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1666199351
transform 1 0 223 0 -1 456
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1666199351
transform 0 1 564 -1 0 1234
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1666199351
transform 0 -1 728 -1 0 1760
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1666199351
transform 0 -1 376 -1 0 1760
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1666199351
transform 1 0 68 0 1 1576
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1666199351
transform -1 0 82 0 1 1062
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1666199351
transform 0 1 933 1 0 174
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1666199351
transform 0 -1 1065 1 0 218
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1666199351
transform 0 1 1013 1 0 1800
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1666199351
transform 1 0 211 0 1 418
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1666199351
transform 1 0 211 0 1 964
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_0
timestamp 1666199351
transform 0 -1 933 1 0 2558
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_1
timestamp 1666199351
transform 1 0 1105 0 -1 140
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_2
timestamp 1666199351
transform 1 0 1105 0 -1 754
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808276  sky130_fd_pr__via_m1m2__example_55959141808276_0
timestamp 1666199351
transform 1 0 1105 0 -1 1234
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808276  sky130_fd_pr__via_m1m2__example_55959141808276_1
timestamp 1666199351
transform 0 -1 391 1 0 2558
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1666199351
transform 0 1 1170 -1 0 250
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1666199351
transform 0 1 1008 -1 0 2552
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1666199351
transform -1 0 987 0 -1 1029
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1666199351
transform -1 0 311 0 -1 1029
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_4
timestamp 1666199351
transform 0 1 1008 -1 0 1650
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_5
timestamp 1666199351
transform 0 1 1170 -1 0 2552
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1666199351
transform 0 1 743 1 0 2562
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808272  sky130_fd_pr__via_pol1__example_55959141808272_0
timestamp 1666199351
transform 0 1 224 1 0 2562
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1666199351
transform 0 -1 961 1 0 406
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1666199351
transform 0 1 353 1 0 1392
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_1
timestamp 1666199351
transform 0 1 609 1 0 534
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_2
timestamp 1666199351
transform 0 1 609 1 0 1392
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_3
timestamp 1666199351
transform 0 1 353 1 0 534
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808275  sky130_fd_pr__via_pol1__example_55959141808275_0
timestamp 1666199351
transform 0 -1 982 -1 0 77
box 0 0 1 1
<< labels >>
flabel comment s 180 210 180 210 0 FreeSans 300 90 0 0 N<2>
flabel comment s 1190 2501 1190 2501 0 FreeSans 300 0 0 0 INT_RES
flabel metal2 s 211 1402 263 1454 7 FreeSans 300 0 0 0 DRVHI_H
port 1 nsew
flabel metal2 s 919 2558 985 2622 3 FreeSans 300 0 0 0 PUEN_H
port 2 nsew
flabel locali s 357 1408 407 1442 3 FreeSans 300 270 0 0 EN_FAST[0]
port 3 nsew
flabel locali s 761 1408 811 1442 3 FreeSans 300 270 0 0 EN_FAST[1]
port 4 nsew
flabel locali s 613 550 663 584 3 FreeSans 300 270 0 0 EN_FAST[2]
port 5 nsew
flabel locali s 357 550 407 584 3 FreeSans 300 270 0 0 EN_FAST[3]
port 6 nsew
flabel metal1 s 1242 1044 1284 1246 7 FreeSans 300 180 0 0 VGND_IO
port 7 nsew
flabel metal1 s 1247 1570 1284 1772 6 FreeSans 300 180 0 0 VCC_IO
port 8 nsew
flabel metal1 s 1196 1800 1236 1846 7 FreeSans 300 0 0 0 PU_H_N
port 9 nsew
flabel metal1 s 0 1044 36 1246 7 FreeSans 300 0 0 0 VGND_IO
port 7 nsew
flabel metal1 s 0 1570 36 1772 6 FreeSans 300 0 0 0 VCC_IO
port 8 nsew
flabel metal1 s 0 1800 36 1846 3 FreeSans 300 180 0 0 PU_H_N
port 9 nsew
flabel metal1 s 1242 632 1284 762 7 FreeSans 300 180 0 0 VGND_IO
port 7 nsew
flabel metal1 s 0 632 36 762 7 FreeSans 300 0 0 0 VGND_IO
port 7 nsew
<< properties >>
string GDS_END 48850390
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48837118
<< end >>
