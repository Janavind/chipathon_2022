magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 2382 201 2851 203
rect 1236 157 1690 201
rect 2015 157 2851 201
rect 1 21 2851 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 423 47 453 131
rect 618 47 648 131
rect 705 47 735 131
rect 792 47 822 131
rect 887 47 917 119
rect 1000 47 1030 119
rect 1102 47 1132 131
rect 1211 47 1241 131
rect 1312 47 1342 175
rect 1396 47 1426 175
rect 1584 47 1614 175
rect 1684 47 1714 119
rect 1792 47 1822 119
rect 1887 47 1917 131
rect 1974 47 2004 131
rect 2091 47 2121 175
rect 2175 47 2205 175
rect 2363 47 2393 131
rect 2460 47 2490 177
rect 2648 47 2678 131
rect 2743 47 2773 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 363 381 491
rect 423 363 453 491
rect 638 413 668 497
rect 722 413 752 497
rect 806 413 836 497
rect 903 413 933 497
rect 987 413 1017 497
rect 1107 413 1137 497
rect 1213 413 1243 497
rect 1321 329 1351 497
rect 1405 329 1435 497
rect 1542 329 1572 497
rect 1686 413 1716 497
rect 1770 413 1800 497
rect 1888 413 1918 497
rect 1996 413 2026 497
rect 2092 329 2122 497
rect 2164 329 2194 497
rect 2363 301 2393 429
rect 2460 297 2490 497
rect 2648 353 2678 481
rect 2743 297 2773 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 111 351 131
rect 299 77 307 111
rect 341 77 351 111
rect 299 47 351 77
rect 381 47 423 131
rect 453 103 512 131
rect 453 69 470 103
rect 504 69 512 103
rect 453 47 512 69
rect 566 111 618 131
rect 566 77 574 111
rect 608 77 618 111
rect 566 47 618 77
rect 648 89 705 131
rect 648 55 661 89
rect 695 55 705 89
rect 648 47 705 55
rect 735 47 792 131
rect 822 119 872 131
rect 1262 131 1312 175
rect 1045 119 1102 131
rect 822 103 887 119
rect 822 69 832 103
rect 866 69 887 103
rect 822 47 887 69
rect 917 93 1000 119
rect 917 59 927 93
rect 961 59 1000 93
rect 917 47 1000 59
rect 1030 47 1102 119
rect 1132 89 1211 131
rect 1132 55 1167 89
rect 1201 55 1211 89
rect 1132 47 1211 55
rect 1241 93 1312 131
rect 1241 59 1268 93
rect 1302 59 1312 93
rect 1241 47 1312 59
rect 1342 156 1396 175
rect 1342 122 1352 156
rect 1386 122 1396 156
rect 1342 47 1396 122
rect 1426 127 1478 175
rect 1426 93 1436 127
rect 1470 93 1478 127
rect 1426 47 1478 93
rect 1532 93 1584 175
rect 1532 59 1540 93
rect 1574 59 1584 93
rect 1532 47 1584 59
rect 1614 119 1664 175
rect 2041 131 2091 175
rect 1837 119 1887 131
rect 1614 47 1684 119
rect 1714 93 1792 119
rect 1714 59 1739 93
rect 1773 59 1792 93
rect 1714 47 1792 59
rect 1822 47 1887 119
rect 1917 89 1974 131
rect 1917 55 1930 89
rect 1964 55 1974 89
rect 1917 47 1974 55
rect 2004 109 2091 131
rect 2004 75 2032 109
rect 2066 75 2091 109
rect 2004 47 2091 75
rect 2121 153 2175 175
rect 2121 119 2131 153
rect 2165 119 2175 153
rect 2121 47 2175 119
rect 2205 101 2257 175
rect 2408 161 2460 177
rect 2408 131 2416 161
rect 2205 67 2215 101
rect 2249 67 2257 101
rect 2205 47 2257 67
rect 2311 103 2363 131
rect 2311 69 2319 103
rect 2353 69 2363 103
rect 2311 47 2363 69
rect 2393 127 2416 131
rect 2450 127 2460 161
rect 2393 93 2460 127
rect 2393 59 2416 93
rect 2450 59 2460 93
rect 2393 47 2460 59
rect 2490 127 2542 177
rect 2693 131 2743 177
rect 2490 93 2500 127
rect 2534 93 2542 127
rect 2490 47 2542 93
rect 2596 119 2648 131
rect 2596 85 2604 119
rect 2638 85 2648 119
rect 2596 47 2648 85
rect 2678 93 2743 131
rect 2678 59 2699 93
rect 2733 59 2743 93
rect 2678 47 2743 59
rect 2773 129 2825 177
rect 2773 95 2783 129
rect 2817 95 2825 129
rect 2773 47 2825 95
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 479 351 491
rect 299 445 307 479
rect 341 445 351 479
rect 299 411 351 445
rect 299 377 307 411
rect 341 377 351 411
rect 299 363 351 377
rect 381 363 423 491
rect 453 477 505 491
rect 453 443 463 477
rect 497 443 505 477
rect 453 409 505 443
rect 586 477 638 497
rect 586 443 594 477
rect 628 443 638 477
rect 586 413 638 443
rect 668 477 722 497
rect 668 443 678 477
rect 712 443 722 477
rect 668 413 722 443
rect 752 413 806 497
rect 836 477 903 497
rect 836 443 846 477
rect 880 443 903 477
rect 836 413 903 443
rect 933 484 987 497
rect 933 450 943 484
rect 977 450 987 484
rect 933 413 987 450
rect 1017 413 1107 497
rect 1137 475 1213 497
rect 1137 441 1157 475
rect 1191 441 1213 475
rect 1137 413 1213 441
rect 1243 459 1321 497
rect 1243 425 1277 459
rect 1311 425 1321 459
rect 1243 413 1321 425
rect 453 375 463 409
rect 497 375 505 409
rect 453 363 505 375
rect 1259 391 1321 413
rect 1259 357 1277 391
rect 1311 357 1321 391
rect 1259 329 1321 357
rect 1351 329 1405 497
rect 1435 485 1542 497
rect 1435 451 1451 485
rect 1485 451 1542 485
rect 1435 417 1542 451
rect 1435 383 1451 417
rect 1485 383 1542 417
rect 1435 329 1542 383
rect 1572 413 1686 497
rect 1716 484 1770 497
rect 1716 450 1726 484
rect 1760 450 1770 484
rect 1716 413 1770 450
rect 1800 413 1888 497
rect 1918 485 1996 497
rect 1918 451 1940 485
rect 1974 451 1996 485
rect 1918 413 1996 451
rect 2026 459 2092 497
rect 2026 425 2048 459
rect 2082 425 2092 459
rect 2026 413 2092 425
rect 1572 329 1624 413
rect 2041 329 2092 413
rect 2122 329 2164 497
rect 2194 485 2246 497
rect 2194 451 2204 485
rect 2238 451 2246 485
rect 2408 485 2460 497
rect 2194 329 2246 451
rect 2408 451 2416 485
rect 2450 451 2460 485
rect 2408 429 2460 451
rect 2311 349 2363 429
rect 2311 315 2319 349
rect 2353 315 2363 349
rect 2311 301 2363 315
rect 2393 301 2460 429
rect 2410 297 2460 301
rect 2490 448 2542 497
rect 2693 481 2743 497
rect 2490 414 2500 448
rect 2534 414 2542 448
rect 2490 380 2542 414
rect 2490 346 2500 380
rect 2534 346 2542 380
rect 2596 467 2648 481
rect 2596 433 2604 467
rect 2638 433 2648 467
rect 2596 399 2648 433
rect 2596 365 2604 399
rect 2638 365 2648 399
rect 2596 353 2648 365
rect 2678 473 2743 481
rect 2678 439 2699 473
rect 2733 439 2743 473
rect 2678 405 2743 439
rect 2678 371 2698 405
rect 2732 371 2743 405
rect 2678 353 2743 371
rect 2490 297 2542 346
rect 2693 297 2743 353
rect 2773 449 2825 497
rect 2773 415 2783 449
rect 2817 415 2825 449
rect 2773 381 2825 415
rect 2773 347 2783 381
rect 2817 347 2825 381
rect 2773 297 2825 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 77 341 111
rect 470 69 504 103
rect 574 77 608 111
rect 661 55 695 89
rect 832 69 866 103
rect 927 59 961 93
rect 1167 55 1201 89
rect 1268 59 1302 93
rect 1352 122 1386 156
rect 1436 93 1470 127
rect 1540 59 1574 93
rect 1739 59 1773 93
rect 1930 55 1964 89
rect 2032 75 2066 109
rect 2131 119 2165 153
rect 2215 67 2249 101
rect 2319 69 2353 103
rect 2416 127 2450 161
rect 2416 59 2450 93
rect 2500 93 2534 127
rect 2604 85 2638 119
rect 2699 59 2733 93
rect 2783 95 2817 129
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 445 341 479
rect 307 377 341 411
rect 463 443 497 477
rect 594 443 628 477
rect 678 443 712 477
rect 846 443 880 477
rect 943 450 977 484
rect 1157 441 1191 475
rect 1277 425 1311 459
rect 463 375 497 409
rect 1277 357 1311 391
rect 1451 451 1485 485
rect 1451 383 1485 417
rect 1726 450 1760 484
rect 1940 451 1974 485
rect 2048 425 2082 459
rect 2204 451 2238 485
rect 2416 451 2450 485
rect 2319 315 2353 349
rect 2500 414 2534 448
rect 2500 346 2534 380
rect 2604 433 2638 467
rect 2604 365 2638 399
rect 2699 439 2733 473
rect 2698 371 2732 405
rect 2783 415 2817 449
rect 2783 347 2817 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 491 381 517
rect 423 491 453 517
rect 638 497 668 523
rect 722 497 752 523
rect 806 497 836 523
rect 903 497 933 523
rect 987 497 1017 523
rect 1107 497 1137 523
rect 1213 497 1243 523
rect 1321 497 1351 523
rect 1405 497 1435 523
rect 1542 497 1572 523
rect 1686 497 1716 523
rect 1770 497 1800 523
rect 1888 497 1918 523
rect 1996 497 2026 523
rect 2092 497 2122 523
rect 2164 497 2194 523
rect 2460 497 2490 523
rect 638 397 668 413
rect 722 397 752 413
rect 542 365 596 381
rect 79 348 109 363
rect 45 318 109 348
rect 45 280 75 318
rect 21 264 75 280
rect 163 274 193 363
rect 351 331 381 363
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 117 264 193 274
rect 295 315 381 331
rect 423 345 453 363
rect 542 345 552 365
rect 423 331 552 345
rect 586 331 596 365
rect 423 318 596 331
rect 638 367 752 397
rect 423 317 594 318
rect 423 315 592 317
rect 295 281 305 315
rect 339 301 381 315
rect 339 281 349 301
rect 638 281 668 367
rect 806 325 836 413
rect 295 265 349 281
rect 117 230 133 264
rect 167 230 193 264
rect 117 220 193 230
rect 45 176 75 214
rect 45 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 311 176 346 265
rect 618 251 668 281
rect 755 315 836 325
rect 755 281 771 315
rect 805 281 836 315
rect 755 271 836 281
rect 903 279 933 413
rect 987 375 1017 413
rect 1107 381 1137 413
rect 975 365 1041 375
rect 975 331 991 365
rect 1025 331 1041 365
rect 975 321 1041 331
rect 1102 365 1171 381
rect 1102 331 1127 365
rect 1161 331 1171 365
rect 1102 315 1171 331
rect 418 214 479 230
rect 418 180 429 214
rect 463 180 479 214
rect 418 177 479 180
rect 618 177 648 251
rect 311 174 362 176
rect 419 175 648 177
rect 311 172 366 174
rect 420 173 648 175
rect 311 170 369 172
rect 421 170 648 173
rect 311 169 371 170
rect 311 167 373 169
rect 422 167 648 170
rect 311 164 375 167
rect 311 161 377 164
rect 311 157 379 161
rect 311 146 381 157
rect 351 131 381 146
rect 423 147 648 167
rect 696 203 750 219
rect 696 169 706 203
rect 740 169 750 203
rect 696 153 750 169
rect 423 131 453 147
rect 618 131 648 147
rect 705 131 735 153
rect 792 131 822 271
rect 903 249 1041 279
rect 1000 219 1041 249
rect 887 191 958 207
rect 887 157 914 191
rect 948 157 958 191
rect 887 141 958 157
rect 1000 203 1060 219
rect 1000 169 1016 203
rect 1050 169 1060 203
rect 1000 153 1060 169
rect 887 119 917 141
rect 1000 119 1030 153
rect 1102 131 1132 315
rect 1213 229 1243 413
rect 1686 381 1716 413
rect 1662 365 1716 381
rect 1770 375 1800 413
rect 1888 381 1918 413
rect 1662 331 1672 365
rect 1706 331 1716 365
rect 1321 297 1351 329
rect 1285 281 1351 297
rect 1285 247 1295 281
rect 1329 273 1351 281
rect 1405 297 1435 329
rect 1405 281 1491 297
rect 1329 247 1342 273
rect 1405 257 1447 281
rect 1285 231 1342 247
rect 1174 213 1243 229
rect 1174 179 1190 213
rect 1224 179 1241 213
rect 1174 163 1241 179
rect 1312 175 1342 231
rect 1396 247 1447 257
rect 1481 247 1491 281
rect 1396 231 1491 247
rect 1542 263 1572 329
rect 1662 315 1716 331
rect 1758 365 1824 375
rect 1758 331 1774 365
rect 1808 331 1824 365
rect 1758 321 1824 331
rect 1887 365 1954 381
rect 1887 331 1910 365
rect 1944 331 1954 365
rect 1686 279 1716 315
rect 1887 315 1954 331
rect 1542 247 1619 263
rect 1686 249 1822 279
rect 1542 233 1575 247
rect 1396 175 1426 231
rect 1565 213 1575 233
rect 1609 213 1619 247
rect 1565 197 1619 213
rect 1584 175 1614 197
rect 1684 191 1750 207
rect 1211 131 1241 163
rect 1684 157 1706 191
rect 1740 157 1750 191
rect 1684 141 1750 157
rect 1684 119 1714 141
rect 1792 119 1822 249
rect 1887 131 1917 315
rect 1996 229 2026 413
rect 2363 429 2393 455
rect 2092 281 2122 329
rect 1959 213 2026 229
rect 2068 265 2122 281
rect 2164 297 2194 329
rect 2164 281 2260 297
rect 2164 267 2216 281
rect 2068 231 2078 265
rect 2112 231 2122 265
rect 2068 215 2122 231
rect 2175 247 2216 267
rect 2250 247 2260 281
rect 2363 269 2393 301
rect 2648 481 2678 507
rect 2743 497 2773 523
rect 2648 337 2678 353
rect 2623 307 2678 337
rect 2175 231 2260 247
rect 2313 253 2393 269
rect 2460 265 2490 297
rect 1959 179 1969 213
rect 2003 179 2026 213
rect 1959 163 2026 179
rect 2091 175 2121 215
rect 2175 175 2205 231
rect 2313 219 2323 253
rect 2357 219 2393 253
rect 2313 203 2393 219
rect 1974 131 2004 163
rect 2363 131 2393 203
rect 2441 259 2490 265
rect 2623 259 2653 307
rect 2743 265 2773 297
rect 2441 249 2653 259
rect 2441 215 2451 249
rect 2485 215 2653 249
rect 2441 205 2653 215
rect 2441 199 2490 205
rect 2460 177 2490 199
rect 2623 176 2653 205
rect 2715 249 2773 265
rect 2715 215 2725 249
rect 2759 215 2773 249
rect 2715 199 2773 215
rect 2743 177 2773 199
rect 2623 146 2678 176
rect 2648 131 2678 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 423 21 453 47
rect 618 21 648 47
rect 705 21 735 47
rect 792 21 822 47
rect 887 21 917 47
rect 1000 21 1030 47
rect 1102 21 1132 47
rect 1211 21 1241 47
rect 1312 21 1342 47
rect 1396 21 1426 47
rect 1584 21 1614 47
rect 1684 21 1714 47
rect 1792 21 1822 47
rect 1887 21 1917 47
rect 1974 21 2004 47
rect 2091 21 2121 47
rect 2175 21 2205 47
rect 2363 21 2393 47
rect 2460 21 2490 47
rect 2648 21 2678 47
rect 2743 21 2773 47
<< polycont >>
rect 31 230 65 264
rect 552 331 586 365
rect 305 281 339 315
rect 133 230 167 264
rect 771 281 805 315
rect 991 331 1025 365
rect 1127 331 1161 365
rect 429 180 463 214
rect 706 169 740 203
rect 914 157 948 191
rect 1016 169 1050 203
rect 1672 331 1706 365
rect 1295 247 1329 281
rect 1190 179 1224 213
rect 1447 247 1481 281
rect 1774 331 1808 365
rect 1910 331 1944 365
rect 1575 213 1609 247
rect 1706 157 1740 191
rect 2078 231 2112 265
rect 2216 247 2250 281
rect 1969 179 2003 213
rect 2323 219 2357 253
rect 2451 215 2485 249
rect 2725 215 2759 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 19 477 69 493
rect 19 443 35 477
rect 19 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 247 493
rect 237 443 247 477
rect 19 375 35 409
rect 203 409 247 443
rect 69 375 167 393
rect 19 359 167 375
rect 17 264 87 325
rect 17 230 31 264
rect 65 230 87 264
rect 17 195 87 230
rect 121 264 167 359
rect 121 230 133 264
rect 121 187 167 230
rect 19 153 121 161
rect 155 153 167 187
rect 19 127 167 153
rect 237 391 247 409
rect 286 479 357 527
rect 286 445 307 479
rect 341 445 357 479
rect 594 477 628 493
rect 286 411 357 445
rect 286 377 307 411
rect 341 377 357 411
rect 443 443 463 477
rect 497 443 515 477
rect 443 409 515 443
rect 443 375 463 409
rect 497 375 515 409
rect 662 477 728 527
rect 662 443 678 477
rect 712 443 728 477
rect 846 477 889 493
rect 594 381 628 443
rect 203 357 213 375
rect 19 119 69 127
rect 19 85 35 119
rect 203 119 247 357
rect 283 315 339 337
rect 283 281 305 315
rect 283 205 339 281
rect 387 230 431 339
rect 481 301 515 375
rect 552 365 628 381
rect 586 349 628 365
rect 586 331 721 349
rect 765 335 812 475
rect 880 443 889 477
rect 927 450 943 484
rect 977 450 1093 484
rect 846 427 889 443
rect 552 315 721 331
rect 481 293 521 301
rect 481 286 526 293
rect 481 281 534 286
rect 481 259 615 281
rect 492 255 615 259
rect 492 251 581 255
rect 387 214 463 230
rect 387 180 429 214
rect 387 163 463 180
rect 497 221 581 251
rect 497 215 615 221
rect 686 219 721 315
rect 755 315 812 335
rect 755 281 771 315
rect 805 281 821 315
rect 855 261 889 427
rect 849 255 889 261
rect 845 247 846 255
rect 790 221 846 247
rect 880 235 889 255
rect 923 357 949 391
rect 983 365 1025 391
rect 983 357 991 365
rect 923 331 991 357
rect 923 315 1025 331
rect 880 221 882 235
rect 19 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 247 119
rect 203 69 247 85
rect 286 111 341 127
rect 286 77 307 111
rect 103 17 169 59
rect 286 17 341 77
rect 387 69 431 163
rect 497 119 531 215
rect 686 203 754 219
rect 686 169 706 203
rect 740 169 754 203
rect 686 159 754 169
rect 465 103 531 119
rect 465 69 470 103
rect 504 69 531 103
rect 465 53 531 69
rect 574 153 754 159
rect 790 213 880 221
rect 574 125 729 153
rect 574 111 608 125
rect 790 119 824 213
rect 923 207 958 315
rect 1059 281 1093 450
rect 1141 475 1217 527
rect 1435 485 1501 527
rect 1141 441 1157 475
rect 1191 441 1217 475
rect 1277 459 1311 475
rect 1277 407 1311 425
rect 1435 451 1451 485
rect 1485 451 1501 485
rect 1924 485 2000 527
rect 1435 417 1501 451
rect 1710 450 1726 484
rect 1760 450 1876 484
rect 1924 451 1940 485
rect 1974 451 2000 485
rect 2188 485 2466 527
rect 2048 459 2082 475
rect 1127 391 1397 407
rect 1127 365 1277 391
rect 1161 357 1277 365
rect 1311 357 1397 391
rect 1435 383 1451 417
rect 1485 383 1501 417
rect 1672 391 1719 397
rect 1161 331 1177 357
rect 1127 315 1177 331
rect 1279 281 1329 297
rect 1059 247 1295 281
rect 1059 239 1134 247
rect 914 191 958 207
rect 948 157 958 191
rect 914 141 958 157
rect 1000 169 1016 203
rect 1050 187 1066 203
rect 1000 153 1031 169
rect 1065 153 1066 187
rect 1000 147 1066 153
rect 1100 131 1134 239
rect 1285 231 1329 247
rect 1363 213 1397 357
rect 1672 365 1685 391
rect 1706 331 1719 357
rect 1431 323 1632 331
rect 1431 289 1593 323
rect 1627 289 1632 323
rect 1672 315 1719 331
rect 1767 365 1808 381
rect 1767 331 1774 365
rect 1431 283 1632 289
rect 1431 281 1497 283
rect 1431 247 1447 281
rect 1481 247 1497 281
rect 1767 261 1808 331
rect 1684 255 1808 261
rect 1559 213 1575 247
rect 1609 213 1625 247
rect 1174 179 1190 213
rect 1224 193 1243 213
rect 1363 212 1625 213
rect 1224 187 1259 193
rect 1224 179 1225 187
rect 1174 153 1225 179
rect 1362 179 1625 212
rect 1684 221 1685 255
rect 1719 225 1808 255
rect 1842 281 1876 450
rect 2188 451 2204 485
rect 2238 451 2416 485
rect 2450 451 2466 485
rect 2048 417 2082 425
rect 2500 448 2557 493
rect 1910 383 2466 417
rect 1910 365 1960 383
rect 1944 331 1960 365
rect 1910 315 1960 331
rect 1842 265 2112 281
rect 1842 247 2078 265
rect 1719 221 1741 225
rect 1684 191 1741 221
rect 1362 156 1402 179
rect 1174 147 1259 153
rect 790 103 866 119
rect 574 61 608 77
rect 645 55 661 89
rect 695 55 711 89
rect 790 85 832 103
rect 645 17 711 55
rect 1097 117 1134 131
rect 1336 122 1352 156
rect 1386 122 1402 156
rect 1684 157 1706 191
rect 1740 157 1741 191
rect 1436 127 1470 143
rect 1684 141 1741 157
rect 1097 93 1131 117
rect 832 53 866 69
rect 911 59 927 93
rect 961 59 1131 93
rect 911 53 1131 59
rect 1167 89 1201 105
rect 1842 93 1876 247
rect 2068 231 2078 247
rect 2068 215 2112 231
rect 1951 187 1969 213
rect 1951 153 1961 187
rect 2003 179 2026 213
rect 1995 153 2026 179
rect 2146 156 2181 383
rect 1951 147 2026 153
rect 2115 153 2181 156
rect 2115 119 2131 153
rect 2165 119 2181 153
rect 2216 323 2319 349
rect 2216 289 2237 323
rect 2271 315 2319 323
rect 2353 315 2371 349
rect 2216 281 2271 289
rect 2250 247 2271 281
rect 2432 265 2466 383
rect 2534 414 2557 448
rect 2500 380 2557 414
rect 2534 346 2557 380
rect 2500 326 2557 346
rect 2216 185 2271 247
rect 2307 253 2398 265
rect 2307 219 2323 253
rect 2357 219 2398 253
rect 2432 249 2485 265
rect 2432 215 2451 249
rect 2432 199 2485 215
rect 2216 151 2355 185
rect 1167 17 1201 55
rect 1252 59 1268 93
rect 1302 85 1318 93
rect 1436 85 1470 93
rect 1302 59 1470 85
rect 1252 51 1470 59
rect 1524 59 1540 93
rect 1574 59 1595 93
rect 1524 17 1595 59
rect 1723 59 1739 93
rect 1773 59 1876 93
rect 1723 53 1876 59
rect 1912 89 1964 105
rect 1912 55 1930 89
rect 1912 17 1964 55
rect 2016 75 2032 109
rect 2066 85 2082 109
rect 2215 101 2250 117
rect 2066 75 2215 85
rect 2016 67 2215 75
rect 2249 67 2250 101
rect 2016 51 2250 67
rect 2313 103 2355 151
rect 2313 69 2319 103
rect 2353 69 2355 103
rect 2313 53 2355 69
rect 2400 127 2416 161
rect 2450 127 2466 161
rect 2521 143 2557 326
rect 2400 93 2466 127
rect 2400 59 2416 93
rect 2450 59 2466 93
rect 2400 17 2466 59
rect 2500 127 2557 143
rect 2534 93 2557 127
rect 2500 51 2557 93
rect 2592 467 2655 483
rect 2592 433 2604 467
rect 2638 433 2655 467
rect 2592 399 2655 433
rect 2592 365 2604 399
rect 2638 365 2655 399
rect 2592 265 2655 365
rect 2691 473 2748 527
rect 2691 439 2699 473
rect 2733 439 2748 473
rect 2691 405 2748 439
rect 2691 371 2698 405
rect 2732 371 2748 405
rect 2691 353 2748 371
rect 2783 449 2835 493
rect 2817 415 2835 449
rect 2783 381 2835 415
rect 2817 347 2835 381
rect 2783 294 2835 347
rect 2592 249 2759 265
rect 2592 215 2725 249
rect 2592 199 2759 215
rect 2592 119 2655 199
rect 2793 157 2835 294
rect 2592 85 2604 119
rect 2638 85 2655 119
rect 2783 129 2835 157
rect 2592 51 2655 85
rect 2691 93 2749 109
rect 2691 59 2699 93
rect 2733 59 2749 93
rect 2691 17 2749 59
rect 2817 95 2835 129
rect 2783 51 2835 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 121 153 155 187
rect 213 375 237 391
rect 237 375 247 391
rect 213 357 247 375
rect 581 221 615 255
rect 846 221 880 255
rect 949 357 983 391
rect 1031 169 1050 187
rect 1050 169 1065 187
rect 1031 153 1065 169
rect 1685 365 1719 391
rect 1685 357 1706 365
rect 1706 357 1719 365
rect 1593 289 1627 323
rect 1225 153 1259 187
rect 1685 221 1719 255
rect 1961 179 1969 187
rect 1969 179 1995 187
rect 1961 153 1995 179
rect 2237 289 2271 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 937 391 995 397
rect 937 388 949 391
rect 247 360 949 388
rect 247 357 259 360
rect 201 351 259 357
rect 937 357 949 360
rect 983 388 995 391
rect 1673 391 1731 397
rect 1673 388 1685 391
rect 983 360 1685 388
rect 983 357 995 360
rect 937 351 995 357
rect 1673 357 1685 360
rect 1719 357 1731 391
rect 1673 351 1731 357
rect 1581 323 1639 329
rect 1581 289 1593 323
rect 1627 320 1639 323
rect 2225 323 2283 329
rect 2225 320 2237 323
rect 1627 292 2237 320
rect 1627 289 1639 292
rect 1581 283 1639 289
rect 2225 289 2237 292
rect 2271 289 2283 323
rect 2225 283 2283 289
rect 569 255 627 261
rect 569 221 581 255
rect 615 252 627 255
rect 834 255 892 261
rect 834 252 846 255
rect 615 224 846 252
rect 615 221 627 224
rect 569 215 627 221
rect 834 221 846 224
rect 880 221 892 255
rect 1673 255 1731 261
rect 1673 252 1685 255
rect 834 215 892 221
rect 1034 224 1685 252
rect 1034 193 1077 224
rect 1673 221 1685 224
rect 1719 221 1731 255
rect 1673 215 1731 221
rect 109 187 167 193
rect 109 153 121 187
rect 155 184 167 187
rect 1019 187 1077 193
rect 1019 184 1031 187
rect 155 156 1031 184
rect 155 153 167 156
rect 109 147 167 153
rect 1019 153 1031 156
rect 1065 153 1077 187
rect 1019 147 1077 153
rect 1213 187 1271 193
rect 1213 153 1225 187
rect 1259 184 1271 187
rect 1949 187 2007 193
rect 1949 184 1961 187
rect 1259 156 1961 184
rect 1259 153 1271 156
rect 1213 147 1271 153
rect 1949 153 1961 156
rect 1995 153 2007 187
rect 1949 147 2007 153
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< labels >>
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 SCD
port 4 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 SCD
port 4 nsew signal input
flabel locali s 397 289 431 323 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel locali s 397 85 431 119 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel locali s 2329 221 2363 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 1225 153 1259 187 0 FreeSans 400 0 0 0 SET_B
port 6 nsew signal input
flabel locali s 2789 85 2823 119 0 FreeSans 400 0 0 0 Q
port 11 nsew signal output
flabel locali s 2789 357 2823 391 0 FreeSans 400 0 0 0 Q
port 11 nsew signal output
flabel locali s 2789 425 2823 459 0 FreeSans 400 0 0 0 Q
port 11 nsew signal output
flabel locali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel locali s 765 289 799 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 765 425 799 459 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2513 425 2547 459 0 FreeSans 400 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2513 357 2547 391 0 FreeSans 400 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2513 85 2547 119 0 FreeSans 400 0 0 0 Q_N
port 12 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 3 FreeSans 400 0 0 0 VPB
port 9 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel pwell s 29 -17 63 17 3 FreeSans 400 0 0 0 VNB
port 8 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfbbn_1
rlabel locali s 1951 147 2026 213 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1949 184 2007 193 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1949 147 2007 156 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 184 1271 193 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 156 2007 184 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 147 1271 156 1 SET_B
port 6 nsew signal input
rlabel metal1 s 0 -48 2852 48 1 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2852 592 1 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2852 544
string GDS_END 241634
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 218692
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
