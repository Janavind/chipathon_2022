magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< pwell >>
rect -26 -26 824 362
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
rect 384 0 414 336
rect 492 0 522 336
rect 600 0 630 336
rect 708 0 738 336
<< ndiff >>
rect 0 185 60 336
rect 0 151 8 185
rect 42 151 60 185
rect 0 0 60 151
rect 90 185 168 336
rect 90 151 112 185
rect 146 151 168 185
rect 90 0 168 151
rect 198 185 276 336
rect 198 151 220 185
rect 254 151 276 185
rect 198 0 276 151
rect 306 185 384 336
rect 306 151 328 185
rect 362 151 384 185
rect 306 0 384 151
rect 414 185 492 336
rect 414 151 436 185
rect 470 151 492 185
rect 414 0 492 151
rect 522 185 600 336
rect 522 151 544 185
rect 578 151 600 185
rect 522 0 600 151
rect 630 185 708 336
rect 630 151 652 185
rect 686 151 708 185
rect 630 0 708 151
rect 738 185 798 336
rect 738 151 756 185
rect 790 151 798 185
rect 738 0 798 151
<< ndiffc >>
rect 8 151 42 185
rect 112 151 146 185
rect 220 151 254 185
rect 328 151 362 185
rect 436 151 470 185
rect 544 151 578 185
rect 652 151 686 185
rect 756 151 790 185
<< poly >>
rect 60 362 738 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 384 336 414 362
rect 492 336 522 362
rect 600 336 630 362
rect 708 336 738 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
<< locali >>
rect 112 235 790 269
rect 8 185 42 201
rect 8 135 42 151
rect 112 185 146 235
rect 112 135 146 151
rect 220 185 254 201
rect 220 135 254 151
rect 328 185 362 235
rect 328 135 362 151
rect 436 185 470 201
rect 436 135 470 151
rect 544 185 578 235
rect 544 135 578 151
rect 652 185 686 201
rect 652 135 686 151
rect 756 185 790 235
rect 756 135 790 151
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_0
timestamp 1666199351
transform 1 0 748 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_1
timestamp 1666199351
transform 1 0 644 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_2
timestamp 1666199351
transform 1 0 536 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_3
timestamp 1666199351
transform 1 0 428 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_4
timestamp 1666199351
transform 1 0 320 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_5
timestamp 1666199351
transform 1 0 212 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_6
timestamp 1666199351
transform 1 0 104 0 1 135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_7
timestamp 1666199351
transform 1 0 0 0 1 135
box 0 0 1 1
<< labels >>
rlabel locali s 669 168 669 168 4 S
port 1 nsew
rlabel locali s 25 168 25 168 4 S
port 1 nsew
rlabel locali s 237 168 237 168 4 S
port 1 nsew
rlabel locali s 453 168 453 168 4 S
port 1 nsew
rlabel locali s 451 252 451 252 4 D
port 2 nsew
rlabel poly s 399 377 399 377 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -25 -26 823 392
string GDS_END 37750
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 35546
<< end >>
