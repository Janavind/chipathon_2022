magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect 7295 4707 8101 6839
rect 7445 2944 8095 4476
rect 17560 4144 19398 4322
rect 12748 3038 20068 4144
rect 12748 3012 19938 3038
rect 15236 2962 16666 3012
rect 20028 3012 20068 3038
<< pwell >>
rect 12094 4883 12372 5599
rect 12094 4863 13432 4883
rect 11434 4605 13432 4863
rect 11502 4537 13432 4605
rect 11502 4285 13508 4537
rect 12408 3146 12688 4104
rect 19938 2861 20028 3038
<< mvnmos >>
rect 11460 4684 12060 4784
rect 12173 4573 12293 5573
rect 12406 4684 13406 4804
rect 11581 4311 11781 4511
rect 11837 4311 12037 4511
rect 12093 4311 12293 4511
rect 12349 4311 12549 4511
rect 12605 4311 12725 4511
rect 12781 4311 12901 4511
rect 12957 4311 13077 4511
rect 13133 4311 13253 4511
rect 13309 4311 13429 4511
rect 12434 3225 12518 4025
rect 12578 3225 12662 4025
<< mvpmos >>
rect 7414 4773 7514 6773
rect 7570 4773 7670 6773
rect 7726 4773 7826 6773
rect 7882 4773 7982 6773
rect 7564 3010 7664 4410
rect 7720 3010 7820 4410
rect 7876 3010 7976 4410
rect 17679 4172 19279 4256
rect 12906 3225 12990 4025
rect 13247 3873 13347 4073
rect 13403 3873 13503 4073
rect 13755 3078 13855 4078
rect 13911 3078 14011 4078
rect 14067 3078 14167 4078
rect 14223 3078 14323 4078
rect 14379 3078 14479 4078
rect 14535 3078 14635 4078
rect 14691 3078 14791 4078
rect 14847 3078 14947 4078
rect 15003 3078 15103 4078
rect 15355 3028 15455 4028
rect 15511 3028 15611 4028
rect 15667 3028 15767 4028
rect 15823 3028 15923 4028
rect 15979 3028 16079 4028
rect 16135 3028 16235 4028
rect 16291 3028 16391 4028
rect 16447 3028 16547 4028
rect 16799 3078 16899 4078
rect 16955 3078 17055 4078
rect 17111 3078 17211 4078
rect 17267 3078 17367 4078
rect 17423 3078 17523 4078
rect 17579 3078 17679 4078
rect 17735 3078 17835 4078
rect 17891 3078 17991 4078
rect 18243 3078 18343 4078
rect 18399 3078 18499 4078
rect 18555 3078 18655 4078
rect 18711 3078 18811 4078
rect 18867 3078 18967 4078
rect 19023 3078 19123 4078
rect 19179 3078 19279 4078
rect 19335 3078 19435 4078
rect 19601 3078 19701 4078
rect 19757 3078 19857 4078
<< mvndiff >>
rect 12120 5503 12173 5573
rect 12120 5469 12128 5503
rect 12162 5469 12173 5503
rect 12120 5435 12173 5469
rect 12120 5401 12128 5435
rect 12162 5401 12173 5435
rect 12120 5367 12173 5401
rect 12120 5333 12128 5367
rect 12162 5333 12173 5367
rect 12120 5299 12173 5333
rect 12120 5265 12128 5299
rect 12162 5265 12173 5299
rect 12120 5231 12173 5265
rect 12120 5197 12128 5231
rect 12162 5197 12173 5231
rect 12120 5163 12173 5197
rect 12120 5129 12128 5163
rect 12162 5129 12173 5163
rect 12120 5095 12173 5129
rect 12120 5061 12128 5095
rect 12162 5061 12173 5095
rect 12120 5027 12173 5061
rect 12120 4993 12128 5027
rect 12162 4993 12173 5027
rect 12120 4959 12173 4993
rect 12120 4925 12128 4959
rect 12162 4925 12173 4959
rect 12120 4891 12173 4925
rect 12120 4857 12128 4891
rect 12162 4857 12173 4891
rect 11460 4829 12060 4837
rect 11460 4795 11538 4829
rect 11572 4795 11606 4829
rect 11640 4795 11674 4829
rect 11708 4795 11742 4829
rect 11776 4795 11810 4829
rect 11844 4795 11878 4829
rect 11912 4795 11946 4829
rect 11980 4795 12014 4829
rect 12048 4795 12060 4829
rect 11460 4784 12060 4795
rect 12120 4823 12173 4857
rect 12120 4789 12128 4823
rect 12162 4789 12173 4823
rect 12120 4755 12173 4789
rect 12120 4721 12128 4755
rect 12162 4721 12173 4755
rect 12120 4687 12173 4721
rect 11460 4673 12060 4684
rect 11460 4639 11538 4673
rect 11572 4639 11606 4673
rect 11640 4639 11674 4673
rect 11708 4639 11742 4673
rect 11776 4639 11810 4673
rect 11844 4639 11878 4673
rect 11912 4639 11946 4673
rect 11980 4639 12014 4673
rect 12048 4639 12060 4673
rect 11460 4631 12060 4639
rect 12120 4653 12128 4687
rect 12162 4653 12173 4687
rect 12120 4619 12173 4653
rect 12120 4585 12128 4619
rect 12162 4585 12173 4619
rect 12120 4573 12173 4585
rect 12293 5503 12346 5573
rect 12293 5469 12304 5503
rect 12338 5469 12346 5503
rect 12293 5435 12346 5469
rect 12293 5401 12304 5435
rect 12338 5401 12346 5435
rect 12293 5367 12346 5401
rect 12293 5333 12304 5367
rect 12338 5333 12346 5367
rect 12293 5299 12346 5333
rect 12293 5265 12304 5299
rect 12338 5265 12346 5299
rect 12293 5231 12346 5265
rect 12293 5197 12304 5231
rect 12338 5197 12346 5231
rect 12293 5163 12346 5197
rect 12293 5129 12304 5163
rect 12338 5129 12346 5163
rect 12293 5095 12346 5129
rect 12293 5061 12304 5095
rect 12338 5061 12346 5095
rect 12293 5027 12346 5061
rect 12293 4993 12304 5027
rect 12338 4993 12346 5027
rect 12293 4959 12346 4993
rect 12293 4925 12304 4959
rect 12338 4925 12346 4959
rect 12293 4891 12346 4925
rect 12293 4857 12304 4891
rect 12338 4857 12346 4891
rect 12293 4823 12346 4857
rect 12293 4789 12304 4823
rect 12338 4789 12346 4823
rect 12406 4849 13406 4857
rect 12406 4815 12418 4849
rect 12452 4815 12486 4849
rect 12520 4815 12554 4849
rect 12588 4815 12622 4849
rect 12656 4815 12690 4849
rect 12724 4815 12758 4849
rect 12792 4815 12826 4849
rect 12860 4815 12894 4849
rect 12928 4815 12962 4849
rect 12996 4815 13030 4849
rect 13064 4815 13098 4849
rect 13132 4815 13166 4849
rect 13200 4815 13234 4849
rect 13268 4815 13302 4849
rect 13336 4815 13406 4849
rect 12406 4804 13406 4815
rect 12293 4755 12346 4789
rect 12293 4721 12304 4755
rect 12338 4721 12346 4755
rect 12293 4687 12346 4721
rect 12293 4653 12304 4687
rect 12338 4653 12346 4687
rect 12293 4619 12346 4653
rect 12406 4673 13406 4684
rect 12406 4639 12418 4673
rect 12452 4639 12486 4673
rect 12520 4639 12554 4673
rect 12588 4639 12622 4673
rect 12656 4639 12690 4673
rect 12724 4639 12758 4673
rect 12792 4639 12826 4673
rect 12860 4639 12894 4673
rect 12928 4639 12962 4673
rect 12996 4639 13030 4673
rect 13064 4639 13098 4673
rect 13132 4639 13166 4673
rect 13200 4639 13234 4673
rect 13268 4639 13302 4673
rect 13336 4639 13406 4673
rect 12406 4631 13406 4639
rect 12293 4585 12304 4619
rect 12338 4585 12346 4619
rect 12293 4573 12346 4585
rect 11528 4493 11581 4511
rect 11528 4459 11536 4493
rect 11570 4459 11581 4493
rect 11528 4425 11581 4459
rect 11528 4391 11536 4425
rect 11570 4391 11581 4425
rect 11528 4357 11581 4391
rect 11528 4323 11536 4357
rect 11570 4323 11581 4357
rect 11528 4311 11581 4323
rect 11781 4493 11837 4511
rect 11781 4459 11792 4493
rect 11826 4459 11837 4493
rect 11781 4425 11837 4459
rect 11781 4391 11792 4425
rect 11826 4391 11837 4425
rect 11781 4357 11837 4391
rect 11781 4323 11792 4357
rect 11826 4323 11837 4357
rect 11781 4311 11837 4323
rect 12037 4493 12093 4511
rect 12037 4459 12048 4493
rect 12082 4459 12093 4493
rect 12037 4425 12093 4459
rect 12037 4391 12048 4425
rect 12082 4391 12093 4425
rect 12037 4357 12093 4391
rect 12037 4323 12048 4357
rect 12082 4323 12093 4357
rect 12037 4311 12093 4323
rect 12293 4493 12349 4511
rect 12293 4459 12304 4493
rect 12338 4459 12349 4493
rect 12293 4425 12349 4459
rect 12293 4391 12304 4425
rect 12338 4391 12349 4425
rect 12293 4357 12349 4391
rect 12293 4323 12304 4357
rect 12338 4323 12349 4357
rect 12293 4311 12349 4323
rect 12549 4493 12605 4511
rect 12549 4459 12560 4493
rect 12594 4459 12605 4493
rect 12549 4425 12605 4459
rect 12549 4391 12560 4425
rect 12594 4391 12605 4425
rect 12549 4357 12605 4391
rect 12549 4323 12560 4357
rect 12594 4323 12605 4357
rect 12549 4311 12605 4323
rect 12725 4493 12781 4511
rect 12725 4459 12736 4493
rect 12770 4459 12781 4493
rect 12725 4425 12781 4459
rect 12725 4391 12736 4425
rect 12770 4391 12781 4425
rect 12725 4357 12781 4391
rect 12725 4323 12736 4357
rect 12770 4323 12781 4357
rect 12725 4311 12781 4323
rect 12901 4493 12957 4511
rect 12901 4459 12912 4493
rect 12946 4459 12957 4493
rect 12901 4425 12957 4459
rect 12901 4391 12912 4425
rect 12946 4391 12957 4425
rect 12901 4357 12957 4391
rect 12901 4323 12912 4357
rect 12946 4323 12957 4357
rect 12901 4311 12957 4323
rect 13077 4493 13133 4511
rect 13077 4459 13088 4493
rect 13122 4459 13133 4493
rect 13077 4425 13133 4459
rect 13077 4391 13088 4425
rect 13122 4391 13133 4425
rect 13077 4357 13133 4391
rect 13077 4323 13088 4357
rect 13122 4323 13133 4357
rect 13077 4311 13133 4323
rect 13253 4493 13309 4511
rect 13253 4459 13264 4493
rect 13298 4459 13309 4493
rect 13253 4425 13309 4459
rect 13253 4391 13264 4425
rect 13298 4391 13309 4425
rect 13253 4357 13309 4391
rect 13253 4323 13264 4357
rect 13298 4323 13309 4357
rect 13253 4311 13309 4323
rect 13429 4493 13482 4511
rect 13429 4459 13440 4493
rect 13474 4459 13482 4493
rect 13429 4425 13482 4459
rect 13429 4391 13440 4425
rect 13474 4391 13482 4425
rect 13429 4357 13482 4391
rect 13429 4323 13440 4357
rect 13474 4323 13482 4357
rect 13429 4311 13482 4323
rect 12434 4070 12518 4078
rect 12434 4036 12472 4070
rect 12506 4036 12518 4070
rect 12434 4025 12518 4036
rect 12578 4070 12662 4078
rect 12578 4036 12616 4070
rect 12650 4036 12662 4070
rect 12578 4025 12662 4036
rect 12434 3214 12518 3225
rect 12434 3180 12472 3214
rect 12506 3180 12518 3214
rect 12434 3172 12518 3180
rect 12578 3214 12662 3225
rect 12578 3180 12616 3214
rect 12650 3180 12662 3214
rect 12578 3172 12662 3180
<< mvpdiff >>
rect 7361 6723 7414 6773
rect 7361 6689 7369 6723
rect 7403 6689 7414 6723
rect 7361 6655 7414 6689
rect 7361 6621 7369 6655
rect 7403 6621 7414 6655
rect 7361 6587 7414 6621
rect 7361 6553 7369 6587
rect 7403 6553 7414 6587
rect 7361 6519 7414 6553
rect 7361 6485 7369 6519
rect 7403 6485 7414 6519
rect 7361 6451 7414 6485
rect 7361 6417 7369 6451
rect 7403 6417 7414 6451
rect 7361 6383 7414 6417
rect 7361 6349 7369 6383
rect 7403 6349 7414 6383
rect 7361 6315 7414 6349
rect 7361 6281 7369 6315
rect 7403 6281 7414 6315
rect 7361 6247 7414 6281
rect 7361 6213 7369 6247
rect 7403 6213 7414 6247
rect 7361 6179 7414 6213
rect 7361 6145 7369 6179
rect 7403 6145 7414 6179
rect 7361 6111 7414 6145
rect 7361 6077 7369 6111
rect 7403 6077 7414 6111
rect 7361 6043 7414 6077
rect 7361 6009 7369 6043
rect 7403 6009 7414 6043
rect 7361 5975 7414 6009
rect 7361 5941 7369 5975
rect 7403 5941 7414 5975
rect 7361 5907 7414 5941
rect 7361 5873 7369 5907
rect 7403 5873 7414 5907
rect 7361 5839 7414 5873
rect 7361 5805 7369 5839
rect 7403 5805 7414 5839
rect 7361 5771 7414 5805
rect 7361 5737 7369 5771
rect 7403 5737 7414 5771
rect 7361 5703 7414 5737
rect 7361 5669 7369 5703
rect 7403 5669 7414 5703
rect 7361 5635 7414 5669
rect 7361 5601 7369 5635
rect 7403 5601 7414 5635
rect 7361 5567 7414 5601
rect 7361 5533 7369 5567
rect 7403 5533 7414 5567
rect 7361 5499 7414 5533
rect 7361 5465 7369 5499
rect 7403 5465 7414 5499
rect 7361 5431 7414 5465
rect 7361 5397 7369 5431
rect 7403 5397 7414 5431
rect 7361 5363 7414 5397
rect 7361 5329 7369 5363
rect 7403 5329 7414 5363
rect 7361 5295 7414 5329
rect 7361 5261 7369 5295
rect 7403 5261 7414 5295
rect 7361 5227 7414 5261
rect 7361 5193 7369 5227
rect 7403 5193 7414 5227
rect 7361 5159 7414 5193
rect 7361 5125 7369 5159
rect 7403 5125 7414 5159
rect 7361 5091 7414 5125
rect 7361 5057 7369 5091
rect 7403 5057 7414 5091
rect 7361 5023 7414 5057
rect 7361 4989 7369 5023
rect 7403 4989 7414 5023
rect 7361 4955 7414 4989
rect 7361 4921 7369 4955
rect 7403 4921 7414 4955
rect 7361 4887 7414 4921
rect 7361 4853 7369 4887
rect 7403 4853 7414 4887
rect 7361 4819 7414 4853
rect 7361 4785 7369 4819
rect 7403 4785 7414 4819
rect 7361 4773 7414 4785
rect 7514 6723 7570 6773
rect 7514 6689 7525 6723
rect 7559 6689 7570 6723
rect 7514 6655 7570 6689
rect 7514 6621 7525 6655
rect 7559 6621 7570 6655
rect 7514 6587 7570 6621
rect 7514 6553 7525 6587
rect 7559 6553 7570 6587
rect 7514 6519 7570 6553
rect 7514 6485 7525 6519
rect 7559 6485 7570 6519
rect 7514 6451 7570 6485
rect 7514 6417 7525 6451
rect 7559 6417 7570 6451
rect 7514 6383 7570 6417
rect 7514 6349 7525 6383
rect 7559 6349 7570 6383
rect 7514 6315 7570 6349
rect 7514 6281 7525 6315
rect 7559 6281 7570 6315
rect 7514 6247 7570 6281
rect 7514 6213 7525 6247
rect 7559 6213 7570 6247
rect 7514 6179 7570 6213
rect 7514 6145 7525 6179
rect 7559 6145 7570 6179
rect 7514 6111 7570 6145
rect 7514 6077 7525 6111
rect 7559 6077 7570 6111
rect 7514 6043 7570 6077
rect 7514 6009 7525 6043
rect 7559 6009 7570 6043
rect 7514 5975 7570 6009
rect 7514 5941 7525 5975
rect 7559 5941 7570 5975
rect 7514 5907 7570 5941
rect 7514 5873 7525 5907
rect 7559 5873 7570 5907
rect 7514 5839 7570 5873
rect 7514 5805 7525 5839
rect 7559 5805 7570 5839
rect 7514 5771 7570 5805
rect 7514 5737 7525 5771
rect 7559 5737 7570 5771
rect 7514 5703 7570 5737
rect 7514 5669 7525 5703
rect 7559 5669 7570 5703
rect 7514 5635 7570 5669
rect 7514 5601 7525 5635
rect 7559 5601 7570 5635
rect 7514 5567 7570 5601
rect 7514 5533 7525 5567
rect 7559 5533 7570 5567
rect 7514 5499 7570 5533
rect 7514 5465 7525 5499
rect 7559 5465 7570 5499
rect 7514 5431 7570 5465
rect 7514 5397 7525 5431
rect 7559 5397 7570 5431
rect 7514 5363 7570 5397
rect 7514 5329 7525 5363
rect 7559 5329 7570 5363
rect 7514 5295 7570 5329
rect 7514 5261 7525 5295
rect 7559 5261 7570 5295
rect 7514 5227 7570 5261
rect 7514 5193 7525 5227
rect 7559 5193 7570 5227
rect 7514 5159 7570 5193
rect 7514 5125 7525 5159
rect 7559 5125 7570 5159
rect 7514 5091 7570 5125
rect 7514 5057 7525 5091
rect 7559 5057 7570 5091
rect 7514 5023 7570 5057
rect 7514 4989 7525 5023
rect 7559 4989 7570 5023
rect 7514 4955 7570 4989
rect 7514 4921 7525 4955
rect 7559 4921 7570 4955
rect 7514 4887 7570 4921
rect 7514 4853 7525 4887
rect 7559 4853 7570 4887
rect 7514 4819 7570 4853
rect 7514 4785 7525 4819
rect 7559 4785 7570 4819
rect 7514 4773 7570 4785
rect 7670 6723 7726 6773
rect 7670 6689 7681 6723
rect 7715 6689 7726 6723
rect 7670 6655 7726 6689
rect 7670 6621 7681 6655
rect 7715 6621 7726 6655
rect 7670 6587 7726 6621
rect 7670 6553 7681 6587
rect 7715 6553 7726 6587
rect 7670 6519 7726 6553
rect 7670 6485 7681 6519
rect 7715 6485 7726 6519
rect 7670 6451 7726 6485
rect 7670 6417 7681 6451
rect 7715 6417 7726 6451
rect 7670 6383 7726 6417
rect 7670 6349 7681 6383
rect 7715 6349 7726 6383
rect 7670 6315 7726 6349
rect 7670 6281 7681 6315
rect 7715 6281 7726 6315
rect 7670 6247 7726 6281
rect 7670 6213 7681 6247
rect 7715 6213 7726 6247
rect 7670 6179 7726 6213
rect 7670 6145 7681 6179
rect 7715 6145 7726 6179
rect 7670 6111 7726 6145
rect 7670 6077 7681 6111
rect 7715 6077 7726 6111
rect 7670 6043 7726 6077
rect 7670 6009 7681 6043
rect 7715 6009 7726 6043
rect 7670 5975 7726 6009
rect 7670 5941 7681 5975
rect 7715 5941 7726 5975
rect 7670 5907 7726 5941
rect 7670 5873 7681 5907
rect 7715 5873 7726 5907
rect 7670 5839 7726 5873
rect 7670 5805 7681 5839
rect 7715 5805 7726 5839
rect 7670 5771 7726 5805
rect 7670 5737 7681 5771
rect 7715 5737 7726 5771
rect 7670 5703 7726 5737
rect 7670 5669 7681 5703
rect 7715 5669 7726 5703
rect 7670 5635 7726 5669
rect 7670 5601 7681 5635
rect 7715 5601 7726 5635
rect 7670 5567 7726 5601
rect 7670 5533 7681 5567
rect 7715 5533 7726 5567
rect 7670 5499 7726 5533
rect 7670 5465 7681 5499
rect 7715 5465 7726 5499
rect 7670 5431 7726 5465
rect 7670 5397 7681 5431
rect 7715 5397 7726 5431
rect 7670 5363 7726 5397
rect 7670 5329 7681 5363
rect 7715 5329 7726 5363
rect 7670 5295 7726 5329
rect 7670 5261 7681 5295
rect 7715 5261 7726 5295
rect 7670 5227 7726 5261
rect 7670 5193 7681 5227
rect 7715 5193 7726 5227
rect 7670 5159 7726 5193
rect 7670 5125 7681 5159
rect 7715 5125 7726 5159
rect 7670 5091 7726 5125
rect 7670 5057 7681 5091
rect 7715 5057 7726 5091
rect 7670 5023 7726 5057
rect 7670 4989 7681 5023
rect 7715 4989 7726 5023
rect 7670 4955 7726 4989
rect 7670 4921 7681 4955
rect 7715 4921 7726 4955
rect 7670 4887 7726 4921
rect 7670 4853 7681 4887
rect 7715 4853 7726 4887
rect 7670 4819 7726 4853
rect 7670 4785 7681 4819
rect 7715 4785 7726 4819
rect 7670 4773 7726 4785
rect 7826 6723 7882 6773
rect 7826 6689 7837 6723
rect 7871 6689 7882 6723
rect 7826 6655 7882 6689
rect 7826 6621 7837 6655
rect 7871 6621 7882 6655
rect 7826 6587 7882 6621
rect 7826 6553 7837 6587
rect 7871 6553 7882 6587
rect 7826 6519 7882 6553
rect 7826 6485 7837 6519
rect 7871 6485 7882 6519
rect 7826 6451 7882 6485
rect 7826 6417 7837 6451
rect 7871 6417 7882 6451
rect 7826 6383 7882 6417
rect 7826 6349 7837 6383
rect 7871 6349 7882 6383
rect 7826 6315 7882 6349
rect 7826 6281 7837 6315
rect 7871 6281 7882 6315
rect 7826 6247 7882 6281
rect 7826 6213 7837 6247
rect 7871 6213 7882 6247
rect 7826 6179 7882 6213
rect 7826 6145 7837 6179
rect 7871 6145 7882 6179
rect 7826 6111 7882 6145
rect 7826 6077 7837 6111
rect 7871 6077 7882 6111
rect 7826 6043 7882 6077
rect 7826 6009 7837 6043
rect 7871 6009 7882 6043
rect 7826 5975 7882 6009
rect 7826 5941 7837 5975
rect 7871 5941 7882 5975
rect 7826 5907 7882 5941
rect 7826 5873 7837 5907
rect 7871 5873 7882 5907
rect 7826 5839 7882 5873
rect 7826 5805 7837 5839
rect 7871 5805 7882 5839
rect 7826 5771 7882 5805
rect 7826 5737 7837 5771
rect 7871 5737 7882 5771
rect 7826 5703 7882 5737
rect 7826 5669 7837 5703
rect 7871 5669 7882 5703
rect 7826 5635 7882 5669
rect 7826 5601 7837 5635
rect 7871 5601 7882 5635
rect 7826 5567 7882 5601
rect 7826 5533 7837 5567
rect 7871 5533 7882 5567
rect 7826 5499 7882 5533
rect 7826 5465 7837 5499
rect 7871 5465 7882 5499
rect 7826 5431 7882 5465
rect 7826 5397 7837 5431
rect 7871 5397 7882 5431
rect 7826 5363 7882 5397
rect 7826 5329 7837 5363
rect 7871 5329 7882 5363
rect 7826 5295 7882 5329
rect 7826 5261 7837 5295
rect 7871 5261 7882 5295
rect 7826 5227 7882 5261
rect 7826 5193 7837 5227
rect 7871 5193 7882 5227
rect 7826 5159 7882 5193
rect 7826 5125 7837 5159
rect 7871 5125 7882 5159
rect 7826 5091 7882 5125
rect 7826 5057 7837 5091
rect 7871 5057 7882 5091
rect 7826 5023 7882 5057
rect 7826 4989 7837 5023
rect 7871 4989 7882 5023
rect 7826 4955 7882 4989
rect 7826 4921 7837 4955
rect 7871 4921 7882 4955
rect 7826 4887 7882 4921
rect 7826 4853 7837 4887
rect 7871 4853 7882 4887
rect 7826 4819 7882 4853
rect 7826 4785 7837 4819
rect 7871 4785 7882 4819
rect 7826 4773 7882 4785
rect 7982 6723 8035 6773
rect 7982 6689 7993 6723
rect 8027 6689 8035 6723
rect 7982 6655 8035 6689
rect 7982 6621 7993 6655
rect 8027 6621 8035 6655
rect 7982 6587 8035 6621
rect 7982 6553 7993 6587
rect 8027 6553 8035 6587
rect 7982 6519 8035 6553
rect 7982 6485 7993 6519
rect 8027 6485 8035 6519
rect 7982 6451 8035 6485
rect 7982 6417 7993 6451
rect 8027 6417 8035 6451
rect 7982 6383 8035 6417
rect 7982 6349 7993 6383
rect 8027 6349 8035 6383
rect 7982 6315 8035 6349
rect 7982 6281 7993 6315
rect 8027 6281 8035 6315
rect 7982 6247 8035 6281
rect 7982 6213 7993 6247
rect 8027 6213 8035 6247
rect 7982 6179 8035 6213
rect 7982 6145 7993 6179
rect 8027 6145 8035 6179
rect 7982 6111 8035 6145
rect 7982 6077 7993 6111
rect 8027 6077 8035 6111
rect 7982 6043 8035 6077
rect 7982 6009 7993 6043
rect 8027 6009 8035 6043
rect 7982 5975 8035 6009
rect 7982 5941 7993 5975
rect 8027 5941 8035 5975
rect 7982 5907 8035 5941
rect 7982 5873 7993 5907
rect 8027 5873 8035 5907
rect 7982 5839 8035 5873
rect 7982 5805 7993 5839
rect 8027 5805 8035 5839
rect 7982 5771 8035 5805
rect 7982 5737 7993 5771
rect 8027 5737 8035 5771
rect 7982 5703 8035 5737
rect 7982 5669 7993 5703
rect 8027 5669 8035 5703
rect 7982 5635 8035 5669
rect 7982 5601 7993 5635
rect 8027 5601 8035 5635
rect 7982 5567 8035 5601
rect 7982 5533 7993 5567
rect 8027 5533 8035 5567
rect 7982 5499 8035 5533
rect 7982 5465 7993 5499
rect 8027 5465 8035 5499
rect 7982 5431 8035 5465
rect 7982 5397 7993 5431
rect 8027 5397 8035 5431
rect 7982 5363 8035 5397
rect 7982 5329 7993 5363
rect 8027 5329 8035 5363
rect 7982 5295 8035 5329
rect 7982 5261 7993 5295
rect 8027 5261 8035 5295
rect 7982 5227 8035 5261
rect 7982 5193 7993 5227
rect 8027 5193 8035 5227
rect 7982 5159 8035 5193
rect 7982 5125 7993 5159
rect 8027 5125 8035 5159
rect 7982 5091 8035 5125
rect 7982 5057 7993 5091
rect 8027 5057 8035 5091
rect 7982 5023 8035 5057
rect 7982 4989 7993 5023
rect 8027 4989 8035 5023
rect 7982 4955 8035 4989
rect 7982 4921 7993 4955
rect 8027 4921 8035 4955
rect 7982 4887 8035 4921
rect 7982 4853 7993 4887
rect 8027 4853 8035 4887
rect 7982 4819 8035 4853
rect 7982 4785 7993 4819
rect 8027 4785 8035 4819
rect 7982 4773 8035 4785
rect 7511 4348 7564 4410
rect 7511 4314 7519 4348
rect 7553 4314 7564 4348
rect 7511 4280 7564 4314
rect 7511 4246 7519 4280
rect 7553 4246 7564 4280
rect 7511 4212 7564 4246
rect 7511 4178 7519 4212
rect 7553 4178 7564 4212
rect 7511 4144 7564 4178
rect 7511 4110 7519 4144
rect 7553 4110 7564 4144
rect 7511 4076 7564 4110
rect 7511 4042 7519 4076
rect 7553 4042 7564 4076
rect 7511 4008 7564 4042
rect 7511 3974 7519 4008
rect 7553 3974 7564 4008
rect 7511 3940 7564 3974
rect 7511 3906 7519 3940
rect 7553 3906 7564 3940
rect 7511 3872 7564 3906
rect 7511 3838 7519 3872
rect 7553 3838 7564 3872
rect 7511 3804 7564 3838
rect 7511 3770 7519 3804
rect 7553 3770 7564 3804
rect 7511 3736 7564 3770
rect 7511 3702 7519 3736
rect 7553 3702 7564 3736
rect 7511 3668 7564 3702
rect 7511 3634 7519 3668
rect 7553 3634 7564 3668
rect 7511 3600 7564 3634
rect 7511 3566 7519 3600
rect 7553 3566 7564 3600
rect 7511 3532 7564 3566
rect 7511 3498 7519 3532
rect 7553 3498 7564 3532
rect 7511 3464 7564 3498
rect 7511 3430 7519 3464
rect 7553 3430 7564 3464
rect 7511 3396 7564 3430
rect 7511 3362 7519 3396
rect 7553 3362 7564 3396
rect 7511 3328 7564 3362
rect 7511 3294 7519 3328
rect 7553 3294 7564 3328
rect 7511 3260 7564 3294
rect 7511 3226 7519 3260
rect 7553 3226 7564 3260
rect 7511 3192 7564 3226
rect 7511 3158 7519 3192
rect 7553 3158 7564 3192
rect 7511 3124 7564 3158
rect 7511 3090 7519 3124
rect 7553 3090 7564 3124
rect 7511 3056 7564 3090
rect 7511 3022 7519 3056
rect 7553 3022 7564 3056
rect 7511 3010 7564 3022
rect 7664 4348 7720 4410
rect 7664 4314 7675 4348
rect 7709 4314 7720 4348
rect 7664 4280 7720 4314
rect 7664 4246 7675 4280
rect 7709 4246 7720 4280
rect 7664 4212 7720 4246
rect 7664 4178 7675 4212
rect 7709 4178 7720 4212
rect 7664 4144 7720 4178
rect 7664 4110 7675 4144
rect 7709 4110 7720 4144
rect 7664 4076 7720 4110
rect 7664 4042 7675 4076
rect 7709 4042 7720 4076
rect 7664 4008 7720 4042
rect 7664 3974 7675 4008
rect 7709 3974 7720 4008
rect 7664 3940 7720 3974
rect 7664 3906 7675 3940
rect 7709 3906 7720 3940
rect 7664 3872 7720 3906
rect 7664 3838 7675 3872
rect 7709 3838 7720 3872
rect 7664 3804 7720 3838
rect 7664 3770 7675 3804
rect 7709 3770 7720 3804
rect 7664 3736 7720 3770
rect 7664 3702 7675 3736
rect 7709 3702 7720 3736
rect 7664 3668 7720 3702
rect 7664 3634 7675 3668
rect 7709 3634 7720 3668
rect 7664 3600 7720 3634
rect 7664 3566 7675 3600
rect 7709 3566 7720 3600
rect 7664 3532 7720 3566
rect 7664 3498 7675 3532
rect 7709 3498 7720 3532
rect 7664 3464 7720 3498
rect 7664 3430 7675 3464
rect 7709 3430 7720 3464
rect 7664 3396 7720 3430
rect 7664 3362 7675 3396
rect 7709 3362 7720 3396
rect 7664 3328 7720 3362
rect 7664 3294 7675 3328
rect 7709 3294 7720 3328
rect 7664 3260 7720 3294
rect 7664 3226 7675 3260
rect 7709 3226 7720 3260
rect 7664 3192 7720 3226
rect 7664 3158 7675 3192
rect 7709 3158 7720 3192
rect 7664 3124 7720 3158
rect 7664 3090 7675 3124
rect 7709 3090 7720 3124
rect 7664 3056 7720 3090
rect 7664 3022 7675 3056
rect 7709 3022 7720 3056
rect 7664 3010 7720 3022
rect 7820 4348 7876 4410
rect 7820 4314 7831 4348
rect 7865 4314 7876 4348
rect 7820 4280 7876 4314
rect 7820 4246 7831 4280
rect 7865 4246 7876 4280
rect 7820 4212 7876 4246
rect 7820 4178 7831 4212
rect 7865 4178 7876 4212
rect 7820 4144 7876 4178
rect 7820 4110 7831 4144
rect 7865 4110 7876 4144
rect 7820 4076 7876 4110
rect 7820 4042 7831 4076
rect 7865 4042 7876 4076
rect 7820 4008 7876 4042
rect 7820 3974 7831 4008
rect 7865 3974 7876 4008
rect 7820 3940 7876 3974
rect 7820 3906 7831 3940
rect 7865 3906 7876 3940
rect 7820 3872 7876 3906
rect 7820 3838 7831 3872
rect 7865 3838 7876 3872
rect 7820 3804 7876 3838
rect 7820 3770 7831 3804
rect 7865 3770 7876 3804
rect 7820 3736 7876 3770
rect 7820 3702 7831 3736
rect 7865 3702 7876 3736
rect 7820 3668 7876 3702
rect 7820 3634 7831 3668
rect 7865 3634 7876 3668
rect 7820 3600 7876 3634
rect 7820 3566 7831 3600
rect 7865 3566 7876 3600
rect 7820 3532 7876 3566
rect 7820 3498 7831 3532
rect 7865 3498 7876 3532
rect 7820 3464 7876 3498
rect 7820 3430 7831 3464
rect 7865 3430 7876 3464
rect 7820 3396 7876 3430
rect 7820 3362 7831 3396
rect 7865 3362 7876 3396
rect 7820 3328 7876 3362
rect 7820 3294 7831 3328
rect 7865 3294 7876 3328
rect 7820 3260 7876 3294
rect 7820 3226 7831 3260
rect 7865 3226 7876 3260
rect 7820 3192 7876 3226
rect 7820 3158 7831 3192
rect 7865 3158 7876 3192
rect 7820 3124 7876 3158
rect 7820 3090 7831 3124
rect 7865 3090 7876 3124
rect 7820 3056 7876 3090
rect 7820 3022 7831 3056
rect 7865 3022 7876 3056
rect 7820 3010 7876 3022
rect 7976 4348 8029 4410
rect 7976 4314 7987 4348
rect 8021 4314 8029 4348
rect 7976 4280 8029 4314
rect 7976 4246 7987 4280
rect 8021 4246 8029 4280
rect 7976 4212 8029 4246
rect 7976 4178 7987 4212
rect 8021 4178 8029 4212
rect 7976 4144 8029 4178
rect 17626 4244 17679 4256
rect 17626 4210 17634 4244
rect 17668 4210 17679 4244
rect 17626 4172 17679 4210
rect 19279 4244 19332 4256
rect 19279 4210 19290 4244
rect 19324 4210 19332 4244
rect 19279 4172 19332 4210
rect 7976 4110 7987 4144
rect 8021 4110 8029 4144
rect 7976 4076 8029 4110
rect 7976 4042 7987 4076
rect 8021 4042 8029 4076
rect 7976 4008 8029 4042
rect 7976 3974 7987 4008
rect 8021 3974 8029 4008
rect 7976 3940 8029 3974
rect 7976 3906 7987 3940
rect 8021 3906 8029 3940
rect 7976 3872 8029 3906
rect 7976 3838 7987 3872
rect 8021 3838 8029 3872
rect 7976 3804 8029 3838
rect 7976 3770 7987 3804
rect 8021 3770 8029 3804
rect 7976 3736 8029 3770
rect 7976 3702 7987 3736
rect 8021 3702 8029 3736
rect 7976 3668 8029 3702
rect 7976 3634 7987 3668
rect 8021 3634 8029 3668
rect 7976 3600 8029 3634
rect 7976 3566 7987 3600
rect 8021 3566 8029 3600
rect 7976 3532 8029 3566
rect 7976 3498 7987 3532
rect 8021 3498 8029 3532
rect 7976 3464 8029 3498
rect 7976 3430 7987 3464
rect 8021 3430 8029 3464
rect 7976 3396 8029 3430
rect 7976 3362 7987 3396
rect 8021 3362 8029 3396
rect 7976 3328 8029 3362
rect 7976 3294 7987 3328
rect 8021 3294 8029 3328
rect 7976 3260 8029 3294
rect 7976 3226 7987 3260
rect 8021 3226 8029 3260
rect 7976 3192 8029 3226
rect 12906 4070 12990 4078
rect 12906 4036 12944 4070
rect 12978 4036 12990 4070
rect 12906 4025 12990 4036
rect 13194 4061 13247 4073
rect 13194 4027 13202 4061
rect 13236 4027 13247 4061
rect 7976 3158 7987 3192
rect 8021 3158 8029 3192
rect 13194 3993 13247 4027
rect 13194 3959 13202 3993
rect 13236 3959 13247 3993
rect 13194 3925 13247 3959
rect 13194 3891 13202 3925
rect 13236 3891 13247 3925
rect 13194 3873 13247 3891
rect 13347 4061 13403 4073
rect 13347 4027 13358 4061
rect 13392 4027 13403 4061
rect 13347 3993 13403 4027
rect 13347 3959 13358 3993
rect 13392 3959 13403 3993
rect 13347 3925 13403 3959
rect 13347 3891 13358 3925
rect 13392 3891 13403 3925
rect 13347 3873 13403 3891
rect 13503 4061 13556 4073
rect 13503 4027 13514 4061
rect 13548 4027 13556 4061
rect 13503 3993 13556 4027
rect 13503 3959 13514 3993
rect 13548 3959 13556 3993
rect 13503 3925 13556 3959
rect 13503 3891 13514 3925
rect 13548 3891 13556 3925
rect 13503 3873 13556 3891
rect 7976 3124 8029 3158
rect 7976 3090 7987 3124
rect 8021 3090 8029 3124
rect 7976 3056 8029 3090
rect 12906 3214 12990 3225
rect 12906 3180 12944 3214
rect 12978 3180 12990 3214
rect 12906 3172 12990 3180
rect 13702 4066 13755 4078
rect 13702 4032 13710 4066
rect 13744 4032 13755 4066
rect 13702 3998 13755 4032
rect 13702 3964 13710 3998
rect 13744 3964 13755 3998
rect 13702 3930 13755 3964
rect 13702 3896 13710 3930
rect 13744 3896 13755 3930
rect 13702 3862 13755 3896
rect 13702 3828 13710 3862
rect 13744 3828 13755 3862
rect 13702 3794 13755 3828
rect 13702 3760 13710 3794
rect 13744 3760 13755 3794
rect 13702 3726 13755 3760
rect 13702 3692 13710 3726
rect 13744 3692 13755 3726
rect 13702 3658 13755 3692
rect 13702 3624 13710 3658
rect 13744 3624 13755 3658
rect 13702 3590 13755 3624
rect 13702 3556 13710 3590
rect 13744 3556 13755 3590
rect 13702 3522 13755 3556
rect 13702 3488 13710 3522
rect 13744 3488 13755 3522
rect 13702 3454 13755 3488
rect 13702 3420 13710 3454
rect 13744 3420 13755 3454
rect 13702 3386 13755 3420
rect 13702 3352 13710 3386
rect 13744 3352 13755 3386
rect 13702 3318 13755 3352
rect 13702 3284 13710 3318
rect 13744 3284 13755 3318
rect 13702 3250 13755 3284
rect 13702 3216 13710 3250
rect 13744 3216 13755 3250
rect 13702 3182 13755 3216
rect 13702 3148 13710 3182
rect 13744 3148 13755 3182
rect 13702 3078 13755 3148
rect 13855 4066 13911 4078
rect 13855 4032 13866 4066
rect 13900 4032 13911 4066
rect 13855 3998 13911 4032
rect 13855 3964 13866 3998
rect 13900 3964 13911 3998
rect 13855 3930 13911 3964
rect 13855 3896 13866 3930
rect 13900 3896 13911 3930
rect 13855 3862 13911 3896
rect 13855 3828 13866 3862
rect 13900 3828 13911 3862
rect 13855 3794 13911 3828
rect 13855 3760 13866 3794
rect 13900 3760 13911 3794
rect 13855 3726 13911 3760
rect 13855 3692 13866 3726
rect 13900 3692 13911 3726
rect 13855 3658 13911 3692
rect 13855 3624 13866 3658
rect 13900 3624 13911 3658
rect 13855 3590 13911 3624
rect 13855 3556 13866 3590
rect 13900 3556 13911 3590
rect 13855 3522 13911 3556
rect 13855 3488 13866 3522
rect 13900 3488 13911 3522
rect 13855 3454 13911 3488
rect 13855 3420 13866 3454
rect 13900 3420 13911 3454
rect 13855 3386 13911 3420
rect 13855 3352 13866 3386
rect 13900 3352 13911 3386
rect 13855 3318 13911 3352
rect 13855 3284 13866 3318
rect 13900 3284 13911 3318
rect 13855 3250 13911 3284
rect 13855 3216 13866 3250
rect 13900 3216 13911 3250
rect 13855 3182 13911 3216
rect 13855 3148 13866 3182
rect 13900 3148 13911 3182
rect 13855 3078 13911 3148
rect 14011 4066 14067 4078
rect 14011 4032 14022 4066
rect 14056 4032 14067 4066
rect 14011 3998 14067 4032
rect 14011 3964 14022 3998
rect 14056 3964 14067 3998
rect 14011 3930 14067 3964
rect 14011 3896 14022 3930
rect 14056 3896 14067 3930
rect 14011 3862 14067 3896
rect 14011 3828 14022 3862
rect 14056 3828 14067 3862
rect 14011 3794 14067 3828
rect 14011 3760 14022 3794
rect 14056 3760 14067 3794
rect 14011 3726 14067 3760
rect 14011 3692 14022 3726
rect 14056 3692 14067 3726
rect 14011 3658 14067 3692
rect 14011 3624 14022 3658
rect 14056 3624 14067 3658
rect 14011 3590 14067 3624
rect 14011 3556 14022 3590
rect 14056 3556 14067 3590
rect 14011 3522 14067 3556
rect 14011 3488 14022 3522
rect 14056 3488 14067 3522
rect 14011 3454 14067 3488
rect 14011 3420 14022 3454
rect 14056 3420 14067 3454
rect 14011 3386 14067 3420
rect 14011 3352 14022 3386
rect 14056 3352 14067 3386
rect 14011 3318 14067 3352
rect 14011 3284 14022 3318
rect 14056 3284 14067 3318
rect 14011 3250 14067 3284
rect 14011 3216 14022 3250
rect 14056 3216 14067 3250
rect 14011 3182 14067 3216
rect 14011 3148 14022 3182
rect 14056 3148 14067 3182
rect 14011 3078 14067 3148
rect 14167 4066 14223 4078
rect 14167 4032 14178 4066
rect 14212 4032 14223 4066
rect 14167 3998 14223 4032
rect 14167 3964 14178 3998
rect 14212 3964 14223 3998
rect 14167 3930 14223 3964
rect 14167 3896 14178 3930
rect 14212 3896 14223 3930
rect 14167 3862 14223 3896
rect 14167 3828 14178 3862
rect 14212 3828 14223 3862
rect 14167 3794 14223 3828
rect 14167 3760 14178 3794
rect 14212 3760 14223 3794
rect 14167 3726 14223 3760
rect 14167 3692 14178 3726
rect 14212 3692 14223 3726
rect 14167 3658 14223 3692
rect 14167 3624 14178 3658
rect 14212 3624 14223 3658
rect 14167 3590 14223 3624
rect 14167 3556 14178 3590
rect 14212 3556 14223 3590
rect 14167 3522 14223 3556
rect 14167 3488 14178 3522
rect 14212 3488 14223 3522
rect 14167 3454 14223 3488
rect 14167 3420 14178 3454
rect 14212 3420 14223 3454
rect 14167 3386 14223 3420
rect 14167 3352 14178 3386
rect 14212 3352 14223 3386
rect 14167 3318 14223 3352
rect 14167 3284 14178 3318
rect 14212 3284 14223 3318
rect 14167 3250 14223 3284
rect 14167 3216 14178 3250
rect 14212 3216 14223 3250
rect 14167 3182 14223 3216
rect 14167 3148 14178 3182
rect 14212 3148 14223 3182
rect 14167 3078 14223 3148
rect 14323 4066 14379 4078
rect 14323 4032 14334 4066
rect 14368 4032 14379 4066
rect 14323 3998 14379 4032
rect 14323 3964 14334 3998
rect 14368 3964 14379 3998
rect 14323 3930 14379 3964
rect 14323 3896 14334 3930
rect 14368 3896 14379 3930
rect 14323 3862 14379 3896
rect 14323 3828 14334 3862
rect 14368 3828 14379 3862
rect 14323 3794 14379 3828
rect 14323 3760 14334 3794
rect 14368 3760 14379 3794
rect 14323 3726 14379 3760
rect 14323 3692 14334 3726
rect 14368 3692 14379 3726
rect 14323 3658 14379 3692
rect 14323 3624 14334 3658
rect 14368 3624 14379 3658
rect 14323 3590 14379 3624
rect 14323 3556 14334 3590
rect 14368 3556 14379 3590
rect 14323 3522 14379 3556
rect 14323 3488 14334 3522
rect 14368 3488 14379 3522
rect 14323 3454 14379 3488
rect 14323 3420 14334 3454
rect 14368 3420 14379 3454
rect 14323 3386 14379 3420
rect 14323 3352 14334 3386
rect 14368 3352 14379 3386
rect 14323 3318 14379 3352
rect 14323 3284 14334 3318
rect 14368 3284 14379 3318
rect 14323 3250 14379 3284
rect 14323 3216 14334 3250
rect 14368 3216 14379 3250
rect 14323 3182 14379 3216
rect 14323 3148 14334 3182
rect 14368 3148 14379 3182
rect 14323 3078 14379 3148
rect 14479 4066 14535 4078
rect 14479 4032 14490 4066
rect 14524 4032 14535 4066
rect 14479 3998 14535 4032
rect 14479 3964 14490 3998
rect 14524 3964 14535 3998
rect 14479 3930 14535 3964
rect 14479 3896 14490 3930
rect 14524 3896 14535 3930
rect 14479 3862 14535 3896
rect 14479 3828 14490 3862
rect 14524 3828 14535 3862
rect 14479 3794 14535 3828
rect 14479 3760 14490 3794
rect 14524 3760 14535 3794
rect 14479 3726 14535 3760
rect 14479 3692 14490 3726
rect 14524 3692 14535 3726
rect 14479 3658 14535 3692
rect 14479 3624 14490 3658
rect 14524 3624 14535 3658
rect 14479 3590 14535 3624
rect 14479 3556 14490 3590
rect 14524 3556 14535 3590
rect 14479 3522 14535 3556
rect 14479 3488 14490 3522
rect 14524 3488 14535 3522
rect 14479 3454 14535 3488
rect 14479 3420 14490 3454
rect 14524 3420 14535 3454
rect 14479 3386 14535 3420
rect 14479 3352 14490 3386
rect 14524 3352 14535 3386
rect 14479 3318 14535 3352
rect 14479 3284 14490 3318
rect 14524 3284 14535 3318
rect 14479 3250 14535 3284
rect 14479 3216 14490 3250
rect 14524 3216 14535 3250
rect 14479 3182 14535 3216
rect 14479 3148 14490 3182
rect 14524 3148 14535 3182
rect 14479 3078 14535 3148
rect 14635 4066 14691 4078
rect 14635 4032 14646 4066
rect 14680 4032 14691 4066
rect 14635 3998 14691 4032
rect 14635 3964 14646 3998
rect 14680 3964 14691 3998
rect 14635 3930 14691 3964
rect 14635 3896 14646 3930
rect 14680 3896 14691 3930
rect 14635 3862 14691 3896
rect 14635 3828 14646 3862
rect 14680 3828 14691 3862
rect 14635 3794 14691 3828
rect 14635 3760 14646 3794
rect 14680 3760 14691 3794
rect 14635 3726 14691 3760
rect 14635 3692 14646 3726
rect 14680 3692 14691 3726
rect 14635 3658 14691 3692
rect 14635 3624 14646 3658
rect 14680 3624 14691 3658
rect 14635 3590 14691 3624
rect 14635 3556 14646 3590
rect 14680 3556 14691 3590
rect 14635 3522 14691 3556
rect 14635 3488 14646 3522
rect 14680 3488 14691 3522
rect 14635 3454 14691 3488
rect 14635 3420 14646 3454
rect 14680 3420 14691 3454
rect 14635 3386 14691 3420
rect 14635 3352 14646 3386
rect 14680 3352 14691 3386
rect 14635 3318 14691 3352
rect 14635 3284 14646 3318
rect 14680 3284 14691 3318
rect 14635 3250 14691 3284
rect 14635 3216 14646 3250
rect 14680 3216 14691 3250
rect 14635 3182 14691 3216
rect 14635 3148 14646 3182
rect 14680 3148 14691 3182
rect 14635 3078 14691 3148
rect 14791 4066 14847 4078
rect 14791 4032 14802 4066
rect 14836 4032 14847 4066
rect 14791 3998 14847 4032
rect 14791 3964 14802 3998
rect 14836 3964 14847 3998
rect 14791 3930 14847 3964
rect 14791 3896 14802 3930
rect 14836 3896 14847 3930
rect 14791 3862 14847 3896
rect 14791 3828 14802 3862
rect 14836 3828 14847 3862
rect 14791 3794 14847 3828
rect 14791 3760 14802 3794
rect 14836 3760 14847 3794
rect 14791 3726 14847 3760
rect 14791 3692 14802 3726
rect 14836 3692 14847 3726
rect 14791 3658 14847 3692
rect 14791 3624 14802 3658
rect 14836 3624 14847 3658
rect 14791 3590 14847 3624
rect 14791 3556 14802 3590
rect 14836 3556 14847 3590
rect 14791 3522 14847 3556
rect 14791 3488 14802 3522
rect 14836 3488 14847 3522
rect 14791 3454 14847 3488
rect 14791 3420 14802 3454
rect 14836 3420 14847 3454
rect 14791 3386 14847 3420
rect 14791 3352 14802 3386
rect 14836 3352 14847 3386
rect 14791 3318 14847 3352
rect 14791 3284 14802 3318
rect 14836 3284 14847 3318
rect 14791 3250 14847 3284
rect 14791 3216 14802 3250
rect 14836 3216 14847 3250
rect 14791 3182 14847 3216
rect 14791 3148 14802 3182
rect 14836 3148 14847 3182
rect 14791 3078 14847 3148
rect 14947 4066 15003 4078
rect 14947 4032 14958 4066
rect 14992 4032 15003 4066
rect 14947 3998 15003 4032
rect 14947 3964 14958 3998
rect 14992 3964 15003 3998
rect 14947 3930 15003 3964
rect 14947 3896 14958 3930
rect 14992 3896 15003 3930
rect 14947 3862 15003 3896
rect 14947 3828 14958 3862
rect 14992 3828 15003 3862
rect 14947 3794 15003 3828
rect 14947 3760 14958 3794
rect 14992 3760 15003 3794
rect 14947 3726 15003 3760
rect 14947 3692 14958 3726
rect 14992 3692 15003 3726
rect 14947 3658 15003 3692
rect 14947 3624 14958 3658
rect 14992 3624 15003 3658
rect 14947 3590 15003 3624
rect 14947 3556 14958 3590
rect 14992 3556 15003 3590
rect 14947 3522 15003 3556
rect 14947 3488 14958 3522
rect 14992 3488 15003 3522
rect 14947 3454 15003 3488
rect 14947 3420 14958 3454
rect 14992 3420 15003 3454
rect 14947 3386 15003 3420
rect 14947 3352 14958 3386
rect 14992 3352 15003 3386
rect 14947 3318 15003 3352
rect 14947 3284 14958 3318
rect 14992 3284 15003 3318
rect 14947 3250 15003 3284
rect 14947 3216 14958 3250
rect 14992 3216 15003 3250
rect 14947 3182 15003 3216
rect 14947 3148 14958 3182
rect 14992 3148 15003 3182
rect 14947 3078 15003 3148
rect 15103 4066 15156 4078
rect 15103 4032 15114 4066
rect 15148 4032 15156 4066
rect 15103 3998 15156 4032
rect 15103 3964 15114 3998
rect 15148 3964 15156 3998
rect 15103 3930 15156 3964
rect 15103 3896 15114 3930
rect 15148 3896 15156 3930
rect 15103 3862 15156 3896
rect 15103 3828 15114 3862
rect 15148 3828 15156 3862
rect 15103 3794 15156 3828
rect 15103 3760 15114 3794
rect 15148 3760 15156 3794
rect 15103 3726 15156 3760
rect 15103 3692 15114 3726
rect 15148 3692 15156 3726
rect 15103 3658 15156 3692
rect 15103 3624 15114 3658
rect 15148 3624 15156 3658
rect 15103 3590 15156 3624
rect 15103 3556 15114 3590
rect 15148 3556 15156 3590
rect 15103 3522 15156 3556
rect 15103 3488 15114 3522
rect 15148 3488 15156 3522
rect 15103 3454 15156 3488
rect 15103 3420 15114 3454
rect 15148 3420 15156 3454
rect 15103 3386 15156 3420
rect 15103 3352 15114 3386
rect 15148 3352 15156 3386
rect 15103 3318 15156 3352
rect 15103 3284 15114 3318
rect 15148 3284 15156 3318
rect 15103 3250 15156 3284
rect 15103 3216 15114 3250
rect 15148 3216 15156 3250
rect 15103 3182 15156 3216
rect 15103 3148 15114 3182
rect 15148 3148 15156 3182
rect 15103 3078 15156 3148
rect 15302 4016 15355 4028
rect 15302 3982 15310 4016
rect 15344 3982 15355 4016
rect 15302 3948 15355 3982
rect 15302 3914 15310 3948
rect 15344 3914 15355 3948
rect 15302 3880 15355 3914
rect 15302 3846 15310 3880
rect 15344 3846 15355 3880
rect 15302 3812 15355 3846
rect 15302 3778 15310 3812
rect 15344 3778 15355 3812
rect 15302 3744 15355 3778
rect 15302 3710 15310 3744
rect 15344 3710 15355 3744
rect 15302 3676 15355 3710
rect 15302 3642 15310 3676
rect 15344 3642 15355 3676
rect 15302 3608 15355 3642
rect 15302 3574 15310 3608
rect 15344 3574 15355 3608
rect 15302 3540 15355 3574
rect 15302 3506 15310 3540
rect 15344 3506 15355 3540
rect 15302 3472 15355 3506
rect 15302 3438 15310 3472
rect 15344 3438 15355 3472
rect 15302 3404 15355 3438
rect 15302 3370 15310 3404
rect 15344 3370 15355 3404
rect 15302 3336 15355 3370
rect 15302 3302 15310 3336
rect 15344 3302 15355 3336
rect 15302 3268 15355 3302
rect 15302 3234 15310 3268
rect 15344 3234 15355 3268
rect 15302 3200 15355 3234
rect 15302 3166 15310 3200
rect 15344 3166 15355 3200
rect 15302 3132 15355 3166
rect 15302 3098 15310 3132
rect 15344 3098 15355 3132
rect 7976 3022 7987 3056
rect 8021 3022 8029 3056
rect 7976 3010 8029 3022
rect 15302 3028 15355 3098
rect 15455 4016 15511 4028
rect 15455 3982 15466 4016
rect 15500 3982 15511 4016
rect 15455 3948 15511 3982
rect 15455 3914 15466 3948
rect 15500 3914 15511 3948
rect 15455 3880 15511 3914
rect 15455 3846 15466 3880
rect 15500 3846 15511 3880
rect 15455 3812 15511 3846
rect 15455 3778 15466 3812
rect 15500 3778 15511 3812
rect 15455 3744 15511 3778
rect 15455 3710 15466 3744
rect 15500 3710 15511 3744
rect 15455 3676 15511 3710
rect 15455 3642 15466 3676
rect 15500 3642 15511 3676
rect 15455 3608 15511 3642
rect 15455 3574 15466 3608
rect 15500 3574 15511 3608
rect 15455 3540 15511 3574
rect 15455 3506 15466 3540
rect 15500 3506 15511 3540
rect 15455 3472 15511 3506
rect 15455 3438 15466 3472
rect 15500 3438 15511 3472
rect 15455 3404 15511 3438
rect 15455 3370 15466 3404
rect 15500 3370 15511 3404
rect 15455 3336 15511 3370
rect 15455 3302 15466 3336
rect 15500 3302 15511 3336
rect 15455 3268 15511 3302
rect 15455 3234 15466 3268
rect 15500 3234 15511 3268
rect 15455 3200 15511 3234
rect 15455 3166 15466 3200
rect 15500 3166 15511 3200
rect 15455 3132 15511 3166
rect 15455 3098 15466 3132
rect 15500 3098 15511 3132
rect 15455 3028 15511 3098
rect 15611 4016 15667 4028
rect 15611 3982 15622 4016
rect 15656 3982 15667 4016
rect 15611 3948 15667 3982
rect 15611 3914 15622 3948
rect 15656 3914 15667 3948
rect 15611 3880 15667 3914
rect 15611 3846 15622 3880
rect 15656 3846 15667 3880
rect 15611 3812 15667 3846
rect 15611 3778 15622 3812
rect 15656 3778 15667 3812
rect 15611 3744 15667 3778
rect 15611 3710 15622 3744
rect 15656 3710 15667 3744
rect 15611 3676 15667 3710
rect 15611 3642 15622 3676
rect 15656 3642 15667 3676
rect 15611 3608 15667 3642
rect 15611 3574 15622 3608
rect 15656 3574 15667 3608
rect 15611 3540 15667 3574
rect 15611 3506 15622 3540
rect 15656 3506 15667 3540
rect 15611 3472 15667 3506
rect 15611 3438 15622 3472
rect 15656 3438 15667 3472
rect 15611 3404 15667 3438
rect 15611 3370 15622 3404
rect 15656 3370 15667 3404
rect 15611 3336 15667 3370
rect 15611 3302 15622 3336
rect 15656 3302 15667 3336
rect 15611 3268 15667 3302
rect 15611 3234 15622 3268
rect 15656 3234 15667 3268
rect 15611 3200 15667 3234
rect 15611 3166 15622 3200
rect 15656 3166 15667 3200
rect 15611 3132 15667 3166
rect 15611 3098 15622 3132
rect 15656 3098 15667 3132
rect 15611 3028 15667 3098
rect 15767 4016 15823 4028
rect 15767 3982 15778 4016
rect 15812 3982 15823 4016
rect 15767 3948 15823 3982
rect 15767 3914 15778 3948
rect 15812 3914 15823 3948
rect 15767 3880 15823 3914
rect 15767 3846 15778 3880
rect 15812 3846 15823 3880
rect 15767 3812 15823 3846
rect 15767 3778 15778 3812
rect 15812 3778 15823 3812
rect 15767 3744 15823 3778
rect 15767 3710 15778 3744
rect 15812 3710 15823 3744
rect 15767 3676 15823 3710
rect 15767 3642 15778 3676
rect 15812 3642 15823 3676
rect 15767 3608 15823 3642
rect 15767 3574 15778 3608
rect 15812 3574 15823 3608
rect 15767 3540 15823 3574
rect 15767 3506 15778 3540
rect 15812 3506 15823 3540
rect 15767 3472 15823 3506
rect 15767 3438 15778 3472
rect 15812 3438 15823 3472
rect 15767 3404 15823 3438
rect 15767 3370 15778 3404
rect 15812 3370 15823 3404
rect 15767 3336 15823 3370
rect 15767 3302 15778 3336
rect 15812 3302 15823 3336
rect 15767 3268 15823 3302
rect 15767 3234 15778 3268
rect 15812 3234 15823 3268
rect 15767 3200 15823 3234
rect 15767 3166 15778 3200
rect 15812 3166 15823 3200
rect 15767 3132 15823 3166
rect 15767 3098 15778 3132
rect 15812 3098 15823 3132
rect 15767 3028 15823 3098
rect 15923 4016 15979 4028
rect 15923 3982 15934 4016
rect 15968 3982 15979 4016
rect 15923 3948 15979 3982
rect 15923 3914 15934 3948
rect 15968 3914 15979 3948
rect 15923 3880 15979 3914
rect 15923 3846 15934 3880
rect 15968 3846 15979 3880
rect 15923 3812 15979 3846
rect 15923 3778 15934 3812
rect 15968 3778 15979 3812
rect 15923 3744 15979 3778
rect 15923 3710 15934 3744
rect 15968 3710 15979 3744
rect 15923 3676 15979 3710
rect 15923 3642 15934 3676
rect 15968 3642 15979 3676
rect 15923 3608 15979 3642
rect 15923 3574 15934 3608
rect 15968 3574 15979 3608
rect 15923 3540 15979 3574
rect 15923 3506 15934 3540
rect 15968 3506 15979 3540
rect 15923 3472 15979 3506
rect 15923 3438 15934 3472
rect 15968 3438 15979 3472
rect 15923 3404 15979 3438
rect 15923 3370 15934 3404
rect 15968 3370 15979 3404
rect 15923 3336 15979 3370
rect 15923 3302 15934 3336
rect 15968 3302 15979 3336
rect 15923 3268 15979 3302
rect 15923 3234 15934 3268
rect 15968 3234 15979 3268
rect 15923 3200 15979 3234
rect 15923 3166 15934 3200
rect 15968 3166 15979 3200
rect 15923 3132 15979 3166
rect 15923 3098 15934 3132
rect 15968 3098 15979 3132
rect 15923 3028 15979 3098
rect 16079 4016 16135 4028
rect 16079 3982 16090 4016
rect 16124 3982 16135 4016
rect 16079 3948 16135 3982
rect 16079 3914 16090 3948
rect 16124 3914 16135 3948
rect 16079 3880 16135 3914
rect 16079 3846 16090 3880
rect 16124 3846 16135 3880
rect 16079 3812 16135 3846
rect 16079 3778 16090 3812
rect 16124 3778 16135 3812
rect 16079 3744 16135 3778
rect 16079 3710 16090 3744
rect 16124 3710 16135 3744
rect 16079 3676 16135 3710
rect 16079 3642 16090 3676
rect 16124 3642 16135 3676
rect 16079 3608 16135 3642
rect 16079 3574 16090 3608
rect 16124 3574 16135 3608
rect 16079 3540 16135 3574
rect 16079 3506 16090 3540
rect 16124 3506 16135 3540
rect 16079 3472 16135 3506
rect 16079 3438 16090 3472
rect 16124 3438 16135 3472
rect 16079 3404 16135 3438
rect 16079 3370 16090 3404
rect 16124 3370 16135 3404
rect 16079 3336 16135 3370
rect 16079 3302 16090 3336
rect 16124 3302 16135 3336
rect 16079 3268 16135 3302
rect 16079 3234 16090 3268
rect 16124 3234 16135 3268
rect 16079 3200 16135 3234
rect 16079 3166 16090 3200
rect 16124 3166 16135 3200
rect 16079 3132 16135 3166
rect 16079 3098 16090 3132
rect 16124 3098 16135 3132
rect 16079 3028 16135 3098
rect 16235 4016 16291 4028
rect 16235 3982 16246 4016
rect 16280 3982 16291 4016
rect 16235 3948 16291 3982
rect 16235 3914 16246 3948
rect 16280 3914 16291 3948
rect 16235 3880 16291 3914
rect 16235 3846 16246 3880
rect 16280 3846 16291 3880
rect 16235 3812 16291 3846
rect 16235 3778 16246 3812
rect 16280 3778 16291 3812
rect 16235 3744 16291 3778
rect 16235 3710 16246 3744
rect 16280 3710 16291 3744
rect 16235 3676 16291 3710
rect 16235 3642 16246 3676
rect 16280 3642 16291 3676
rect 16235 3608 16291 3642
rect 16235 3574 16246 3608
rect 16280 3574 16291 3608
rect 16235 3540 16291 3574
rect 16235 3506 16246 3540
rect 16280 3506 16291 3540
rect 16235 3472 16291 3506
rect 16235 3438 16246 3472
rect 16280 3438 16291 3472
rect 16235 3404 16291 3438
rect 16235 3370 16246 3404
rect 16280 3370 16291 3404
rect 16235 3336 16291 3370
rect 16235 3302 16246 3336
rect 16280 3302 16291 3336
rect 16235 3268 16291 3302
rect 16235 3234 16246 3268
rect 16280 3234 16291 3268
rect 16235 3200 16291 3234
rect 16235 3166 16246 3200
rect 16280 3166 16291 3200
rect 16235 3132 16291 3166
rect 16235 3098 16246 3132
rect 16280 3098 16291 3132
rect 16235 3028 16291 3098
rect 16391 4016 16447 4028
rect 16391 3982 16402 4016
rect 16436 3982 16447 4016
rect 16391 3948 16447 3982
rect 16391 3914 16402 3948
rect 16436 3914 16447 3948
rect 16391 3880 16447 3914
rect 16391 3846 16402 3880
rect 16436 3846 16447 3880
rect 16391 3812 16447 3846
rect 16391 3778 16402 3812
rect 16436 3778 16447 3812
rect 16391 3744 16447 3778
rect 16391 3710 16402 3744
rect 16436 3710 16447 3744
rect 16391 3676 16447 3710
rect 16391 3642 16402 3676
rect 16436 3642 16447 3676
rect 16391 3608 16447 3642
rect 16391 3574 16402 3608
rect 16436 3574 16447 3608
rect 16391 3540 16447 3574
rect 16391 3506 16402 3540
rect 16436 3506 16447 3540
rect 16391 3472 16447 3506
rect 16391 3438 16402 3472
rect 16436 3438 16447 3472
rect 16391 3404 16447 3438
rect 16391 3370 16402 3404
rect 16436 3370 16447 3404
rect 16391 3336 16447 3370
rect 16391 3302 16402 3336
rect 16436 3302 16447 3336
rect 16391 3268 16447 3302
rect 16391 3234 16402 3268
rect 16436 3234 16447 3268
rect 16391 3200 16447 3234
rect 16391 3166 16402 3200
rect 16436 3166 16447 3200
rect 16391 3132 16447 3166
rect 16391 3098 16402 3132
rect 16436 3098 16447 3132
rect 16391 3028 16447 3098
rect 16547 4016 16600 4028
rect 16547 3982 16558 4016
rect 16592 3982 16600 4016
rect 16547 3948 16600 3982
rect 16547 3914 16558 3948
rect 16592 3914 16600 3948
rect 16547 3880 16600 3914
rect 16547 3846 16558 3880
rect 16592 3846 16600 3880
rect 16547 3812 16600 3846
rect 16547 3778 16558 3812
rect 16592 3778 16600 3812
rect 16547 3744 16600 3778
rect 16547 3710 16558 3744
rect 16592 3710 16600 3744
rect 16547 3676 16600 3710
rect 16547 3642 16558 3676
rect 16592 3642 16600 3676
rect 16547 3608 16600 3642
rect 16547 3574 16558 3608
rect 16592 3574 16600 3608
rect 16547 3540 16600 3574
rect 16547 3506 16558 3540
rect 16592 3506 16600 3540
rect 16547 3472 16600 3506
rect 16547 3438 16558 3472
rect 16592 3438 16600 3472
rect 16547 3404 16600 3438
rect 16547 3370 16558 3404
rect 16592 3370 16600 3404
rect 16547 3336 16600 3370
rect 16547 3302 16558 3336
rect 16592 3302 16600 3336
rect 16547 3268 16600 3302
rect 16547 3234 16558 3268
rect 16592 3234 16600 3268
rect 16547 3200 16600 3234
rect 16547 3166 16558 3200
rect 16592 3166 16600 3200
rect 16547 3132 16600 3166
rect 16547 3098 16558 3132
rect 16592 3098 16600 3132
rect 16547 3028 16600 3098
rect 16746 4066 16799 4078
rect 16746 4032 16754 4066
rect 16788 4032 16799 4066
rect 16746 3998 16799 4032
rect 16746 3964 16754 3998
rect 16788 3964 16799 3998
rect 16746 3930 16799 3964
rect 16746 3896 16754 3930
rect 16788 3896 16799 3930
rect 16746 3862 16799 3896
rect 16746 3828 16754 3862
rect 16788 3828 16799 3862
rect 16746 3794 16799 3828
rect 16746 3760 16754 3794
rect 16788 3760 16799 3794
rect 16746 3726 16799 3760
rect 16746 3692 16754 3726
rect 16788 3692 16799 3726
rect 16746 3658 16799 3692
rect 16746 3624 16754 3658
rect 16788 3624 16799 3658
rect 16746 3590 16799 3624
rect 16746 3556 16754 3590
rect 16788 3556 16799 3590
rect 16746 3522 16799 3556
rect 16746 3488 16754 3522
rect 16788 3488 16799 3522
rect 16746 3454 16799 3488
rect 16746 3420 16754 3454
rect 16788 3420 16799 3454
rect 16746 3386 16799 3420
rect 16746 3352 16754 3386
rect 16788 3352 16799 3386
rect 16746 3318 16799 3352
rect 16746 3284 16754 3318
rect 16788 3284 16799 3318
rect 16746 3250 16799 3284
rect 16746 3216 16754 3250
rect 16788 3216 16799 3250
rect 16746 3182 16799 3216
rect 16746 3148 16754 3182
rect 16788 3148 16799 3182
rect 16746 3078 16799 3148
rect 16899 4066 16955 4078
rect 16899 4032 16910 4066
rect 16944 4032 16955 4066
rect 16899 3998 16955 4032
rect 16899 3964 16910 3998
rect 16944 3964 16955 3998
rect 16899 3930 16955 3964
rect 16899 3896 16910 3930
rect 16944 3896 16955 3930
rect 16899 3862 16955 3896
rect 16899 3828 16910 3862
rect 16944 3828 16955 3862
rect 16899 3794 16955 3828
rect 16899 3760 16910 3794
rect 16944 3760 16955 3794
rect 16899 3726 16955 3760
rect 16899 3692 16910 3726
rect 16944 3692 16955 3726
rect 16899 3658 16955 3692
rect 16899 3624 16910 3658
rect 16944 3624 16955 3658
rect 16899 3590 16955 3624
rect 16899 3556 16910 3590
rect 16944 3556 16955 3590
rect 16899 3522 16955 3556
rect 16899 3488 16910 3522
rect 16944 3488 16955 3522
rect 16899 3454 16955 3488
rect 16899 3420 16910 3454
rect 16944 3420 16955 3454
rect 16899 3386 16955 3420
rect 16899 3352 16910 3386
rect 16944 3352 16955 3386
rect 16899 3318 16955 3352
rect 16899 3284 16910 3318
rect 16944 3284 16955 3318
rect 16899 3250 16955 3284
rect 16899 3216 16910 3250
rect 16944 3216 16955 3250
rect 16899 3182 16955 3216
rect 16899 3148 16910 3182
rect 16944 3148 16955 3182
rect 16899 3078 16955 3148
rect 17055 4066 17111 4078
rect 17055 4032 17066 4066
rect 17100 4032 17111 4066
rect 17055 3998 17111 4032
rect 17055 3964 17066 3998
rect 17100 3964 17111 3998
rect 17055 3930 17111 3964
rect 17055 3896 17066 3930
rect 17100 3896 17111 3930
rect 17055 3862 17111 3896
rect 17055 3828 17066 3862
rect 17100 3828 17111 3862
rect 17055 3794 17111 3828
rect 17055 3760 17066 3794
rect 17100 3760 17111 3794
rect 17055 3726 17111 3760
rect 17055 3692 17066 3726
rect 17100 3692 17111 3726
rect 17055 3658 17111 3692
rect 17055 3624 17066 3658
rect 17100 3624 17111 3658
rect 17055 3590 17111 3624
rect 17055 3556 17066 3590
rect 17100 3556 17111 3590
rect 17055 3522 17111 3556
rect 17055 3488 17066 3522
rect 17100 3488 17111 3522
rect 17055 3454 17111 3488
rect 17055 3420 17066 3454
rect 17100 3420 17111 3454
rect 17055 3386 17111 3420
rect 17055 3352 17066 3386
rect 17100 3352 17111 3386
rect 17055 3318 17111 3352
rect 17055 3284 17066 3318
rect 17100 3284 17111 3318
rect 17055 3250 17111 3284
rect 17055 3216 17066 3250
rect 17100 3216 17111 3250
rect 17055 3182 17111 3216
rect 17055 3148 17066 3182
rect 17100 3148 17111 3182
rect 17055 3078 17111 3148
rect 17211 4066 17267 4078
rect 17211 4032 17222 4066
rect 17256 4032 17267 4066
rect 17211 3998 17267 4032
rect 17211 3964 17222 3998
rect 17256 3964 17267 3998
rect 17211 3930 17267 3964
rect 17211 3896 17222 3930
rect 17256 3896 17267 3930
rect 17211 3862 17267 3896
rect 17211 3828 17222 3862
rect 17256 3828 17267 3862
rect 17211 3794 17267 3828
rect 17211 3760 17222 3794
rect 17256 3760 17267 3794
rect 17211 3726 17267 3760
rect 17211 3692 17222 3726
rect 17256 3692 17267 3726
rect 17211 3658 17267 3692
rect 17211 3624 17222 3658
rect 17256 3624 17267 3658
rect 17211 3590 17267 3624
rect 17211 3556 17222 3590
rect 17256 3556 17267 3590
rect 17211 3522 17267 3556
rect 17211 3488 17222 3522
rect 17256 3488 17267 3522
rect 17211 3454 17267 3488
rect 17211 3420 17222 3454
rect 17256 3420 17267 3454
rect 17211 3386 17267 3420
rect 17211 3352 17222 3386
rect 17256 3352 17267 3386
rect 17211 3318 17267 3352
rect 17211 3284 17222 3318
rect 17256 3284 17267 3318
rect 17211 3250 17267 3284
rect 17211 3216 17222 3250
rect 17256 3216 17267 3250
rect 17211 3182 17267 3216
rect 17211 3148 17222 3182
rect 17256 3148 17267 3182
rect 17211 3078 17267 3148
rect 17367 4066 17423 4078
rect 17367 4032 17378 4066
rect 17412 4032 17423 4066
rect 17367 3998 17423 4032
rect 17367 3964 17378 3998
rect 17412 3964 17423 3998
rect 17367 3930 17423 3964
rect 17367 3896 17378 3930
rect 17412 3896 17423 3930
rect 17367 3862 17423 3896
rect 17367 3828 17378 3862
rect 17412 3828 17423 3862
rect 17367 3794 17423 3828
rect 17367 3760 17378 3794
rect 17412 3760 17423 3794
rect 17367 3726 17423 3760
rect 17367 3692 17378 3726
rect 17412 3692 17423 3726
rect 17367 3658 17423 3692
rect 17367 3624 17378 3658
rect 17412 3624 17423 3658
rect 17367 3590 17423 3624
rect 17367 3556 17378 3590
rect 17412 3556 17423 3590
rect 17367 3522 17423 3556
rect 17367 3488 17378 3522
rect 17412 3488 17423 3522
rect 17367 3454 17423 3488
rect 17367 3420 17378 3454
rect 17412 3420 17423 3454
rect 17367 3386 17423 3420
rect 17367 3352 17378 3386
rect 17412 3352 17423 3386
rect 17367 3318 17423 3352
rect 17367 3284 17378 3318
rect 17412 3284 17423 3318
rect 17367 3250 17423 3284
rect 17367 3216 17378 3250
rect 17412 3216 17423 3250
rect 17367 3182 17423 3216
rect 17367 3148 17378 3182
rect 17412 3148 17423 3182
rect 17367 3078 17423 3148
rect 17523 4066 17579 4078
rect 17523 4032 17534 4066
rect 17568 4032 17579 4066
rect 17523 3998 17579 4032
rect 17523 3964 17534 3998
rect 17568 3964 17579 3998
rect 17523 3930 17579 3964
rect 17523 3896 17534 3930
rect 17568 3896 17579 3930
rect 17523 3862 17579 3896
rect 17523 3828 17534 3862
rect 17568 3828 17579 3862
rect 17523 3794 17579 3828
rect 17523 3760 17534 3794
rect 17568 3760 17579 3794
rect 17523 3726 17579 3760
rect 17523 3692 17534 3726
rect 17568 3692 17579 3726
rect 17523 3658 17579 3692
rect 17523 3624 17534 3658
rect 17568 3624 17579 3658
rect 17523 3590 17579 3624
rect 17523 3556 17534 3590
rect 17568 3556 17579 3590
rect 17523 3522 17579 3556
rect 17523 3488 17534 3522
rect 17568 3488 17579 3522
rect 17523 3454 17579 3488
rect 17523 3420 17534 3454
rect 17568 3420 17579 3454
rect 17523 3386 17579 3420
rect 17523 3352 17534 3386
rect 17568 3352 17579 3386
rect 17523 3318 17579 3352
rect 17523 3284 17534 3318
rect 17568 3284 17579 3318
rect 17523 3250 17579 3284
rect 17523 3216 17534 3250
rect 17568 3216 17579 3250
rect 17523 3182 17579 3216
rect 17523 3148 17534 3182
rect 17568 3148 17579 3182
rect 17523 3078 17579 3148
rect 17679 4066 17735 4078
rect 17679 4032 17690 4066
rect 17724 4032 17735 4066
rect 17679 3998 17735 4032
rect 17679 3964 17690 3998
rect 17724 3964 17735 3998
rect 17679 3930 17735 3964
rect 17679 3896 17690 3930
rect 17724 3896 17735 3930
rect 17679 3862 17735 3896
rect 17679 3828 17690 3862
rect 17724 3828 17735 3862
rect 17679 3794 17735 3828
rect 17679 3760 17690 3794
rect 17724 3760 17735 3794
rect 17679 3726 17735 3760
rect 17679 3692 17690 3726
rect 17724 3692 17735 3726
rect 17679 3658 17735 3692
rect 17679 3624 17690 3658
rect 17724 3624 17735 3658
rect 17679 3590 17735 3624
rect 17679 3556 17690 3590
rect 17724 3556 17735 3590
rect 17679 3522 17735 3556
rect 17679 3488 17690 3522
rect 17724 3488 17735 3522
rect 17679 3454 17735 3488
rect 17679 3420 17690 3454
rect 17724 3420 17735 3454
rect 17679 3386 17735 3420
rect 17679 3352 17690 3386
rect 17724 3352 17735 3386
rect 17679 3318 17735 3352
rect 17679 3284 17690 3318
rect 17724 3284 17735 3318
rect 17679 3250 17735 3284
rect 17679 3216 17690 3250
rect 17724 3216 17735 3250
rect 17679 3182 17735 3216
rect 17679 3148 17690 3182
rect 17724 3148 17735 3182
rect 17679 3078 17735 3148
rect 17835 4066 17891 4078
rect 17835 4032 17846 4066
rect 17880 4032 17891 4066
rect 17835 3998 17891 4032
rect 17835 3964 17846 3998
rect 17880 3964 17891 3998
rect 17835 3930 17891 3964
rect 17835 3896 17846 3930
rect 17880 3896 17891 3930
rect 17835 3862 17891 3896
rect 17835 3828 17846 3862
rect 17880 3828 17891 3862
rect 17835 3794 17891 3828
rect 17835 3760 17846 3794
rect 17880 3760 17891 3794
rect 17835 3726 17891 3760
rect 17835 3692 17846 3726
rect 17880 3692 17891 3726
rect 17835 3658 17891 3692
rect 17835 3624 17846 3658
rect 17880 3624 17891 3658
rect 17835 3590 17891 3624
rect 17835 3556 17846 3590
rect 17880 3556 17891 3590
rect 17835 3522 17891 3556
rect 17835 3488 17846 3522
rect 17880 3488 17891 3522
rect 17835 3454 17891 3488
rect 17835 3420 17846 3454
rect 17880 3420 17891 3454
rect 17835 3386 17891 3420
rect 17835 3352 17846 3386
rect 17880 3352 17891 3386
rect 17835 3318 17891 3352
rect 17835 3284 17846 3318
rect 17880 3284 17891 3318
rect 17835 3250 17891 3284
rect 17835 3216 17846 3250
rect 17880 3216 17891 3250
rect 17835 3182 17891 3216
rect 17835 3148 17846 3182
rect 17880 3148 17891 3182
rect 17835 3078 17891 3148
rect 17991 4066 18044 4078
rect 17991 4032 18002 4066
rect 18036 4032 18044 4066
rect 17991 3998 18044 4032
rect 17991 3964 18002 3998
rect 18036 3964 18044 3998
rect 17991 3930 18044 3964
rect 17991 3896 18002 3930
rect 18036 3896 18044 3930
rect 17991 3862 18044 3896
rect 17991 3828 18002 3862
rect 18036 3828 18044 3862
rect 17991 3794 18044 3828
rect 17991 3760 18002 3794
rect 18036 3760 18044 3794
rect 17991 3726 18044 3760
rect 17991 3692 18002 3726
rect 18036 3692 18044 3726
rect 17991 3658 18044 3692
rect 17991 3624 18002 3658
rect 18036 3624 18044 3658
rect 17991 3590 18044 3624
rect 17991 3556 18002 3590
rect 18036 3556 18044 3590
rect 17991 3522 18044 3556
rect 17991 3488 18002 3522
rect 18036 3488 18044 3522
rect 17991 3454 18044 3488
rect 17991 3420 18002 3454
rect 18036 3420 18044 3454
rect 17991 3386 18044 3420
rect 17991 3352 18002 3386
rect 18036 3352 18044 3386
rect 17991 3318 18044 3352
rect 17991 3284 18002 3318
rect 18036 3284 18044 3318
rect 17991 3250 18044 3284
rect 17991 3216 18002 3250
rect 18036 3216 18044 3250
rect 17991 3182 18044 3216
rect 17991 3148 18002 3182
rect 18036 3148 18044 3182
rect 17991 3078 18044 3148
rect 18190 4066 18243 4078
rect 18190 4032 18198 4066
rect 18232 4032 18243 4066
rect 18190 3998 18243 4032
rect 18190 3964 18198 3998
rect 18232 3964 18243 3998
rect 18190 3930 18243 3964
rect 18190 3896 18198 3930
rect 18232 3896 18243 3930
rect 18190 3862 18243 3896
rect 18190 3828 18198 3862
rect 18232 3828 18243 3862
rect 18190 3794 18243 3828
rect 18190 3760 18198 3794
rect 18232 3760 18243 3794
rect 18190 3726 18243 3760
rect 18190 3692 18198 3726
rect 18232 3692 18243 3726
rect 18190 3658 18243 3692
rect 18190 3624 18198 3658
rect 18232 3624 18243 3658
rect 18190 3590 18243 3624
rect 18190 3556 18198 3590
rect 18232 3556 18243 3590
rect 18190 3522 18243 3556
rect 18190 3488 18198 3522
rect 18232 3488 18243 3522
rect 18190 3454 18243 3488
rect 18190 3420 18198 3454
rect 18232 3420 18243 3454
rect 18190 3386 18243 3420
rect 18190 3352 18198 3386
rect 18232 3352 18243 3386
rect 18190 3318 18243 3352
rect 18190 3284 18198 3318
rect 18232 3284 18243 3318
rect 18190 3250 18243 3284
rect 18190 3216 18198 3250
rect 18232 3216 18243 3250
rect 18190 3182 18243 3216
rect 18190 3148 18198 3182
rect 18232 3148 18243 3182
rect 18190 3078 18243 3148
rect 18343 4066 18399 4078
rect 18343 4032 18354 4066
rect 18388 4032 18399 4066
rect 18343 3998 18399 4032
rect 18343 3964 18354 3998
rect 18388 3964 18399 3998
rect 18343 3930 18399 3964
rect 18343 3896 18354 3930
rect 18388 3896 18399 3930
rect 18343 3862 18399 3896
rect 18343 3828 18354 3862
rect 18388 3828 18399 3862
rect 18343 3794 18399 3828
rect 18343 3760 18354 3794
rect 18388 3760 18399 3794
rect 18343 3726 18399 3760
rect 18343 3692 18354 3726
rect 18388 3692 18399 3726
rect 18343 3658 18399 3692
rect 18343 3624 18354 3658
rect 18388 3624 18399 3658
rect 18343 3590 18399 3624
rect 18343 3556 18354 3590
rect 18388 3556 18399 3590
rect 18343 3522 18399 3556
rect 18343 3488 18354 3522
rect 18388 3488 18399 3522
rect 18343 3454 18399 3488
rect 18343 3420 18354 3454
rect 18388 3420 18399 3454
rect 18343 3386 18399 3420
rect 18343 3352 18354 3386
rect 18388 3352 18399 3386
rect 18343 3318 18399 3352
rect 18343 3284 18354 3318
rect 18388 3284 18399 3318
rect 18343 3250 18399 3284
rect 18343 3216 18354 3250
rect 18388 3216 18399 3250
rect 18343 3182 18399 3216
rect 18343 3148 18354 3182
rect 18388 3148 18399 3182
rect 18343 3078 18399 3148
rect 18499 4066 18555 4078
rect 18499 4032 18510 4066
rect 18544 4032 18555 4066
rect 18499 3998 18555 4032
rect 18499 3964 18510 3998
rect 18544 3964 18555 3998
rect 18499 3930 18555 3964
rect 18499 3896 18510 3930
rect 18544 3896 18555 3930
rect 18499 3862 18555 3896
rect 18499 3828 18510 3862
rect 18544 3828 18555 3862
rect 18499 3794 18555 3828
rect 18499 3760 18510 3794
rect 18544 3760 18555 3794
rect 18499 3726 18555 3760
rect 18499 3692 18510 3726
rect 18544 3692 18555 3726
rect 18499 3658 18555 3692
rect 18499 3624 18510 3658
rect 18544 3624 18555 3658
rect 18499 3590 18555 3624
rect 18499 3556 18510 3590
rect 18544 3556 18555 3590
rect 18499 3522 18555 3556
rect 18499 3488 18510 3522
rect 18544 3488 18555 3522
rect 18499 3454 18555 3488
rect 18499 3420 18510 3454
rect 18544 3420 18555 3454
rect 18499 3386 18555 3420
rect 18499 3352 18510 3386
rect 18544 3352 18555 3386
rect 18499 3318 18555 3352
rect 18499 3284 18510 3318
rect 18544 3284 18555 3318
rect 18499 3250 18555 3284
rect 18499 3216 18510 3250
rect 18544 3216 18555 3250
rect 18499 3182 18555 3216
rect 18499 3148 18510 3182
rect 18544 3148 18555 3182
rect 18499 3078 18555 3148
rect 18655 4066 18711 4078
rect 18655 4032 18666 4066
rect 18700 4032 18711 4066
rect 18655 3998 18711 4032
rect 18655 3964 18666 3998
rect 18700 3964 18711 3998
rect 18655 3930 18711 3964
rect 18655 3896 18666 3930
rect 18700 3896 18711 3930
rect 18655 3862 18711 3896
rect 18655 3828 18666 3862
rect 18700 3828 18711 3862
rect 18655 3794 18711 3828
rect 18655 3760 18666 3794
rect 18700 3760 18711 3794
rect 18655 3726 18711 3760
rect 18655 3692 18666 3726
rect 18700 3692 18711 3726
rect 18655 3658 18711 3692
rect 18655 3624 18666 3658
rect 18700 3624 18711 3658
rect 18655 3590 18711 3624
rect 18655 3556 18666 3590
rect 18700 3556 18711 3590
rect 18655 3522 18711 3556
rect 18655 3488 18666 3522
rect 18700 3488 18711 3522
rect 18655 3454 18711 3488
rect 18655 3420 18666 3454
rect 18700 3420 18711 3454
rect 18655 3386 18711 3420
rect 18655 3352 18666 3386
rect 18700 3352 18711 3386
rect 18655 3318 18711 3352
rect 18655 3284 18666 3318
rect 18700 3284 18711 3318
rect 18655 3250 18711 3284
rect 18655 3216 18666 3250
rect 18700 3216 18711 3250
rect 18655 3182 18711 3216
rect 18655 3148 18666 3182
rect 18700 3148 18711 3182
rect 18655 3078 18711 3148
rect 18811 4066 18867 4078
rect 18811 4032 18822 4066
rect 18856 4032 18867 4066
rect 18811 3998 18867 4032
rect 18811 3964 18822 3998
rect 18856 3964 18867 3998
rect 18811 3930 18867 3964
rect 18811 3896 18822 3930
rect 18856 3896 18867 3930
rect 18811 3862 18867 3896
rect 18811 3828 18822 3862
rect 18856 3828 18867 3862
rect 18811 3794 18867 3828
rect 18811 3760 18822 3794
rect 18856 3760 18867 3794
rect 18811 3726 18867 3760
rect 18811 3692 18822 3726
rect 18856 3692 18867 3726
rect 18811 3658 18867 3692
rect 18811 3624 18822 3658
rect 18856 3624 18867 3658
rect 18811 3590 18867 3624
rect 18811 3556 18822 3590
rect 18856 3556 18867 3590
rect 18811 3522 18867 3556
rect 18811 3488 18822 3522
rect 18856 3488 18867 3522
rect 18811 3454 18867 3488
rect 18811 3420 18822 3454
rect 18856 3420 18867 3454
rect 18811 3386 18867 3420
rect 18811 3352 18822 3386
rect 18856 3352 18867 3386
rect 18811 3318 18867 3352
rect 18811 3284 18822 3318
rect 18856 3284 18867 3318
rect 18811 3250 18867 3284
rect 18811 3216 18822 3250
rect 18856 3216 18867 3250
rect 18811 3182 18867 3216
rect 18811 3148 18822 3182
rect 18856 3148 18867 3182
rect 18811 3078 18867 3148
rect 18967 4066 19023 4078
rect 18967 4032 18978 4066
rect 19012 4032 19023 4066
rect 18967 3998 19023 4032
rect 18967 3964 18978 3998
rect 19012 3964 19023 3998
rect 18967 3930 19023 3964
rect 18967 3896 18978 3930
rect 19012 3896 19023 3930
rect 18967 3862 19023 3896
rect 18967 3828 18978 3862
rect 19012 3828 19023 3862
rect 18967 3794 19023 3828
rect 18967 3760 18978 3794
rect 19012 3760 19023 3794
rect 18967 3726 19023 3760
rect 18967 3692 18978 3726
rect 19012 3692 19023 3726
rect 18967 3658 19023 3692
rect 18967 3624 18978 3658
rect 19012 3624 19023 3658
rect 18967 3590 19023 3624
rect 18967 3556 18978 3590
rect 19012 3556 19023 3590
rect 18967 3522 19023 3556
rect 18967 3488 18978 3522
rect 19012 3488 19023 3522
rect 18967 3454 19023 3488
rect 18967 3420 18978 3454
rect 19012 3420 19023 3454
rect 18967 3386 19023 3420
rect 18967 3352 18978 3386
rect 19012 3352 19023 3386
rect 18967 3318 19023 3352
rect 18967 3284 18978 3318
rect 19012 3284 19023 3318
rect 18967 3250 19023 3284
rect 18967 3216 18978 3250
rect 19012 3216 19023 3250
rect 18967 3182 19023 3216
rect 18967 3148 18978 3182
rect 19012 3148 19023 3182
rect 18967 3078 19023 3148
rect 19123 4066 19179 4078
rect 19123 4032 19134 4066
rect 19168 4032 19179 4066
rect 19123 3998 19179 4032
rect 19123 3964 19134 3998
rect 19168 3964 19179 3998
rect 19123 3930 19179 3964
rect 19123 3896 19134 3930
rect 19168 3896 19179 3930
rect 19123 3862 19179 3896
rect 19123 3828 19134 3862
rect 19168 3828 19179 3862
rect 19123 3794 19179 3828
rect 19123 3760 19134 3794
rect 19168 3760 19179 3794
rect 19123 3726 19179 3760
rect 19123 3692 19134 3726
rect 19168 3692 19179 3726
rect 19123 3658 19179 3692
rect 19123 3624 19134 3658
rect 19168 3624 19179 3658
rect 19123 3590 19179 3624
rect 19123 3556 19134 3590
rect 19168 3556 19179 3590
rect 19123 3522 19179 3556
rect 19123 3488 19134 3522
rect 19168 3488 19179 3522
rect 19123 3454 19179 3488
rect 19123 3420 19134 3454
rect 19168 3420 19179 3454
rect 19123 3386 19179 3420
rect 19123 3352 19134 3386
rect 19168 3352 19179 3386
rect 19123 3318 19179 3352
rect 19123 3284 19134 3318
rect 19168 3284 19179 3318
rect 19123 3250 19179 3284
rect 19123 3216 19134 3250
rect 19168 3216 19179 3250
rect 19123 3182 19179 3216
rect 19123 3148 19134 3182
rect 19168 3148 19179 3182
rect 19123 3078 19179 3148
rect 19279 4066 19335 4078
rect 19279 4032 19290 4066
rect 19324 4032 19335 4066
rect 19279 3998 19335 4032
rect 19279 3964 19290 3998
rect 19324 3964 19335 3998
rect 19279 3930 19335 3964
rect 19279 3896 19290 3930
rect 19324 3896 19335 3930
rect 19279 3862 19335 3896
rect 19279 3828 19290 3862
rect 19324 3828 19335 3862
rect 19279 3794 19335 3828
rect 19279 3760 19290 3794
rect 19324 3760 19335 3794
rect 19279 3726 19335 3760
rect 19279 3692 19290 3726
rect 19324 3692 19335 3726
rect 19279 3658 19335 3692
rect 19279 3624 19290 3658
rect 19324 3624 19335 3658
rect 19279 3590 19335 3624
rect 19279 3556 19290 3590
rect 19324 3556 19335 3590
rect 19279 3522 19335 3556
rect 19279 3488 19290 3522
rect 19324 3488 19335 3522
rect 19279 3454 19335 3488
rect 19279 3420 19290 3454
rect 19324 3420 19335 3454
rect 19279 3386 19335 3420
rect 19279 3352 19290 3386
rect 19324 3352 19335 3386
rect 19279 3318 19335 3352
rect 19279 3284 19290 3318
rect 19324 3284 19335 3318
rect 19279 3250 19335 3284
rect 19279 3216 19290 3250
rect 19324 3216 19335 3250
rect 19279 3182 19335 3216
rect 19279 3148 19290 3182
rect 19324 3148 19335 3182
rect 19279 3078 19335 3148
rect 19435 4066 19488 4078
rect 19435 4032 19446 4066
rect 19480 4032 19488 4066
rect 19435 3998 19488 4032
rect 19435 3964 19446 3998
rect 19480 3964 19488 3998
rect 19435 3930 19488 3964
rect 19435 3896 19446 3930
rect 19480 3896 19488 3930
rect 19435 3862 19488 3896
rect 19435 3828 19446 3862
rect 19480 3828 19488 3862
rect 19435 3794 19488 3828
rect 19435 3760 19446 3794
rect 19480 3760 19488 3794
rect 19435 3726 19488 3760
rect 19435 3692 19446 3726
rect 19480 3692 19488 3726
rect 19435 3658 19488 3692
rect 19435 3624 19446 3658
rect 19480 3624 19488 3658
rect 19435 3590 19488 3624
rect 19435 3556 19446 3590
rect 19480 3556 19488 3590
rect 19435 3522 19488 3556
rect 19435 3488 19446 3522
rect 19480 3488 19488 3522
rect 19435 3454 19488 3488
rect 19435 3420 19446 3454
rect 19480 3420 19488 3454
rect 19435 3386 19488 3420
rect 19435 3352 19446 3386
rect 19480 3352 19488 3386
rect 19435 3318 19488 3352
rect 19435 3284 19446 3318
rect 19480 3284 19488 3318
rect 19435 3250 19488 3284
rect 19435 3216 19446 3250
rect 19480 3216 19488 3250
rect 19435 3182 19488 3216
rect 19435 3148 19446 3182
rect 19480 3148 19488 3182
rect 19435 3078 19488 3148
rect 19548 4066 19601 4078
rect 19548 4032 19556 4066
rect 19590 4032 19601 4066
rect 19548 3998 19601 4032
rect 19548 3964 19556 3998
rect 19590 3964 19601 3998
rect 19548 3930 19601 3964
rect 19548 3896 19556 3930
rect 19590 3896 19601 3930
rect 19548 3862 19601 3896
rect 19548 3828 19556 3862
rect 19590 3828 19601 3862
rect 19548 3794 19601 3828
rect 19548 3760 19556 3794
rect 19590 3760 19601 3794
rect 19548 3726 19601 3760
rect 19548 3692 19556 3726
rect 19590 3692 19601 3726
rect 19548 3658 19601 3692
rect 19548 3624 19556 3658
rect 19590 3624 19601 3658
rect 19548 3590 19601 3624
rect 19548 3556 19556 3590
rect 19590 3556 19601 3590
rect 19548 3522 19601 3556
rect 19548 3488 19556 3522
rect 19590 3488 19601 3522
rect 19548 3454 19601 3488
rect 19548 3420 19556 3454
rect 19590 3420 19601 3454
rect 19548 3386 19601 3420
rect 19548 3352 19556 3386
rect 19590 3352 19601 3386
rect 19548 3318 19601 3352
rect 19548 3284 19556 3318
rect 19590 3284 19601 3318
rect 19548 3250 19601 3284
rect 19548 3216 19556 3250
rect 19590 3216 19601 3250
rect 19548 3182 19601 3216
rect 19548 3148 19556 3182
rect 19590 3148 19601 3182
rect 19548 3078 19601 3148
rect 19701 4066 19757 4078
rect 19701 4032 19712 4066
rect 19746 4032 19757 4066
rect 19701 3998 19757 4032
rect 19701 3964 19712 3998
rect 19746 3964 19757 3998
rect 19701 3930 19757 3964
rect 19701 3896 19712 3930
rect 19746 3896 19757 3930
rect 19701 3862 19757 3896
rect 19701 3828 19712 3862
rect 19746 3828 19757 3862
rect 19701 3794 19757 3828
rect 19701 3760 19712 3794
rect 19746 3760 19757 3794
rect 19701 3726 19757 3760
rect 19701 3692 19712 3726
rect 19746 3692 19757 3726
rect 19701 3658 19757 3692
rect 19701 3624 19712 3658
rect 19746 3624 19757 3658
rect 19701 3590 19757 3624
rect 19701 3556 19712 3590
rect 19746 3556 19757 3590
rect 19701 3522 19757 3556
rect 19701 3488 19712 3522
rect 19746 3488 19757 3522
rect 19701 3454 19757 3488
rect 19701 3420 19712 3454
rect 19746 3420 19757 3454
rect 19701 3386 19757 3420
rect 19701 3352 19712 3386
rect 19746 3352 19757 3386
rect 19701 3318 19757 3352
rect 19701 3284 19712 3318
rect 19746 3284 19757 3318
rect 19701 3250 19757 3284
rect 19701 3216 19712 3250
rect 19746 3216 19757 3250
rect 19701 3182 19757 3216
rect 19701 3148 19712 3182
rect 19746 3148 19757 3182
rect 19701 3078 19757 3148
rect 19857 4066 19910 4078
rect 19857 4032 19868 4066
rect 19902 4032 19910 4066
rect 19857 3998 19910 4032
rect 19857 3964 19868 3998
rect 19902 3964 19910 3998
rect 19857 3930 19910 3964
rect 19857 3896 19868 3930
rect 19902 3896 19910 3930
rect 19857 3862 19910 3896
rect 19857 3828 19868 3862
rect 19902 3828 19910 3862
rect 19857 3794 19910 3828
rect 19857 3760 19868 3794
rect 19902 3760 19910 3794
rect 19857 3726 19910 3760
rect 19857 3692 19868 3726
rect 19902 3692 19910 3726
rect 19857 3658 19910 3692
rect 19857 3624 19868 3658
rect 19902 3624 19910 3658
rect 19857 3590 19910 3624
rect 19857 3556 19868 3590
rect 19902 3556 19910 3590
rect 19857 3522 19910 3556
rect 19857 3488 19868 3522
rect 19902 3488 19910 3522
rect 19857 3454 19910 3488
rect 19857 3420 19868 3454
rect 19902 3420 19910 3454
rect 19857 3386 19910 3420
rect 19857 3352 19868 3386
rect 19902 3352 19910 3386
rect 19857 3318 19910 3352
rect 19857 3284 19868 3318
rect 19902 3284 19910 3318
rect 19857 3250 19910 3284
rect 19857 3216 19868 3250
rect 19902 3216 19910 3250
rect 19857 3182 19910 3216
rect 19857 3148 19868 3182
rect 19902 3148 19910 3182
rect 19857 3078 19910 3148
<< mvndiffc >>
rect 12128 5469 12162 5503
rect 12128 5401 12162 5435
rect 12128 5333 12162 5367
rect 12128 5265 12162 5299
rect 12128 5197 12162 5231
rect 12128 5129 12162 5163
rect 12128 5061 12162 5095
rect 12128 4993 12162 5027
rect 12128 4925 12162 4959
rect 12128 4857 12162 4891
rect 11538 4795 11572 4829
rect 11606 4795 11640 4829
rect 11674 4795 11708 4829
rect 11742 4795 11776 4829
rect 11810 4795 11844 4829
rect 11878 4795 11912 4829
rect 11946 4795 11980 4829
rect 12014 4795 12048 4829
rect 12128 4789 12162 4823
rect 12128 4721 12162 4755
rect 11538 4639 11572 4673
rect 11606 4639 11640 4673
rect 11674 4639 11708 4673
rect 11742 4639 11776 4673
rect 11810 4639 11844 4673
rect 11878 4639 11912 4673
rect 11946 4639 11980 4673
rect 12014 4639 12048 4673
rect 12128 4653 12162 4687
rect 12128 4585 12162 4619
rect 12304 5469 12338 5503
rect 12304 5401 12338 5435
rect 12304 5333 12338 5367
rect 12304 5265 12338 5299
rect 12304 5197 12338 5231
rect 12304 5129 12338 5163
rect 12304 5061 12338 5095
rect 12304 4993 12338 5027
rect 12304 4925 12338 4959
rect 12304 4857 12338 4891
rect 12304 4789 12338 4823
rect 12418 4815 12452 4849
rect 12486 4815 12520 4849
rect 12554 4815 12588 4849
rect 12622 4815 12656 4849
rect 12690 4815 12724 4849
rect 12758 4815 12792 4849
rect 12826 4815 12860 4849
rect 12894 4815 12928 4849
rect 12962 4815 12996 4849
rect 13030 4815 13064 4849
rect 13098 4815 13132 4849
rect 13166 4815 13200 4849
rect 13234 4815 13268 4849
rect 13302 4815 13336 4849
rect 12304 4721 12338 4755
rect 12304 4653 12338 4687
rect 12418 4639 12452 4673
rect 12486 4639 12520 4673
rect 12554 4639 12588 4673
rect 12622 4639 12656 4673
rect 12690 4639 12724 4673
rect 12758 4639 12792 4673
rect 12826 4639 12860 4673
rect 12894 4639 12928 4673
rect 12962 4639 12996 4673
rect 13030 4639 13064 4673
rect 13098 4639 13132 4673
rect 13166 4639 13200 4673
rect 13234 4639 13268 4673
rect 13302 4639 13336 4673
rect 12304 4585 12338 4619
rect 11536 4459 11570 4493
rect 11536 4391 11570 4425
rect 11536 4323 11570 4357
rect 11792 4459 11826 4493
rect 11792 4391 11826 4425
rect 11792 4323 11826 4357
rect 12048 4459 12082 4493
rect 12048 4391 12082 4425
rect 12048 4323 12082 4357
rect 12304 4459 12338 4493
rect 12304 4391 12338 4425
rect 12304 4323 12338 4357
rect 12560 4459 12594 4493
rect 12560 4391 12594 4425
rect 12560 4323 12594 4357
rect 12736 4459 12770 4493
rect 12736 4391 12770 4425
rect 12736 4323 12770 4357
rect 12912 4459 12946 4493
rect 12912 4391 12946 4425
rect 12912 4323 12946 4357
rect 13088 4459 13122 4493
rect 13088 4391 13122 4425
rect 13088 4323 13122 4357
rect 13264 4459 13298 4493
rect 13264 4391 13298 4425
rect 13264 4323 13298 4357
rect 13440 4459 13474 4493
rect 13440 4391 13474 4425
rect 13440 4323 13474 4357
rect 12472 4036 12506 4070
rect 12616 4036 12650 4070
rect 12472 3180 12506 3214
rect 12616 3180 12650 3214
<< mvpdiffc >>
rect 7369 6689 7403 6723
rect 7369 6621 7403 6655
rect 7369 6553 7403 6587
rect 7369 6485 7403 6519
rect 7369 6417 7403 6451
rect 7369 6349 7403 6383
rect 7369 6281 7403 6315
rect 7369 6213 7403 6247
rect 7369 6145 7403 6179
rect 7369 6077 7403 6111
rect 7369 6009 7403 6043
rect 7369 5941 7403 5975
rect 7369 5873 7403 5907
rect 7369 5805 7403 5839
rect 7369 5737 7403 5771
rect 7369 5669 7403 5703
rect 7369 5601 7403 5635
rect 7369 5533 7403 5567
rect 7369 5465 7403 5499
rect 7369 5397 7403 5431
rect 7369 5329 7403 5363
rect 7369 5261 7403 5295
rect 7369 5193 7403 5227
rect 7369 5125 7403 5159
rect 7369 5057 7403 5091
rect 7369 4989 7403 5023
rect 7369 4921 7403 4955
rect 7369 4853 7403 4887
rect 7369 4785 7403 4819
rect 7525 6689 7559 6723
rect 7525 6621 7559 6655
rect 7525 6553 7559 6587
rect 7525 6485 7559 6519
rect 7525 6417 7559 6451
rect 7525 6349 7559 6383
rect 7525 6281 7559 6315
rect 7525 6213 7559 6247
rect 7525 6145 7559 6179
rect 7525 6077 7559 6111
rect 7525 6009 7559 6043
rect 7525 5941 7559 5975
rect 7525 5873 7559 5907
rect 7525 5805 7559 5839
rect 7525 5737 7559 5771
rect 7525 5669 7559 5703
rect 7525 5601 7559 5635
rect 7525 5533 7559 5567
rect 7525 5465 7559 5499
rect 7525 5397 7559 5431
rect 7525 5329 7559 5363
rect 7525 5261 7559 5295
rect 7525 5193 7559 5227
rect 7525 5125 7559 5159
rect 7525 5057 7559 5091
rect 7525 4989 7559 5023
rect 7525 4921 7559 4955
rect 7525 4853 7559 4887
rect 7525 4785 7559 4819
rect 7681 6689 7715 6723
rect 7681 6621 7715 6655
rect 7681 6553 7715 6587
rect 7681 6485 7715 6519
rect 7681 6417 7715 6451
rect 7681 6349 7715 6383
rect 7681 6281 7715 6315
rect 7681 6213 7715 6247
rect 7681 6145 7715 6179
rect 7681 6077 7715 6111
rect 7681 6009 7715 6043
rect 7681 5941 7715 5975
rect 7681 5873 7715 5907
rect 7681 5805 7715 5839
rect 7681 5737 7715 5771
rect 7681 5669 7715 5703
rect 7681 5601 7715 5635
rect 7681 5533 7715 5567
rect 7681 5465 7715 5499
rect 7681 5397 7715 5431
rect 7681 5329 7715 5363
rect 7681 5261 7715 5295
rect 7681 5193 7715 5227
rect 7681 5125 7715 5159
rect 7681 5057 7715 5091
rect 7681 4989 7715 5023
rect 7681 4921 7715 4955
rect 7681 4853 7715 4887
rect 7681 4785 7715 4819
rect 7837 6689 7871 6723
rect 7837 6621 7871 6655
rect 7837 6553 7871 6587
rect 7837 6485 7871 6519
rect 7837 6417 7871 6451
rect 7837 6349 7871 6383
rect 7837 6281 7871 6315
rect 7837 6213 7871 6247
rect 7837 6145 7871 6179
rect 7837 6077 7871 6111
rect 7837 6009 7871 6043
rect 7837 5941 7871 5975
rect 7837 5873 7871 5907
rect 7837 5805 7871 5839
rect 7837 5737 7871 5771
rect 7837 5669 7871 5703
rect 7837 5601 7871 5635
rect 7837 5533 7871 5567
rect 7837 5465 7871 5499
rect 7837 5397 7871 5431
rect 7837 5329 7871 5363
rect 7837 5261 7871 5295
rect 7837 5193 7871 5227
rect 7837 5125 7871 5159
rect 7837 5057 7871 5091
rect 7837 4989 7871 5023
rect 7837 4921 7871 4955
rect 7837 4853 7871 4887
rect 7837 4785 7871 4819
rect 7993 6689 8027 6723
rect 7993 6621 8027 6655
rect 7993 6553 8027 6587
rect 7993 6485 8027 6519
rect 7993 6417 8027 6451
rect 7993 6349 8027 6383
rect 7993 6281 8027 6315
rect 7993 6213 8027 6247
rect 7993 6145 8027 6179
rect 7993 6077 8027 6111
rect 7993 6009 8027 6043
rect 7993 5941 8027 5975
rect 7993 5873 8027 5907
rect 7993 5805 8027 5839
rect 7993 5737 8027 5771
rect 7993 5669 8027 5703
rect 7993 5601 8027 5635
rect 7993 5533 8027 5567
rect 7993 5465 8027 5499
rect 7993 5397 8027 5431
rect 7993 5329 8027 5363
rect 7993 5261 8027 5295
rect 7993 5193 8027 5227
rect 7993 5125 8027 5159
rect 7993 5057 8027 5091
rect 7993 4989 8027 5023
rect 7993 4921 8027 4955
rect 7993 4853 8027 4887
rect 7993 4785 8027 4819
rect 7519 4314 7553 4348
rect 7519 4246 7553 4280
rect 7519 4178 7553 4212
rect 7519 4110 7553 4144
rect 7519 4042 7553 4076
rect 7519 3974 7553 4008
rect 7519 3906 7553 3940
rect 7519 3838 7553 3872
rect 7519 3770 7553 3804
rect 7519 3702 7553 3736
rect 7519 3634 7553 3668
rect 7519 3566 7553 3600
rect 7519 3498 7553 3532
rect 7519 3430 7553 3464
rect 7519 3362 7553 3396
rect 7519 3294 7553 3328
rect 7519 3226 7553 3260
rect 7519 3158 7553 3192
rect 7519 3090 7553 3124
rect 7519 3022 7553 3056
rect 7675 4314 7709 4348
rect 7675 4246 7709 4280
rect 7675 4178 7709 4212
rect 7675 4110 7709 4144
rect 7675 4042 7709 4076
rect 7675 3974 7709 4008
rect 7675 3906 7709 3940
rect 7675 3838 7709 3872
rect 7675 3770 7709 3804
rect 7675 3702 7709 3736
rect 7675 3634 7709 3668
rect 7675 3566 7709 3600
rect 7675 3498 7709 3532
rect 7675 3430 7709 3464
rect 7675 3362 7709 3396
rect 7675 3294 7709 3328
rect 7675 3226 7709 3260
rect 7675 3158 7709 3192
rect 7675 3090 7709 3124
rect 7675 3022 7709 3056
rect 7831 4314 7865 4348
rect 7831 4246 7865 4280
rect 7831 4178 7865 4212
rect 7831 4110 7865 4144
rect 7831 4042 7865 4076
rect 7831 3974 7865 4008
rect 7831 3906 7865 3940
rect 7831 3838 7865 3872
rect 7831 3770 7865 3804
rect 7831 3702 7865 3736
rect 7831 3634 7865 3668
rect 7831 3566 7865 3600
rect 7831 3498 7865 3532
rect 7831 3430 7865 3464
rect 7831 3362 7865 3396
rect 7831 3294 7865 3328
rect 7831 3226 7865 3260
rect 7831 3158 7865 3192
rect 7831 3090 7865 3124
rect 7831 3022 7865 3056
rect 7987 4314 8021 4348
rect 7987 4246 8021 4280
rect 7987 4178 8021 4212
rect 17634 4210 17668 4244
rect 19290 4210 19324 4244
rect 7987 4110 8021 4144
rect 7987 4042 8021 4076
rect 7987 3974 8021 4008
rect 7987 3906 8021 3940
rect 7987 3838 8021 3872
rect 7987 3770 8021 3804
rect 7987 3702 8021 3736
rect 7987 3634 8021 3668
rect 7987 3566 8021 3600
rect 7987 3498 8021 3532
rect 7987 3430 8021 3464
rect 7987 3362 8021 3396
rect 7987 3294 8021 3328
rect 7987 3226 8021 3260
rect 12944 4036 12978 4070
rect 13202 4027 13236 4061
rect 7987 3158 8021 3192
rect 13202 3959 13236 3993
rect 13202 3891 13236 3925
rect 13358 4027 13392 4061
rect 13358 3959 13392 3993
rect 13358 3891 13392 3925
rect 13514 4027 13548 4061
rect 13514 3959 13548 3993
rect 13514 3891 13548 3925
rect 7987 3090 8021 3124
rect 12944 3180 12978 3214
rect 13710 4032 13744 4066
rect 13710 3964 13744 3998
rect 13710 3896 13744 3930
rect 13710 3828 13744 3862
rect 13710 3760 13744 3794
rect 13710 3692 13744 3726
rect 13710 3624 13744 3658
rect 13710 3556 13744 3590
rect 13710 3488 13744 3522
rect 13710 3420 13744 3454
rect 13710 3352 13744 3386
rect 13710 3284 13744 3318
rect 13710 3216 13744 3250
rect 13710 3148 13744 3182
rect 13866 4032 13900 4066
rect 13866 3964 13900 3998
rect 13866 3896 13900 3930
rect 13866 3828 13900 3862
rect 13866 3760 13900 3794
rect 13866 3692 13900 3726
rect 13866 3624 13900 3658
rect 13866 3556 13900 3590
rect 13866 3488 13900 3522
rect 13866 3420 13900 3454
rect 13866 3352 13900 3386
rect 13866 3284 13900 3318
rect 13866 3216 13900 3250
rect 13866 3148 13900 3182
rect 14022 4032 14056 4066
rect 14022 3964 14056 3998
rect 14022 3896 14056 3930
rect 14022 3828 14056 3862
rect 14022 3760 14056 3794
rect 14022 3692 14056 3726
rect 14022 3624 14056 3658
rect 14022 3556 14056 3590
rect 14022 3488 14056 3522
rect 14022 3420 14056 3454
rect 14022 3352 14056 3386
rect 14022 3284 14056 3318
rect 14022 3216 14056 3250
rect 14022 3148 14056 3182
rect 14178 4032 14212 4066
rect 14178 3964 14212 3998
rect 14178 3896 14212 3930
rect 14178 3828 14212 3862
rect 14178 3760 14212 3794
rect 14178 3692 14212 3726
rect 14178 3624 14212 3658
rect 14178 3556 14212 3590
rect 14178 3488 14212 3522
rect 14178 3420 14212 3454
rect 14178 3352 14212 3386
rect 14178 3284 14212 3318
rect 14178 3216 14212 3250
rect 14178 3148 14212 3182
rect 14334 4032 14368 4066
rect 14334 3964 14368 3998
rect 14334 3896 14368 3930
rect 14334 3828 14368 3862
rect 14334 3760 14368 3794
rect 14334 3692 14368 3726
rect 14334 3624 14368 3658
rect 14334 3556 14368 3590
rect 14334 3488 14368 3522
rect 14334 3420 14368 3454
rect 14334 3352 14368 3386
rect 14334 3284 14368 3318
rect 14334 3216 14368 3250
rect 14334 3148 14368 3182
rect 14490 4032 14524 4066
rect 14490 3964 14524 3998
rect 14490 3896 14524 3930
rect 14490 3828 14524 3862
rect 14490 3760 14524 3794
rect 14490 3692 14524 3726
rect 14490 3624 14524 3658
rect 14490 3556 14524 3590
rect 14490 3488 14524 3522
rect 14490 3420 14524 3454
rect 14490 3352 14524 3386
rect 14490 3284 14524 3318
rect 14490 3216 14524 3250
rect 14490 3148 14524 3182
rect 14646 4032 14680 4066
rect 14646 3964 14680 3998
rect 14646 3896 14680 3930
rect 14646 3828 14680 3862
rect 14646 3760 14680 3794
rect 14646 3692 14680 3726
rect 14646 3624 14680 3658
rect 14646 3556 14680 3590
rect 14646 3488 14680 3522
rect 14646 3420 14680 3454
rect 14646 3352 14680 3386
rect 14646 3284 14680 3318
rect 14646 3216 14680 3250
rect 14646 3148 14680 3182
rect 14802 4032 14836 4066
rect 14802 3964 14836 3998
rect 14802 3896 14836 3930
rect 14802 3828 14836 3862
rect 14802 3760 14836 3794
rect 14802 3692 14836 3726
rect 14802 3624 14836 3658
rect 14802 3556 14836 3590
rect 14802 3488 14836 3522
rect 14802 3420 14836 3454
rect 14802 3352 14836 3386
rect 14802 3284 14836 3318
rect 14802 3216 14836 3250
rect 14802 3148 14836 3182
rect 14958 4032 14992 4066
rect 14958 3964 14992 3998
rect 14958 3896 14992 3930
rect 14958 3828 14992 3862
rect 14958 3760 14992 3794
rect 14958 3692 14992 3726
rect 14958 3624 14992 3658
rect 14958 3556 14992 3590
rect 14958 3488 14992 3522
rect 14958 3420 14992 3454
rect 14958 3352 14992 3386
rect 14958 3284 14992 3318
rect 14958 3216 14992 3250
rect 14958 3148 14992 3182
rect 15114 4032 15148 4066
rect 15114 3964 15148 3998
rect 15114 3896 15148 3930
rect 15114 3828 15148 3862
rect 15114 3760 15148 3794
rect 15114 3692 15148 3726
rect 15114 3624 15148 3658
rect 15114 3556 15148 3590
rect 15114 3488 15148 3522
rect 15114 3420 15148 3454
rect 15114 3352 15148 3386
rect 15114 3284 15148 3318
rect 15114 3216 15148 3250
rect 15114 3148 15148 3182
rect 15310 3982 15344 4016
rect 15310 3914 15344 3948
rect 15310 3846 15344 3880
rect 15310 3778 15344 3812
rect 15310 3710 15344 3744
rect 15310 3642 15344 3676
rect 15310 3574 15344 3608
rect 15310 3506 15344 3540
rect 15310 3438 15344 3472
rect 15310 3370 15344 3404
rect 15310 3302 15344 3336
rect 15310 3234 15344 3268
rect 15310 3166 15344 3200
rect 15310 3098 15344 3132
rect 7987 3022 8021 3056
rect 15466 3982 15500 4016
rect 15466 3914 15500 3948
rect 15466 3846 15500 3880
rect 15466 3778 15500 3812
rect 15466 3710 15500 3744
rect 15466 3642 15500 3676
rect 15466 3574 15500 3608
rect 15466 3506 15500 3540
rect 15466 3438 15500 3472
rect 15466 3370 15500 3404
rect 15466 3302 15500 3336
rect 15466 3234 15500 3268
rect 15466 3166 15500 3200
rect 15466 3098 15500 3132
rect 15622 3982 15656 4016
rect 15622 3914 15656 3948
rect 15622 3846 15656 3880
rect 15622 3778 15656 3812
rect 15622 3710 15656 3744
rect 15622 3642 15656 3676
rect 15622 3574 15656 3608
rect 15622 3506 15656 3540
rect 15622 3438 15656 3472
rect 15622 3370 15656 3404
rect 15622 3302 15656 3336
rect 15622 3234 15656 3268
rect 15622 3166 15656 3200
rect 15622 3098 15656 3132
rect 15778 3982 15812 4016
rect 15778 3914 15812 3948
rect 15778 3846 15812 3880
rect 15778 3778 15812 3812
rect 15778 3710 15812 3744
rect 15778 3642 15812 3676
rect 15778 3574 15812 3608
rect 15778 3506 15812 3540
rect 15778 3438 15812 3472
rect 15778 3370 15812 3404
rect 15778 3302 15812 3336
rect 15778 3234 15812 3268
rect 15778 3166 15812 3200
rect 15778 3098 15812 3132
rect 15934 3982 15968 4016
rect 15934 3914 15968 3948
rect 15934 3846 15968 3880
rect 15934 3778 15968 3812
rect 15934 3710 15968 3744
rect 15934 3642 15968 3676
rect 15934 3574 15968 3608
rect 15934 3506 15968 3540
rect 15934 3438 15968 3472
rect 15934 3370 15968 3404
rect 15934 3302 15968 3336
rect 15934 3234 15968 3268
rect 15934 3166 15968 3200
rect 15934 3098 15968 3132
rect 16090 3982 16124 4016
rect 16090 3914 16124 3948
rect 16090 3846 16124 3880
rect 16090 3778 16124 3812
rect 16090 3710 16124 3744
rect 16090 3642 16124 3676
rect 16090 3574 16124 3608
rect 16090 3506 16124 3540
rect 16090 3438 16124 3472
rect 16090 3370 16124 3404
rect 16090 3302 16124 3336
rect 16090 3234 16124 3268
rect 16090 3166 16124 3200
rect 16090 3098 16124 3132
rect 16246 3982 16280 4016
rect 16246 3914 16280 3948
rect 16246 3846 16280 3880
rect 16246 3778 16280 3812
rect 16246 3710 16280 3744
rect 16246 3642 16280 3676
rect 16246 3574 16280 3608
rect 16246 3506 16280 3540
rect 16246 3438 16280 3472
rect 16246 3370 16280 3404
rect 16246 3302 16280 3336
rect 16246 3234 16280 3268
rect 16246 3166 16280 3200
rect 16246 3098 16280 3132
rect 16402 3982 16436 4016
rect 16402 3914 16436 3948
rect 16402 3846 16436 3880
rect 16402 3778 16436 3812
rect 16402 3710 16436 3744
rect 16402 3642 16436 3676
rect 16402 3574 16436 3608
rect 16402 3506 16436 3540
rect 16402 3438 16436 3472
rect 16402 3370 16436 3404
rect 16402 3302 16436 3336
rect 16402 3234 16436 3268
rect 16402 3166 16436 3200
rect 16402 3098 16436 3132
rect 16558 3982 16592 4016
rect 16558 3914 16592 3948
rect 16558 3846 16592 3880
rect 16558 3778 16592 3812
rect 16558 3710 16592 3744
rect 16558 3642 16592 3676
rect 16558 3574 16592 3608
rect 16558 3506 16592 3540
rect 16558 3438 16592 3472
rect 16558 3370 16592 3404
rect 16558 3302 16592 3336
rect 16558 3234 16592 3268
rect 16558 3166 16592 3200
rect 16558 3098 16592 3132
rect 16754 4032 16788 4066
rect 16754 3964 16788 3998
rect 16754 3896 16788 3930
rect 16754 3828 16788 3862
rect 16754 3760 16788 3794
rect 16754 3692 16788 3726
rect 16754 3624 16788 3658
rect 16754 3556 16788 3590
rect 16754 3488 16788 3522
rect 16754 3420 16788 3454
rect 16754 3352 16788 3386
rect 16754 3284 16788 3318
rect 16754 3216 16788 3250
rect 16754 3148 16788 3182
rect 16910 4032 16944 4066
rect 16910 3964 16944 3998
rect 16910 3896 16944 3930
rect 16910 3828 16944 3862
rect 16910 3760 16944 3794
rect 16910 3692 16944 3726
rect 16910 3624 16944 3658
rect 16910 3556 16944 3590
rect 16910 3488 16944 3522
rect 16910 3420 16944 3454
rect 16910 3352 16944 3386
rect 16910 3284 16944 3318
rect 16910 3216 16944 3250
rect 16910 3148 16944 3182
rect 17066 4032 17100 4066
rect 17066 3964 17100 3998
rect 17066 3896 17100 3930
rect 17066 3828 17100 3862
rect 17066 3760 17100 3794
rect 17066 3692 17100 3726
rect 17066 3624 17100 3658
rect 17066 3556 17100 3590
rect 17066 3488 17100 3522
rect 17066 3420 17100 3454
rect 17066 3352 17100 3386
rect 17066 3284 17100 3318
rect 17066 3216 17100 3250
rect 17066 3148 17100 3182
rect 17222 4032 17256 4066
rect 17222 3964 17256 3998
rect 17222 3896 17256 3930
rect 17222 3828 17256 3862
rect 17222 3760 17256 3794
rect 17222 3692 17256 3726
rect 17222 3624 17256 3658
rect 17222 3556 17256 3590
rect 17222 3488 17256 3522
rect 17222 3420 17256 3454
rect 17222 3352 17256 3386
rect 17222 3284 17256 3318
rect 17222 3216 17256 3250
rect 17222 3148 17256 3182
rect 17378 4032 17412 4066
rect 17378 3964 17412 3998
rect 17378 3896 17412 3930
rect 17378 3828 17412 3862
rect 17378 3760 17412 3794
rect 17378 3692 17412 3726
rect 17378 3624 17412 3658
rect 17378 3556 17412 3590
rect 17378 3488 17412 3522
rect 17378 3420 17412 3454
rect 17378 3352 17412 3386
rect 17378 3284 17412 3318
rect 17378 3216 17412 3250
rect 17378 3148 17412 3182
rect 17534 4032 17568 4066
rect 17534 3964 17568 3998
rect 17534 3896 17568 3930
rect 17534 3828 17568 3862
rect 17534 3760 17568 3794
rect 17534 3692 17568 3726
rect 17534 3624 17568 3658
rect 17534 3556 17568 3590
rect 17534 3488 17568 3522
rect 17534 3420 17568 3454
rect 17534 3352 17568 3386
rect 17534 3284 17568 3318
rect 17534 3216 17568 3250
rect 17534 3148 17568 3182
rect 17690 4032 17724 4066
rect 17690 3964 17724 3998
rect 17690 3896 17724 3930
rect 17690 3828 17724 3862
rect 17690 3760 17724 3794
rect 17690 3692 17724 3726
rect 17690 3624 17724 3658
rect 17690 3556 17724 3590
rect 17690 3488 17724 3522
rect 17690 3420 17724 3454
rect 17690 3352 17724 3386
rect 17690 3284 17724 3318
rect 17690 3216 17724 3250
rect 17690 3148 17724 3182
rect 17846 4032 17880 4066
rect 17846 3964 17880 3998
rect 17846 3896 17880 3930
rect 17846 3828 17880 3862
rect 17846 3760 17880 3794
rect 17846 3692 17880 3726
rect 17846 3624 17880 3658
rect 17846 3556 17880 3590
rect 17846 3488 17880 3522
rect 17846 3420 17880 3454
rect 17846 3352 17880 3386
rect 17846 3284 17880 3318
rect 17846 3216 17880 3250
rect 17846 3148 17880 3182
rect 18002 4032 18036 4066
rect 18002 3964 18036 3998
rect 18002 3896 18036 3930
rect 18002 3828 18036 3862
rect 18002 3760 18036 3794
rect 18002 3692 18036 3726
rect 18002 3624 18036 3658
rect 18002 3556 18036 3590
rect 18002 3488 18036 3522
rect 18002 3420 18036 3454
rect 18002 3352 18036 3386
rect 18002 3284 18036 3318
rect 18002 3216 18036 3250
rect 18002 3148 18036 3182
rect 18198 4032 18232 4066
rect 18198 3964 18232 3998
rect 18198 3896 18232 3930
rect 18198 3828 18232 3862
rect 18198 3760 18232 3794
rect 18198 3692 18232 3726
rect 18198 3624 18232 3658
rect 18198 3556 18232 3590
rect 18198 3488 18232 3522
rect 18198 3420 18232 3454
rect 18198 3352 18232 3386
rect 18198 3284 18232 3318
rect 18198 3216 18232 3250
rect 18198 3148 18232 3182
rect 18354 4032 18388 4066
rect 18354 3964 18388 3998
rect 18354 3896 18388 3930
rect 18354 3828 18388 3862
rect 18354 3760 18388 3794
rect 18354 3692 18388 3726
rect 18354 3624 18388 3658
rect 18354 3556 18388 3590
rect 18354 3488 18388 3522
rect 18354 3420 18388 3454
rect 18354 3352 18388 3386
rect 18354 3284 18388 3318
rect 18354 3216 18388 3250
rect 18354 3148 18388 3182
rect 18510 4032 18544 4066
rect 18510 3964 18544 3998
rect 18510 3896 18544 3930
rect 18510 3828 18544 3862
rect 18510 3760 18544 3794
rect 18510 3692 18544 3726
rect 18510 3624 18544 3658
rect 18510 3556 18544 3590
rect 18510 3488 18544 3522
rect 18510 3420 18544 3454
rect 18510 3352 18544 3386
rect 18510 3284 18544 3318
rect 18510 3216 18544 3250
rect 18510 3148 18544 3182
rect 18666 4032 18700 4066
rect 18666 3964 18700 3998
rect 18666 3896 18700 3930
rect 18666 3828 18700 3862
rect 18666 3760 18700 3794
rect 18666 3692 18700 3726
rect 18666 3624 18700 3658
rect 18666 3556 18700 3590
rect 18666 3488 18700 3522
rect 18666 3420 18700 3454
rect 18666 3352 18700 3386
rect 18666 3284 18700 3318
rect 18666 3216 18700 3250
rect 18666 3148 18700 3182
rect 18822 4032 18856 4066
rect 18822 3964 18856 3998
rect 18822 3896 18856 3930
rect 18822 3828 18856 3862
rect 18822 3760 18856 3794
rect 18822 3692 18856 3726
rect 18822 3624 18856 3658
rect 18822 3556 18856 3590
rect 18822 3488 18856 3522
rect 18822 3420 18856 3454
rect 18822 3352 18856 3386
rect 18822 3284 18856 3318
rect 18822 3216 18856 3250
rect 18822 3148 18856 3182
rect 18978 4032 19012 4066
rect 18978 3964 19012 3998
rect 18978 3896 19012 3930
rect 18978 3828 19012 3862
rect 18978 3760 19012 3794
rect 18978 3692 19012 3726
rect 18978 3624 19012 3658
rect 18978 3556 19012 3590
rect 18978 3488 19012 3522
rect 18978 3420 19012 3454
rect 18978 3352 19012 3386
rect 18978 3284 19012 3318
rect 18978 3216 19012 3250
rect 18978 3148 19012 3182
rect 19134 4032 19168 4066
rect 19134 3964 19168 3998
rect 19134 3896 19168 3930
rect 19134 3828 19168 3862
rect 19134 3760 19168 3794
rect 19134 3692 19168 3726
rect 19134 3624 19168 3658
rect 19134 3556 19168 3590
rect 19134 3488 19168 3522
rect 19134 3420 19168 3454
rect 19134 3352 19168 3386
rect 19134 3284 19168 3318
rect 19134 3216 19168 3250
rect 19134 3148 19168 3182
rect 19290 4032 19324 4066
rect 19290 3964 19324 3998
rect 19290 3896 19324 3930
rect 19290 3828 19324 3862
rect 19290 3760 19324 3794
rect 19290 3692 19324 3726
rect 19290 3624 19324 3658
rect 19290 3556 19324 3590
rect 19290 3488 19324 3522
rect 19290 3420 19324 3454
rect 19290 3352 19324 3386
rect 19290 3284 19324 3318
rect 19290 3216 19324 3250
rect 19290 3148 19324 3182
rect 19446 4032 19480 4066
rect 19446 3964 19480 3998
rect 19446 3896 19480 3930
rect 19446 3828 19480 3862
rect 19446 3760 19480 3794
rect 19446 3692 19480 3726
rect 19446 3624 19480 3658
rect 19446 3556 19480 3590
rect 19446 3488 19480 3522
rect 19446 3420 19480 3454
rect 19446 3352 19480 3386
rect 19446 3284 19480 3318
rect 19446 3216 19480 3250
rect 19446 3148 19480 3182
rect 19556 4032 19590 4066
rect 19556 3964 19590 3998
rect 19556 3896 19590 3930
rect 19556 3828 19590 3862
rect 19556 3760 19590 3794
rect 19556 3692 19590 3726
rect 19556 3624 19590 3658
rect 19556 3556 19590 3590
rect 19556 3488 19590 3522
rect 19556 3420 19590 3454
rect 19556 3352 19590 3386
rect 19556 3284 19590 3318
rect 19556 3216 19590 3250
rect 19556 3148 19590 3182
rect 19712 4032 19746 4066
rect 19712 3964 19746 3998
rect 19712 3896 19746 3930
rect 19712 3828 19746 3862
rect 19712 3760 19746 3794
rect 19712 3692 19746 3726
rect 19712 3624 19746 3658
rect 19712 3556 19746 3590
rect 19712 3488 19746 3522
rect 19712 3420 19746 3454
rect 19712 3352 19746 3386
rect 19712 3284 19746 3318
rect 19712 3216 19746 3250
rect 19712 3148 19746 3182
rect 19868 4032 19902 4066
rect 19868 3964 19902 3998
rect 19868 3896 19902 3930
rect 19868 3828 19902 3862
rect 19868 3760 19902 3794
rect 19868 3692 19902 3726
rect 19868 3624 19902 3658
rect 19868 3556 19902 3590
rect 19868 3488 19902 3522
rect 19868 3420 19902 3454
rect 19868 3352 19902 3386
rect 19868 3284 19902 3318
rect 19868 3216 19902 3250
rect 19868 3148 19902 3182
<< mvnsubdiff >>
rect 12814 4035 12852 4078
rect 12814 4001 12816 4035
rect 12850 4001 12852 4035
rect 12814 3967 12852 4001
rect 12814 3933 12816 3967
rect 12850 3933 12852 3967
rect 12814 3899 12852 3933
rect 12814 3865 12816 3899
rect 12850 3865 12852 3899
rect 12814 3831 12852 3865
rect 12814 3797 12816 3831
rect 12850 3797 12852 3831
rect 12814 3763 12852 3797
rect 12814 3729 12816 3763
rect 12850 3729 12852 3763
rect 12814 3695 12852 3729
rect 12814 3661 12816 3695
rect 12850 3661 12852 3695
rect 12814 3627 12852 3661
rect 12814 3593 12816 3627
rect 12850 3593 12852 3627
rect 12814 3559 12852 3593
rect 12814 3525 12816 3559
rect 12850 3525 12852 3559
rect 12814 3491 12852 3525
rect 12814 3457 12816 3491
rect 12850 3457 12852 3491
rect 12814 3423 12852 3457
rect 12814 3389 12816 3423
rect 12850 3389 12852 3423
rect 12814 3355 12852 3389
rect 12814 3321 12816 3355
rect 12850 3321 12852 3355
rect 12814 3287 12852 3321
rect 12814 3253 12816 3287
rect 12850 3253 12852 3287
rect 12814 3219 12852 3253
rect 13610 4035 13648 4078
rect 13610 4001 13612 4035
rect 13646 4001 13648 4035
rect 13610 3967 13648 4001
rect 13610 3933 13612 3967
rect 13646 3933 13648 3967
rect 13610 3899 13648 3933
rect 13610 3865 13612 3899
rect 13646 3865 13648 3899
rect 13610 3831 13648 3865
rect 13610 3797 13612 3831
rect 13646 3797 13648 3831
rect 13610 3763 13648 3797
rect 13610 3729 13612 3763
rect 13646 3729 13648 3763
rect 13610 3695 13648 3729
rect 13610 3661 13612 3695
rect 13646 3661 13648 3695
rect 13610 3627 13648 3661
rect 13610 3593 13612 3627
rect 13646 3593 13648 3627
rect 13610 3559 13648 3593
rect 13610 3525 13612 3559
rect 13646 3525 13648 3559
rect 13610 3491 13648 3525
rect 13610 3457 13612 3491
rect 13646 3457 13648 3491
rect 13610 3423 13648 3457
rect 13610 3389 13612 3423
rect 13646 3389 13648 3423
rect 13610 3355 13648 3389
rect 13610 3321 13612 3355
rect 13646 3321 13648 3355
rect 13610 3287 13648 3321
rect 13610 3253 13612 3287
rect 13646 3253 13648 3287
rect 12814 3185 12816 3219
rect 12850 3185 12852 3219
rect 12814 3151 12852 3185
rect 13610 3219 13648 3253
rect 13610 3185 13612 3219
rect 13646 3185 13648 3219
rect 12814 3117 12816 3151
rect 12850 3117 12852 3151
rect 12814 3078 12852 3117
rect 13610 3151 13648 3185
rect 13610 3117 13612 3151
rect 13646 3117 13648 3151
rect 13610 3078 13648 3117
rect 15210 4035 15248 4078
rect 15210 4001 15212 4035
rect 15246 4001 15248 4035
rect 16654 4035 16692 4078
rect 15210 3967 15248 4001
rect 15210 3933 15212 3967
rect 15246 3933 15248 3967
rect 15210 3899 15248 3933
rect 15210 3865 15212 3899
rect 15246 3865 15248 3899
rect 15210 3831 15248 3865
rect 15210 3797 15212 3831
rect 15246 3797 15248 3831
rect 15210 3763 15248 3797
rect 15210 3729 15212 3763
rect 15246 3729 15248 3763
rect 15210 3695 15248 3729
rect 15210 3661 15212 3695
rect 15246 3661 15248 3695
rect 15210 3627 15248 3661
rect 15210 3593 15212 3627
rect 15246 3593 15248 3627
rect 15210 3559 15248 3593
rect 15210 3525 15212 3559
rect 15246 3525 15248 3559
rect 15210 3491 15248 3525
rect 15210 3457 15212 3491
rect 15246 3457 15248 3491
rect 15210 3423 15248 3457
rect 15210 3389 15212 3423
rect 15246 3389 15248 3423
rect 15210 3355 15248 3389
rect 15210 3321 15212 3355
rect 15246 3321 15248 3355
rect 15210 3287 15248 3321
rect 15210 3253 15212 3287
rect 15246 3253 15248 3287
rect 15210 3219 15248 3253
rect 15210 3185 15212 3219
rect 15246 3185 15248 3219
rect 15210 3151 15248 3185
rect 15210 3117 15212 3151
rect 15246 3117 15248 3151
rect 15210 3078 15248 3117
rect 16654 4001 16656 4035
rect 16690 4001 16692 4035
rect 16654 3967 16692 4001
rect 16654 3933 16656 3967
rect 16690 3933 16692 3967
rect 16654 3899 16692 3933
rect 16654 3865 16656 3899
rect 16690 3865 16692 3899
rect 16654 3831 16692 3865
rect 16654 3797 16656 3831
rect 16690 3797 16692 3831
rect 16654 3763 16692 3797
rect 16654 3729 16656 3763
rect 16690 3729 16692 3763
rect 16654 3695 16692 3729
rect 16654 3661 16656 3695
rect 16690 3661 16692 3695
rect 16654 3627 16692 3661
rect 16654 3593 16656 3627
rect 16690 3593 16692 3627
rect 16654 3559 16692 3593
rect 16654 3525 16656 3559
rect 16690 3525 16692 3559
rect 16654 3491 16692 3525
rect 16654 3457 16656 3491
rect 16690 3457 16692 3491
rect 16654 3423 16692 3457
rect 16654 3389 16656 3423
rect 16690 3389 16692 3423
rect 16654 3355 16692 3389
rect 16654 3321 16656 3355
rect 16690 3321 16692 3355
rect 16654 3287 16692 3321
rect 16654 3253 16656 3287
rect 16690 3253 16692 3287
rect 16654 3219 16692 3253
rect 16654 3185 16656 3219
rect 16690 3185 16692 3219
rect 16654 3151 16692 3185
rect 16654 3117 16656 3151
rect 16690 3117 16692 3151
rect 16654 3078 16692 3117
rect 18098 4035 18136 4078
rect 18098 4001 18100 4035
rect 18134 4001 18136 4035
rect 18098 3967 18136 4001
rect 18098 3933 18100 3967
rect 18134 3933 18136 3967
rect 18098 3899 18136 3933
rect 18098 3865 18100 3899
rect 18134 3865 18136 3899
rect 18098 3831 18136 3865
rect 18098 3797 18100 3831
rect 18134 3797 18136 3831
rect 18098 3763 18136 3797
rect 18098 3729 18100 3763
rect 18134 3729 18136 3763
rect 18098 3695 18136 3729
rect 18098 3661 18100 3695
rect 18134 3661 18136 3695
rect 18098 3627 18136 3661
rect 18098 3593 18100 3627
rect 18134 3593 18136 3627
rect 18098 3559 18136 3593
rect 18098 3525 18100 3559
rect 18134 3525 18136 3559
rect 18098 3491 18136 3525
rect 18098 3457 18100 3491
rect 18134 3457 18136 3491
rect 18098 3423 18136 3457
rect 18098 3389 18100 3423
rect 18134 3389 18136 3423
rect 18098 3355 18136 3389
rect 18098 3321 18100 3355
rect 18134 3321 18136 3355
rect 18098 3287 18136 3321
rect 18098 3253 18100 3287
rect 18134 3253 18136 3287
rect 18098 3219 18136 3253
rect 18098 3185 18100 3219
rect 18134 3185 18136 3219
rect 18098 3151 18136 3185
rect 18098 3117 18100 3151
rect 18134 3117 18136 3151
rect 18098 3078 18136 3117
rect 19964 3287 20002 3344
rect 19964 3253 19966 3287
rect 20000 3253 20002 3287
rect 19964 3219 20002 3253
rect 19964 3185 19966 3219
rect 20000 3185 20002 3219
rect 19964 3151 20002 3185
rect 19964 3117 19966 3151
rect 20000 3117 20002 3151
rect 19964 3083 20002 3117
rect 19964 3049 19966 3083
rect 20000 3049 20002 3083
rect 19964 3015 20002 3049
rect 19964 3012 19966 3015
rect 20000 3012 20002 3015
rect 19964 2912 20002 3012
<< mvnsubdiffcont >>
rect 12816 4001 12850 4035
rect 12816 3933 12850 3967
rect 12816 3865 12850 3899
rect 12816 3797 12850 3831
rect 12816 3729 12850 3763
rect 12816 3661 12850 3695
rect 12816 3593 12850 3627
rect 12816 3525 12850 3559
rect 12816 3457 12850 3491
rect 12816 3389 12850 3423
rect 12816 3321 12850 3355
rect 12816 3253 12850 3287
rect 13612 4001 13646 4035
rect 13612 3933 13646 3967
rect 13612 3865 13646 3899
rect 13612 3797 13646 3831
rect 13612 3729 13646 3763
rect 13612 3661 13646 3695
rect 13612 3593 13646 3627
rect 13612 3525 13646 3559
rect 13612 3457 13646 3491
rect 13612 3389 13646 3423
rect 13612 3321 13646 3355
rect 13612 3253 13646 3287
rect 12816 3185 12850 3219
rect 13612 3185 13646 3219
rect 12816 3117 12850 3151
rect 13612 3117 13646 3151
rect 15212 4001 15246 4035
rect 15212 3933 15246 3967
rect 15212 3865 15246 3899
rect 15212 3797 15246 3831
rect 15212 3729 15246 3763
rect 15212 3661 15246 3695
rect 15212 3593 15246 3627
rect 15212 3525 15246 3559
rect 15212 3457 15246 3491
rect 15212 3389 15246 3423
rect 15212 3321 15246 3355
rect 15212 3253 15246 3287
rect 15212 3185 15246 3219
rect 15212 3117 15246 3151
rect 16656 4001 16690 4035
rect 16656 3933 16690 3967
rect 16656 3865 16690 3899
rect 16656 3797 16690 3831
rect 16656 3729 16690 3763
rect 16656 3661 16690 3695
rect 16656 3593 16690 3627
rect 16656 3525 16690 3559
rect 16656 3457 16690 3491
rect 16656 3389 16690 3423
rect 16656 3321 16690 3355
rect 16656 3253 16690 3287
rect 16656 3185 16690 3219
rect 16656 3117 16690 3151
rect 18100 4001 18134 4035
rect 18100 3933 18134 3967
rect 18100 3865 18134 3899
rect 18100 3797 18134 3831
rect 18100 3729 18134 3763
rect 18100 3661 18134 3695
rect 18100 3593 18134 3627
rect 18100 3525 18134 3559
rect 18100 3457 18134 3491
rect 18100 3389 18134 3423
rect 18100 3321 18134 3355
rect 18100 3253 18134 3287
rect 18100 3185 18134 3219
rect 18100 3117 18134 3151
rect 19966 3253 20000 3287
rect 19966 3185 20000 3219
rect 19966 3117 20000 3151
rect 19966 3049 20000 3083
rect 19966 3012 20000 3015
<< poly >>
rect 7414 6773 7514 6805
rect 7570 6773 7670 6805
rect 7726 6773 7826 6805
rect 7882 6773 7982 6805
rect 12159 5655 12293 5671
rect 12159 5621 12175 5655
rect 12209 5621 12243 5655
rect 12277 5621 12293 5655
rect 12159 5599 12293 5621
rect 12173 5573 12293 5599
rect 11368 4784 11434 4786
rect 7414 4741 7514 4773
rect 7570 4741 7670 4773
rect 7414 4725 7670 4741
rect 7414 4691 7430 4725
rect 7464 4691 7525 4725
rect 7559 4691 7620 4725
rect 7654 4691 7670 4725
rect 7414 4675 7670 4691
rect 7726 4741 7826 4773
rect 7882 4741 7982 4773
rect 7726 4725 7982 4741
rect 7726 4691 7742 4725
rect 7776 4691 7837 4725
rect 7871 4691 7932 4725
rect 7966 4691 7982 4725
rect 7726 4675 7982 4691
rect 11368 4770 11460 4784
rect 11368 4736 11384 4770
rect 11418 4736 11460 4770
rect 11368 4702 11460 4736
rect 11368 4668 11384 4702
rect 11418 4684 11460 4702
rect 12060 4684 12086 4784
rect 11418 4668 11434 4684
rect 11368 4652 11434 4668
rect 12380 4684 12406 4804
rect 13406 4788 13504 4804
rect 13406 4754 13454 4788
rect 13488 4754 13504 4788
rect 13406 4720 13504 4754
rect 13406 4686 13454 4720
rect 13488 4686 13504 4720
rect 13406 4684 13504 4686
rect 13432 4670 13504 4684
rect 12770 4593 12904 4609
rect 12173 4547 12293 4573
rect 11581 4511 11781 4537
rect 11837 4511 12037 4537
rect 12093 4511 12293 4547
rect 12770 4559 12786 4593
rect 12820 4559 12854 4593
rect 12888 4559 12904 4593
rect 12770 4537 12904 4559
rect 13122 4593 13256 4609
rect 13122 4559 13138 4593
rect 13172 4559 13206 4593
rect 13240 4559 13256 4593
rect 13122 4537 13256 4559
rect 12349 4511 12549 4537
rect 12605 4511 12725 4537
rect 12781 4511 12901 4537
rect 12957 4511 13077 4537
rect 13133 4511 13253 4537
rect 13309 4511 13429 4537
rect 7564 4492 7976 4508
rect 7564 4458 7580 4492
rect 7614 4458 7649 4492
rect 7683 4458 7718 4492
rect 7752 4458 7787 4492
rect 7821 4458 7856 4492
rect 7890 4458 7926 4492
rect 7960 4458 7976 4492
rect 7564 4442 7976 4458
rect 7564 4410 7664 4442
rect 7720 4410 7820 4442
rect 7876 4410 7976 4442
rect 17679 4338 19279 4354
rect 11581 4285 11781 4311
rect 11837 4285 12037 4311
rect 12093 4285 12293 4311
rect 12349 4285 12549 4311
rect 11581 4263 12549 4285
rect 11581 4229 11606 4263
rect 11640 4229 11674 4263
rect 11708 4229 11742 4263
rect 11776 4229 11810 4263
rect 11844 4229 11878 4263
rect 11912 4229 11946 4263
rect 11980 4229 12014 4263
rect 12048 4229 12082 4263
rect 12116 4229 12150 4263
rect 12184 4229 12218 4263
rect 12252 4229 12286 4263
rect 12320 4229 12354 4263
rect 12388 4229 12549 4263
rect 11581 4213 12549 4229
rect 12605 4285 12725 4311
rect 12781 4285 12901 4311
rect 12957 4285 13077 4311
rect 13133 4285 13253 4311
rect 13309 4285 13429 4311
rect 12605 4263 12739 4285
rect 12605 4229 12621 4263
rect 12655 4229 12689 4263
rect 12723 4229 12739 4263
rect 12605 4213 12739 4229
rect 12957 4263 13091 4285
rect 12957 4229 12973 4263
rect 13007 4229 13041 4263
rect 13075 4229 13091 4263
rect 12957 4213 13091 4229
rect 13295 4263 13429 4285
rect 13295 4229 13311 4263
rect 13345 4229 13379 4263
rect 13413 4229 13429 4263
rect 17679 4304 17719 4338
rect 17753 4304 17787 4338
rect 17821 4304 17855 4338
rect 17889 4304 17923 4338
rect 17957 4304 17991 4338
rect 18025 4304 18059 4338
rect 18093 4304 18127 4338
rect 18161 4304 18195 4338
rect 18229 4304 18263 4338
rect 18297 4304 18331 4338
rect 18365 4304 18399 4338
rect 18433 4304 18467 4338
rect 18501 4304 18535 4338
rect 18569 4304 18603 4338
rect 18637 4304 18671 4338
rect 18705 4304 18739 4338
rect 18773 4304 18807 4338
rect 18841 4304 18875 4338
rect 18909 4304 18943 4338
rect 18977 4304 19011 4338
rect 19045 4304 19079 4338
rect 19113 4304 19147 4338
rect 19181 4304 19215 4338
rect 19249 4304 19279 4338
rect 17679 4256 19279 4304
rect 13295 4171 13429 4229
rect 13155 4155 13503 4171
rect 13155 4121 13171 4155
rect 13205 4121 13239 4155
rect 13273 4121 13307 4155
rect 13341 4121 13503 4155
rect 17679 4146 19279 4172
rect 19583 4160 19857 4176
rect 13155 4099 13503 4121
rect 19583 4126 19599 4160
rect 19633 4126 19667 4160
rect 19701 4126 19735 4160
rect 19769 4126 19803 4160
rect 19837 4126 19857 4160
rect 19583 4104 19857 4126
rect 12336 3982 12434 4025
rect 12336 3948 12352 3982
rect 12386 3948 12434 3982
rect 12336 3914 12434 3948
rect 12336 3880 12352 3914
rect 12386 3880 12434 3914
rect 12336 3846 12434 3880
rect 12336 3812 12352 3846
rect 12386 3812 12434 3846
rect 12336 3778 12434 3812
rect 12336 3744 12352 3778
rect 12386 3744 12434 3778
rect 12336 3710 12434 3744
rect 12336 3676 12352 3710
rect 12386 3676 12434 3710
rect 12336 3642 12434 3676
rect 12336 3608 12352 3642
rect 12386 3608 12434 3642
rect 12336 3574 12434 3608
rect 12336 3540 12352 3574
rect 12386 3540 12434 3574
rect 12336 3506 12434 3540
rect 12336 3472 12352 3506
rect 12386 3472 12434 3506
rect 12336 3438 12434 3472
rect 12336 3404 12352 3438
rect 12386 3404 12434 3438
rect 12336 3370 12434 3404
rect 12336 3336 12352 3370
rect 12386 3336 12434 3370
rect 12336 3302 12434 3336
rect 12336 3268 12352 3302
rect 12386 3268 12434 3302
rect 12336 3225 12434 3268
rect 12518 3225 12578 4025
rect 12662 3225 12688 4025
rect 13247 4073 13347 4099
rect 13403 4073 13503 4099
rect 13755 4078 13855 4104
rect 13911 4078 14011 4104
rect 14067 4078 14167 4104
rect 14223 4078 14323 4104
rect 14379 4078 14479 4104
rect 14535 4078 14635 4104
rect 14691 4078 14791 4104
rect 14847 4078 14947 4104
rect 15003 4078 15103 4104
rect 16799 4078 16899 4104
rect 16955 4078 17055 4104
rect 17111 4078 17211 4104
rect 17267 4078 17367 4104
rect 17423 4078 17523 4104
rect 17579 4078 17679 4104
rect 17735 4078 17835 4104
rect 17891 4078 17991 4104
rect 18243 4078 18343 4104
rect 18399 4078 18499 4104
rect 18555 4078 18655 4104
rect 18711 4078 18811 4104
rect 18867 4078 18967 4104
rect 19023 4078 19123 4104
rect 19179 4078 19279 4104
rect 19335 4078 19435 4104
rect 19601 4078 19701 4104
rect 19757 4078 19857 4104
rect 12880 3225 12906 4025
rect 12990 4000 13088 4025
rect 12990 3966 13038 4000
rect 13072 3966 13088 4000
rect 12990 3928 13088 3966
rect 12990 3894 13038 3928
rect 13072 3894 13088 3928
rect 12990 3856 13088 3894
rect 12990 3822 13038 3856
rect 13072 3822 13088 3856
rect 13247 3847 13347 3873
rect 13403 3847 13503 3873
rect 12990 3784 13088 3822
rect 12990 3750 13038 3784
rect 13072 3750 13088 3784
rect 12990 3712 13088 3750
rect 12990 3678 13038 3712
rect 13072 3678 13088 3712
rect 12990 3640 13088 3678
rect 12990 3606 13038 3640
rect 13072 3606 13088 3640
rect 12990 3568 13088 3606
rect 12990 3534 13038 3568
rect 13072 3534 13088 3568
rect 12990 3496 13088 3534
rect 12990 3462 13038 3496
rect 13072 3462 13088 3496
rect 12990 3424 13088 3462
rect 12990 3390 13038 3424
rect 13072 3390 13088 3424
rect 12990 3352 13088 3390
rect 12990 3318 13038 3352
rect 13072 3318 13088 3352
rect 12990 3280 13088 3318
rect 12990 3246 13038 3280
rect 13072 3246 13088 3280
rect 12990 3225 13088 3246
rect 15355 4028 15455 4054
rect 15511 4028 15611 4054
rect 15667 4028 15767 4054
rect 15823 4028 15923 4054
rect 15979 4028 16079 4054
rect 16135 4028 16235 4054
rect 16291 4028 16391 4054
rect 16447 4028 16547 4054
rect 13755 3052 13855 3078
rect 13721 3030 13855 3052
rect 7564 2978 7664 3010
rect 7720 2978 7820 3010
rect 7876 2978 7976 3010
rect 13721 2996 13737 3030
rect 13771 2996 13805 3030
rect 13839 2996 13855 3030
rect 13721 2980 13855 2996
rect 13911 3052 14011 3078
rect 14067 3052 14167 3078
rect 14223 3052 14323 3078
rect 14379 3052 14479 3078
rect 14535 3052 14635 3078
rect 14691 3052 14791 3078
rect 14847 3052 14947 3078
rect 15003 3052 15103 3078
rect 13911 3030 15103 3052
rect 13911 2996 13944 3030
rect 13978 2996 14012 3030
rect 14046 2996 14080 3030
rect 14114 2996 14148 3030
rect 14182 2996 14216 3030
rect 14250 2996 14284 3030
rect 14318 2996 14352 3030
rect 14386 2996 14420 3030
rect 14454 2996 14488 3030
rect 14522 2996 14556 3030
rect 14590 2996 14624 3030
rect 14658 2996 14692 3030
rect 14726 2996 14760 3030
rect 14794 2996 14828 3030
rect 14862 2996 14896 3030
rect 14930 2996 14964 3030
rect 14998 2996 15032 3030
rect 15066 2996 15103 3030
rect 16799 3052 16899 3078
rect 16955 3052 17055 3078
rect 17111 3052 17211 3078
rect 17267 3052 17367 3078
rect 17423 3052 17523 3078
rect 17579 3052 17679 3078
rect 17735 3052 17835 3078
rect 17891 3052 17991 3078
rect 18243 3052 18343 3078
rect 18399 3052 18499 3078
rect 18555 3052 18655 3078
rect 18711 3052 18811 3078
rect 18867 3052 18967 3078
rect 19023 3052 19123 3078
rect 19179 3052 19279 3078
rect 19335 3052 19435 3078
rect 19601 3052 19701 3078
rect 19757 3052 19857 3078
rect 16799 3030 17991 3052
rect 13911 2980 15103 2996
rect 15355 3002 15455 3028
rect 15511 3002 15611 3028
rect 15667 3002 15767 3028
rect 15823 3002 15923 3028
rect 15979 3002 16079 3028
rect 16135 3002 16235 3028
rect 16291 3002 16391 3028
rect 16447 3002 16547 3028
rect 15355 2980 16547 3002
rect 16799 2996 16833 3030
rect 16867 2996 16901 3030
rect 16935 2996 16969 3030
rect 17003 2996 17037 3030
rect 17071 2996 17105 3030
rect 17139 2996 17173 3030
rect 17207 2996 17241 3030
rect 17275 2996 17309 3030
rect 17343 2996 17377 3030
rect 17411 2996 17445 3030
rect 17479 2996 17513 3030
rect 17547 2996 17581 3030
rect 17615 2996 17649 3030
rect 17683 2996 17717 3030
rect 17751 2996 17785 3030
rect 17819 2996 17853 3030
rect 17887 2996 17921 3030
rect 17955 2996 17991 3030
rect 16799 2980 17991 2996
rect 18244 3030 18811 3052
rect 18244 2996 18273 3030
rect 18307 2996 18341 3030
rect 18375 2996 18409 3030
rect 18443 2996 18477 3030
rect 18511 2996 18545 3030
rect 18579 2996 18613 3030
rect 18647 2996 18681 3030
rect 18715 2996 18749 3030
rect 18783 2996 18811 3030
rect 18244 2980 18811 2996
rect 18868 3030 19435 3052
rect 18868 2996 18897 3030
rect 18931 2996 18965 3030
rect 18999 2996 19033 3030
rect 19067 2996 19101 3030
rect 19135 2996 19169 3030
rect 19203 2996 19237 3030
rect 19271 2996 19305 3030
rect 19339 2996 19373 3030
rect 19407 2996 19435 3030
rect 18868 2980 19435 2996
rect 15355 2946 15389 2980
rect 15423 2946 15457 2980
rect 15491 2946 15525 2980
rect 15559 2946 15593 2980
rect 15627 2946 15661 2980
rect 15695 2946 15729 2980
rect 15763 2946 15797 2980
rect 15831 2946 15865 2980
rect 15899 2946 15933 2980
rect 15967 2946 16001 2980
rect 16035 2946 16069 2980
rect 16103 2946 16137 2980
rect 16171 2946 16205 2980
rect 16239 2946 16273 2980
rect 16307 2946 16341 2980
rect 16375 2946 16409 2980
rect 16443 2946 16477 2980
rect 16511 2946 16547 2980
rect 15355 2930 16547 2946
<< polycont >>
rect 12175 5621 12209 5655
rect 12243 5621 12277 5655
rect 7430 4691 7464 4725
rect 7525 4691 7559 4725
rect 7620 4691 7654 4725
rect 7742 4691 7776 4725
rect 7837 4691 7871 4725
rect 7932 4691 7966 4725
rect 11384 4736 11418 4770
rect 11384 4668 11418 4702
rect 13454 4754 13488 4788
rect 13454 4686 13488 4720
rect 12786 4559 12820 4593
rect 12854 4559 12888 4593
rect 13138 4559 13172 4593
rect 13206 4559 13240 4593
rect 7580 4458 7614 4492
rect 7649 4458 7683 4492
rect 7718 4458 7752 4492
rect 7787 4458 7821 4492
rect 7856 4458 7890 4492
rect 7926 4458 7960 4492
rect 11606 4229 11640 4263
rect 11674 4229 11708 4263
rect 11742 4229 11776 4263
rect 11810 4229 11844 4263
rect 11878 4229 11912 4263
rect 11946 4229 11980 4263
rect 12014 4229 12048 4263
rect 12082 4229 12116 4263
rect 12150 4229 12184 4263
rect 12218 4229 12252 4263
rect 12286 4229 12320 4263
rect 12354 4229 12388 4263
rect 12621 4229 12655 4263
rect 12689 4229 12723 4263
rect 12973 4229 13007 4263
rect 13041 4229 13075 4263
rect 13311 4229 13345 4263
rect 13379 4229 13413 4263
rect 17719 4304 17753 4338
rect 17787 4304 17821 4338
rect 17855 4304 17889 4338
rect 17923 4304 17957 4338
rect 17991 4304 18025 4338
rect 18059 4304 18093 4338
rect 18127 4304 18161 4338
rect 18195 4304 18229 4338
rect 18263 4304 18297 4338
rect 18331 4304 18365 4338
rect 18399 4304 18433 4338
rect 18467 4304 18501 4338
rect 18535 4304 18569 4338
rect 18603 4304 18637 4338
rect 18671 4304 18705 4338
rect 18739 4304 18773 4338
rect 18807 4304 18841 4338
rect 18875 4304 18909 4338
rect 18943 4304 18977 4338
rect 19011 4304 19045 4338
rect 19079 4304 19113 4338
rect 19147 4304 19181 4338
rect 19215 4304 19249 4338
rect 13171 4121 13205 4155
rect 13239 4121 13273 4155
rect 13307 4121 13341 4155
rect 19599 4126 19633 4160
rect 19667 4126 19701 4160
rect 19735 4126 19769 4160
rect 19803 4126 19837 4160
rect 12352 3948 12386 3982
rect 12352 3880 12386 3914
rect 12352 3812 12386 3846
rect 12352 3744 12386 3778
rect 12352 3676 12386 3710
rect 12352 3608 12386 3642
rect 12352 3540 12386 3574
rect 12352 3472 12386 3506
rect 12352 3404 12386 3438
rect 12352 3336 12386 3370
rect 12352 3268 12386 3302
rect 13038 3966 13072 4000
rect 13038 3894 13072 3928
rect 13038 3822 13072 3856
rect 13038 3750 13072 3784
rect 13038 3678 13072 3712
rect 13038 3606 13072 3640
rect 13038 3534 13072 3568
rect 13038 3462 13072 3496
rect 13038 3390 13072 3424
rect 13038 3318 13072 3352
rect 13038 3246 13072 3280
rect 13737 2996 13771 3030
rect 13805 2996 13839 3030
rect 13944 2996 13978 3030
rect 14012 2996 14046 3030
rect 14080 2996 14114 3030
rect 14148 2996 14182 3030
rect 14216 2996 14250 3030
rect 14284 2996 14318 3030
rect 14352 2996 14386 3030
rect 14420 2996 14454 3030
rect 14488 2996 14522 3030
rect 14556 2996 14590 3030
rect 14624 2996 14658 3030
rect 14692 2996 14726 3030
rect 14760 2996 14794 3030
rect 14828 2996 14862 3030
rect 14896 2996 14930 3030
rect 14964 2996 14998 3030
rect 15032 2996 15066 3030
rect 16833 2996 16867 3030
rect 16901 2996 16935 3030
rect 16969 2996 17003 3030
rect 17037 2996 17071 3030
rect 17105 2996 17139 3030
rect 17173 2996 17207 3030
rect 17241 2996 17275 3030
rect 17309 2996 17343 3030
rect 17377 2996 17411 3030
rect 17445 2996 17479 3030
rect 17513 2996 17547 3030
rect 17581 2996 17615 3030
rect 17649 2996 17683 3030
rect 17717 2996 17751 3030
rect 17785 2996 17819 3030
rect 17853 2996 17887 3030
rect 17921 2996 17955 3030
rect 18273 2996 18307 3030
rect 18341 2996 18375 3030
rect 18409 2996 18443 3030
rect 18477 2996 18511 3030
rect 18545 2996 18579 3030
rect 18613 2996 18647 3030
rect 18681 2996 18715 3030
rect 18749 2996 18783 3030
rect 18897 2996 18931 3030
rect 18965 2996 18999 3030
rect 19033 2996 19067 3030
rect 19101 2996 19135 3030
rect 19169 2996 19203 3030
rect 19237 2996 19271 3030
rect 19305 2996 19339 3030
rect 19373 2996 19407 3030
rect 15389 2946 15423 2980
rect 15457 2946 15491 2980
rect 15525 2946 15559 2980
rect 15593 2946 15627 2980
rect 15661 2946 15695 2980
rect 15729 2946 15763 2980
rect 15797 2946 15831 2980
rect 15865 2946 15899 2980
rect 15933 2946 15967 2980
rect 16001 2946 16035 2980
rect 16069 2946 16103 2980
rect 16137 2946 16171 2980
rect 16205 2946 16239 2980
rect 16273 2946 16307 2980
rect 16341 2946 16375 2980
rect 16409 2946 16443 2980
rect 16477 2946 16511 2980
<< locali >>
rect 7369 6723 7403 6739
rect 7369 6655 7403 6689
rect 7369 6587 7403 6621
rect 7369 6519 7403 6553
rect 7369 6451 7403 6485
rect 7369 6416 7403 6417
rect 7369 6344 7403 6349
rect 7369 6272 7403 6281
rect 7369 6179 7403 6213
rect 7369 6111 7403 6145
rect 7369 6043 7403 6077
rect 7369 5975 7403 6009
rect 7369 5907 7403 5941
rect 7369 5839 7403 5873
rect 7369 5771 7403 5805
rect 7369 5703 7403 5737
rect 7369 5635 7403 5669
rect 7369 5567 7403 5601
rect 7369 5499 7403 5533
rect 7369 5431 7403 5465
rect 7369 5363 7403 5397
rect 7369 5295 7403 5329
rect 7369 5227 7403 5261
rect 7369 5159 7403 5193
rect 7369 5091 7403 5125
rect 7369 5023 7403 5057
rect 7369 4955 7403 4989
rect 7369 4887 7403 4921
rect 7369 4819 7403 4853
rect 7369 4769 7403 4785
rect 7525 6723 7559 6739
rect 7525 6655 7559 6689
rect 7525 6587 7559 6621
rect 7525 6519 7559 6553
rect 7525 6451 7559 6485
rect 7525 6383 7559 6417
rect 7525 6315 7559 6349
rect 7525 6247 7559 6281
rect 7525 6179 7559 6213
rect 7525 6111 7559 6145
rect 7525 6043 7559 6077
rect 7525 5975 7559 6009
rect 7525 5907 7559 5941
rect 7525 5839 7559 5873
rect 7525 5771 7559 5805
rect 7525 5703 7559 5737
rect 7525 5635 7559 5669
rect 7525 5580 7559 5601
rect 7525 5504 7559 5533
rect 7525 5431 7559 5465
rect 7525 5363 7559 5394
rect 7525 5295 7559 5317
rect 7525 5227 7559 5240
rect 7525 5159 7559 5163
rect 7525 5120 7559 5125
rect 7525 5043 7559 5057
rect 7525 4966 7559 4989
rect 7525 4889 7559 4921
rect 7525 4819 7559 4853
rect 7525 4769 7559 4785
rect 7681 6723 7715 6739
rect 7681 6655 7715 6689
rect 7681 6587 7715 6621
rect 7681 6519 7715 6553
rect 7681 6451 7715 6485
rect 7681 6416 7715 6417
rect 7681 6344 7715 6349
rect 7681 6272 7715 6281
rect 7681 6179 7715 6213
rect 7681 6111 7715 6145
rect 7681 6043 7715 6077
rect 7681 5975 7715 6009
rect 7681 5907 7715 5941
rect 7681 5839 7715 5873
rect 7681 5771 7715 5805
rect 7681 5703 7715 5737
rect 7681 5635 7715 5669
rect 7681 5567 7715 5601
rect 7681 5499 7715 5533
rect 7681 5431 7715 5465
rect 7681 5363 7715 5397
rect 7681 5295 7715 5329
rect 7681 5227 7715 5261
rect 7837 6723 7871 6739
rect 7837 6655 7871 6689
rect 7837 6587 7871 6621
rect 7837 6519 7871 6553
rect 7837 6451 7871 6485
rect 7837 6383 7871 6417
rect 7837 6315 7871 6349
rect 7837 6247 7871 6281
rect 7837 6179 7871 6213
rect 7837 6111 7871 6145
rect 7837 6043 7871 6077
rect 7837 5975 7871 6009
rect 7837 5907 7871 5933
rect 7837 5839 7871 5861
rect 7837 5771 7871 5789
rect 7837 5703 7871 5737
rect 7837 5635 7871 5669
rect 7837 5567 7871 5601
rect 7837 5499 7871 5533
rect 7837 5431 7871 5465
rect 7837 5363 7871 5397
rect 7837 5295 7871 5329
rect 7837 5227 7871 5261
rect 7681 5159 7715 5193
rect 7681 5091 7715 5125
rect 7681 5023 7715 5057
rect 7681 4955 7715 4989
rect 7681 4887 7715 4921
rect 7681 4819 7715 4853
rect 7681 4769 7715 4785
rect 7749 5163 7757 5197
rect 7791 5163 7803 5197
rect 7749 5125 7803 5163
rect 7749 5091 7757 5125
rect 7791 5091 7803 5125
rect 7749 4725 7803 5091
rect 7993 6723 8027 6739
rect 7993 6655 8027 6689
rect 7993 6587 8027 6621
rect 7993 6519 8027 6553
rect 7993 6451 8027 6485
rect 7993 6416 8027 6417
rect 7993 6344 8027 6349
rect 7993 6272 8027 6281
rect 7993 6179 8027 6213
rect 7993 6111 8027 6145
rect 7993 6043 8027 6077
rect 7993 5975 8027 6009
rect 7993 5907 8027 5941
rect 7993 5839 8027 5873
rect 7993 5771 8027 5805
rect 7993 5703 8027 5737
rect 7993 5635 8027 5669
rect 12159 5621 12175 5655
rect 12209 5621 12243 5655
rect 12277 5621 12293 5655
rect 7993 5567 8027 5601
rect 7993 5499 8027 5533
rect 7993 5431 8027 5465
rect 7993 5363 8027 5397
rect 7993 5295 8027 5329
rect 7993 5227 8027 5261
rect 7837 5159 7871 5193
rect 7837 5091 7871 5125
rect 7837 5023 7871 5057
rect 7837 4955 7871 4989
rect 7837 4887 7871 4921
rect 7837 4819 7871 4853
rect 7837 4769 7871 4785
rect 7905 5163 7913 5197
rect 7947 5163 7959 5197
rect 7905 5125 7959 5163
rect 7905 5091 7913 5125
rect 7947 5091 7959 5125
rect 7905 4725 7959 5091
rect 7993 5159 8027 5193
rect 7993 5091 8027 5125
rect 7993 5023 8027 5057
rect 7993 4955 8027 4989
rect 7993 4887 8027 4921
rect 7993 4819 8027 4853
rect 12128 5503 12162 5519
rect 12128 5435 12162 5469
rect 12128 5367 12162 5401
rect 12128 5299 12162 5333
rect 12128 5231 12162 5265
rect 12128 5163 12162 5197
rect 12128 5095 12162 5129
rect 12128 5027 12162 5061
rect 12128 4959 12162 4993
rect 12304 5503 12338 5519
rect 12304 5441 12338 5469
rect 12304 5369 12338 5401
rect 12304 5299 12338 5333
rect 12304 5231 12338 5263
rect 12304 5163 12338 5197
rect 12304 5095 12338 5129
rect 12304 5027 12338 5061
rect 12304 4959 12338 4993
rect 12128 4891 12162 4925
rect 11522 4795 11538 4829
rect 11572 4795 11606 4829
rect 11640 4805 11674 4829
rect 11708 4805 11742 4829
rect 11776 4805 11810 4829
rect 11844 4805 11878 4829
rect 11912 4805 11946 4829
rect 11980 4805 12014 4829
rect 11644 4795 11674 4805
rect 11716 4795 11742 4805
rect 11788 4795 11810 4805
rect 11860 4795 11878 4805
rect 11932 4795 11946 4805
rect 12004 4795 12014 4805
rect 12048 4795 12064 4829
rect 12128 4823 12162 4857
rect 7993 4769 8027 4785
rect 11384 4770 11418 4786
rect 11572 4771 11610 4795
rect 11644 4771 11682 4795
rect 11716 4771 11754 4795
rect 11788 4771 11826 4795
rect 11860 4771 11898 4795
rect 11932 4771 11970 4795
rect 12296 4849 12841 4851
rect 12875 4849 12913 4879
rect 12947 4849 12985 4879
rect 13019 4849 13352 4851
rect 12296 4823 12418 4849
rect 12296 4815 12304 4823
rect 7414 4691 7430 4725
rect 7472 4691 7525 4725
rect 7564 4691 7620 4725
rect 7657 4691 7670 4725
rect 7726 4691 7742 4725
rect 7776 4691 7837 4725
rect 7871 4691 7932 4725
rect 7966 4691 7982 4725
rect 11384 4702 11418 4736
rect 12128 4755 12162 4789
rect 12128 4687 12162 4721
rect 11418 4668 11538 4673
rect 11384 4639 11538 4668
rect 11572 4639 11606 4673
rect 11640 4663 11674 4673
rect 11708 4663 11742 4673
rect 11776 4663 11810 4673
rect 11844 4663 11878 4673
rect 11912 4663 11946 4673
rect 11980 4663 12014 4673
rect 11644 4639 11674 4663
rect 11716 4639 11742 4663
rect 11788 4639 11810 4663
rect 11860 4639 11878 4663
rect 11932 4639 11946 4663
rect 12004 4639 12014 4663
rect 12048 4639 12064 4673
rect 11572 4629 11610 4639
rect 11644 4629 11682 4639
rect 11716 4629 11754 4639
rect 11788 4629 11826 4639
rect 11860 4629 11898 4639
rect 11932 4629 11970 4639
rect 12128 4619 12162 4653
rect 12090 4553 12128 4587
rect 12338 4815 12418 4823
rect 12452 4815 12486 4849
rect 12520 4815 12554 4849
rect 12588 4815 12622 4849
rect 12656 4815 12690 4849
rect 12724 4815 12758 4849
rect 12792 4815 12826 4849
rect 12875 4845 12894 4849
rect 12947 4845 12962 4849
rect 13019 4845 13030 4849
rect 12860 4815 12894 4845
rect 12928 4815 12962 4845
rect 12996 4815 13030 4845
rect 13064 4815 13098 4849
rect 13132 4815 13166 4849
rect 13200 4815 13234 4849
rect 13268 4815 13302 4849
rect 13336 4815 13352 4849
rect 12304 4755 12338 4789
rect 13420 4788 13458 4805
rect 13420 4771 13454 4788
rect 12304 4687 12338 4721
rect 13454 4720 13488 4754
rect 12304 4619 12338 4653
rect 12304 4569 12338 4585
rect 12372 4639 12418 4673
rect 12452 4639 12486 4673
rect 12520 4639 12554 4673
rect 12588 4639 12622 4673
rect 12656 4639 12690 4673
rect 12724 4639 12758 4673
rect 12792 4639 12826 4673
rect 12860 4639 12894 4673
rect 12928 4639 12962 4673
rect 12996 4639 13030 4673
rect 13064 4639 13098 4673
rect 13132 4639 13166 4673
rect 13200 4639 13234 4673
rect 13268 4639 13302 4673
rect 13336 4639 13352 4673
rect 13454 4670 13488 4686
rect 7618 4492 7671 4508
rect 7705 4492 7758 4508
rect 7792 4492 7846 4508
rect 7880 4492 7934 4508
rect 11536 4493 11570 4509
rect 7564 4458 7580 4492
rect 7618 4474 7649 4492
rect 7705 4474 7718 4492
rect 7614 4458 7649 4474
rect 7683 4458 7718 4474
rect 7752 4474 7758 4492
rect 7821 4474 7846 4492
rect 7752 4458 7787 4474
rect 7821 4458 7856 4474
rect 7890 4458 7926 4492
rect 7968 4474 7976 4492
rect 7960 4458 7976 4474
rect 11536 4425 11570 4459
rect 11792 4493 11826 4509
rect 11792 4425 11826 4459
rect 7519 4348 7553 4364
rect 7519 4280 7553 4314
rect 7519 4212 7553 4246
rect 7519 4174 7553 4178
rect 7519 4076 7553 4110
rect 7519 4033 7553 4042
rect 7519 3940 7553 3974
rect 7519 3872 7553 3906
rect 7519 3804 7553 3838
rect 7519 3736 7553 3770
rect 7519 3668 7553 3702
rect 7519 3600 7553 3634
rect 7519 3532 7553 3566
rect 7519 3464 7553 3498
rect 7519 3396 7553 3430
rect 7519 3328 7553 3362
rect 7519 3260 7553 3294
rect 7519 3192 7553 3226
rect 7519 3124 7553 3158
rect 7519 3056 7553 3090
rect 7519 3006 7553 3022
rect 7675 4349 7709 4387
rect 7977 4388 8015 4422
rect 7675 4280 7709 4314
rect 7675 4212 7709 4246
rect 7675 4144 7709 4178
rect 7675 4076 7709 4110
rect 7675 4008 7709 4042
rect 7675 3940 7709 3974
rect 7675 3872 7709 3906
rect 7675 3804 7709 3838
rect 7675 3736 7709 3770
rect 7675 3668 7709 3702
rect 7675 3600 7709 3634
rect 7675 3532 7709 3566
rect 7675 3464 7709 3498
rect 7675 3396 7709 3430
rect 7675 3328 7709 3362
rect 7675 3260 7709 3294
rect 7675 3192 7709 3226
rect 7675 3124 7709 3158
rect 7675 3056 7709 3090
rect 7675 3006 7709 3022
rect 7831 4348 7865 4364
rect 7831 4280 7865 4314
rect 7831 4212 7865 4246
rect 7831 4174 7865 4178
rect 7831 4076 7865 4110
rect 7831 4033 7865 4042
rect 7831 3940 7865 3974
rect 7831 3872 7865 3906
rect 7831 3804 7865 3838
rect 7831 3736 7865 3770
rect 7831 3668 7865 3702
rect 7831 3600 7865 3634
rect 7831 3532 7865 3566
rect 7831 3464 7865 3498
rect 7831 3396 7865 3430
rect 7831 3328 7865 3362
rect 7831 3260 7865 3294
rect 7831 3192 7865 3226
rect 7831 3124 7865 3158
rect 7831 3056 7865 3090
rect 7831 3006 7865 3022
rect 7943 4348 8049 4388
rect 7943 4314 7987 4348
rect 8021 4314 8049 4348
rect 7943 4280 8049 4314
rect 11752 4391 11790 4425
rect 11536 4357 11570 4391
rect 11792 4357 11826 4391
rect 11536 4313 11548 4323
rect 11582 4313 11620 4347
rect 12048 4493 12082 4509
rect 12048 4425 12082 4459
rect 12304 4493 12338 4509
rect 12304 4425 12338 4459
rect 12048 4357 12082 4391
rect 12266 4387 12304 4421
rect 11536 4307 11570 4313
rect 11792 4307 11826 4323
rect 12304 4357 12338 4387
rect 12082 4323 12086 4347
rect 12048 4313 12086 4323
rect 12048 4307 12082 4313
rect 12304 4307 12338 4323
rect 7943 4246 7987 4280
rect 8021 4246 8049 4280
rect 12372 4263 12430 4639
rect 12664 4571 12702 4605
rect 12630 4509 12736 4571
rect 12770 4559 12786 4593
rect 12822 4559 12854 4593
rect 12894 4559 12904 4593
rect 12980 4509 13088 4639
rect 13188 4593 13226 4602
rect 13122 4559 13138 4593
rect 13188 4568 13206 4593
rect 13260 4568 13298 4602
rect 13172 4559 13206 4568
rect 13240 4559 13256 4568
rect 12560 4493 12594 4509
rect 12560 4425 12594 4459
rect 12560 4357 12594 4391
rect 7943 4212 8049 4246
rect 7943 4178 7987 4212
rect 8021 4178 8049 4212
rect 7943 4144 8049 4178
rect 11590 4229 11606 4263
rect 11640 4229 11674 4263
rect 11708 4229 11742 4263
rect 11776 4229 11810 4263
rect 11844 4229 11878 4263
rect 11912 4229 11946 4263
rect 11980 4229 12014 4263
rect 12048 4229 12082 4263
rect 12116 4229 12150 4263
rect 12184 4229 12218 4263
rect 12252 4229 12286 4263
rect 12320 4229 12354 4263
rect 12388 4229 12430 4263
rect 11590 4189 12430 4229
rect 11590 4155 11623 4189
rect 11657 4155 11695 4189
rect 11729 4155 11767 4189
rect 11801 4155 11839 4189
rect 11873 4155 11911 4189
rect 11945 4155 11983 4189
rect 12017 4155 12055 4189
rect 12089 4155 12127 4189
rect 12161 4155 12199 4189
rect 12233 4155 12271 4189
rect 12305 4155 12343 4189
rect 12377 4155 12430 4189
rect 12464 4307 12488 4341
rect 12522 4307 12560 4341
rect 12630 4493 12770 4509
rect 12630 4459 12736 4493
rect 12630 4425 12770 4459
rect 12630 4391 12736 4425
rect 12630 4357 12770 4391
rect 12630 4323 12736 4357
rect 12912 4493 12946 4509
rect 12912 4425 12946 4459
rect 12912 4357 12946 4391
rect 12630 4307 12770 4323
rect 12874 4313 12912 4347
rect 12912 4307 12946 4313
rect 12980 4493 13122 4509
rect 12980 4459 13088 4493
rect 12980 4425 13122 4459
rect 12980 4391 13088 4425
rect 12980 4357 13122 4391
rect 12980 4323 13088 4357
rect 13264 4493 13298 4509
rect 13264 4425 13298 4459
rect 13264 4357 13298 4391
rect 12980 4307 13122 4323
rect 13440 4493 13497 4509
rect 13474 4459 13497 4493
rect 13440 4425 13497 4459
rect 13474 4391 13497 4425
rect 13440 4357 13497 4391
rect 13298 4323 13302 4347
rect 13264 4313 13302 4323
rect 13474 4323 13497 4357
rect 13264 4307 13298 4313
rect 13440 4307 13497 4323
rect 7943 4110 7987 4144
rect 8021 4110 8049 4144
rect 7943 4076 8049 4110
rect 7943 4042 7987 4076
rect 8021 4042 8049 4076
rect 12464 4070 12530 4307
rect 12605 4229 12621 4263
rect 12655 4229 12689 4263
rect 12723 4229 12973 4263
rect 13007 4229 13041 4263
rect 13075 4229 13311 4263
rect 13345 4229 13379 4263
rect 13413 4229 13429 4263
rect 13148 4189 13412 4229
rect 13463 4195 13497 4307
rect 17703 4304 17719 4338
rect 17753 4304 17787 4338
rect 17825 4304 17855 4338
rect 17897 4304 17923 4338
rect 17969 4304 17991 4338
rect 18041 4304 18059 4338
rect 18113 4304 18127 4338
rect 18185 4304 18195 4338
rect 18257 4304 18263 4338
rect 18329 4304 18331 4338
rect 18365 4304 18367 4338
rect 18433 4304 18439 4338
rect 18501 4304 18511 4338
rect 18569 4304 18583 4338
rect 18637 4304 18655 4338
rect 18705 4304 18727 4338
rect 18773 4304 18799 4338
rect 18841 4304 18871 4338
rect 18909 4304 18943 4338
rect 18977 4304 19011 4338
rect 19049 4304 19079 4338
rect 19121 4304 19147 4338
rect 19193 4304 19215 4338
rect 13024 4155 13062 4189
rect 13096 4155 13108 4189
rect 7943 4008 8049 4042
rect 12456 4036 12472 4070
rect 12506 4036 12530 4070
rect 12602 4036 12616 4070
rect 7943 3974 7987 4008
rect 8021 3974 8049 4008
rect 12816 4035 12850 4070
rect 7943 3940 8049 3974
rect 7943 3906 7987 3940
rect 8021 3906 8049 3940
rect 7943 3872 8049 3906
rect 7943 3838 7987 3872
rect 8021 3838 8049 3872
rect 7943 3804 8049 3838
rect 7943 3770 7987 3804
rect 8021 3770 8049 3804
rect 7943 3736 8049 3770
rect 7943 3702 7987 3736
rect 8021 3702 8049 3736
rect 7943 3668 8049 3702
rect 7943 3634 7987 3668
rect 8021 3634 8049 3668
rect 7943 3600 8049 3634
rect 7943 3566 7987 3600
rect 8021 3566 8049 3600
rect 7943 3532 8049 3566
rect 7943 3498 7987 3532
rect 8021 3498 8049 3532
rect 7943 3464 8049 3498
rect 7943 3430 7987 3464
rect 8021 3430 8049 3464
rect 7943 3396 8049 3430
rect 12352 3982 12386 3998
rect 12352 3914 12386 3948
rect 12352 3846 12386 3880
rect 12352 3778 12386 3812
rect 12352 3710 12386 3744
rect 12352 3642 12386 3676
rect 12352 3574 12386 3608
rect 12352 3506 12386 3540
rect 12352 3438 12386 3472
rect 12816 3967 12850 4001
rect 12884 4036 12944 4070
rect 12978 4036 12994 4070
rect 12884 4013 12990 4036
rect 12918 3979 12956 4013
rect 13038 4000 13108 4155
rect 13182 4155 13220 4189
rect 13254 4155 13412 4189
rect 13148 4121 13171 4155
rect 13205 4121 13239 4155
rect 13273 4121 13307 4155
rect 13341 4121 13412 4155
rect 13446 4189 13497 4195
rect 17634 4258 17668 4260
rect 17634 4244 17724 4258
rect 17668 4210 17724 4244
rect 13446 4155 13475 4189
rect 13509 4155 13547 4189
rect 13446 4141 13497 4155
rect 13446 4087 13480 4141
rect 12816 3899 12850 3933
rect 12816 3831 12850 3865
rect 13072 3966 13108 4000
rect 13038 3928 13108 3966
rect 13072 3894 13108 3928
rect 13038 3856 13108 3894
rect 12888 3816 12994 3828
rect 12816 3627 12850 3638
rect 12816 3559 12850 3593
rect 12816 3491 12850 3525
rect 7943 3362 7987 3396
rect 8021 3362 8049 3396
rect 12333 3404 12352 3429
rect 12333 3395 12371 3404
rect 12816 3423 12850 3457
rect 7943 3328 8049 3362
rect 7943 3294 7987 3328
rect 8021 3294 8049 3328
rect 7943 3260 8049 3294
rect 7943 3226 7987 3260
rect 8021 3226 8049 3260
rect 12352 3370 12386 3395
rect 12352 3302 12386 3336
rect 12352 3252 12386 3268
rect 12816 3355 12850 3389
rect 12816 3287 12850 3321
rect 7943 3192 8049 3226
rect 12816 3219 12850 3253
rect 7943 3158 7987 3192
rect 8021 3158 8049 3192
rect 12456 3180 12472 3214
rect 12506 3180 12616 3214
rect 12650 3180 12666 3214
rect 7943 3124 8049 3158
rect 7943 3090 7987 3124
rect 8021 3090 8049 3124
rect 7943 3056 8049 3090
rect 12816 3151 12850 3185
rect 12888 3214 12994 3638
rect 13072 3822 13108 3856
rect 13038 3784 13108 3822
rect 13072 3750 13108 3784
rect 13038 3712 13108 3750
rect 13072 3678 13108 3712
rect 13038 3640 13108 3678
rect 13072 3606 13108 3640
rect 13192 4061 13236 4077
rect 13192 4027 13202 4061
rect 13192 3993 13236 4027
rect 13192 3959 13202 3993
rect 13358 4061 13480 4087
rect 13392 4053 13480 4061
rect 13514 4061 13548 4077
rect 13358 3993 13392 4027
rect 13192 3925 13236 3959
rect 13320 3942 13358 3976
rect 13192 3891 13202 3925
rect 13192 3875 13236 3891
rect 13358 3925 13392 3942
rect 13358 3875 13392 3891
rect 13710 4066 13744 4082
rect 13514 3993 13548 4027
rect 13514 3925 13548 3959
rect 13192 3816 13226 3875
rect 13514 3816 13548 3891
rect 13612 4035 13646 4051
rect 13612 3967 13646 4001
rect 13612 3899 13646 3933
rect 13612 3831 13646 3865
rect 13710 3998 13744 4032
rect 13710 3930 13744 3940
rect 13710 3862 13744 3868
rect 13192 3744 13226 3782
rect 13192 3672 13226 3710
rect 13710 3794 13744 3828
rect 13710 3726 13744 3760
rect 13710 3658 13744 3692
rect 13192 3631 13226 3638
rect 13514 3616 13548 3638
rect 13612 3627 13646 3638
rect 13038 3568 13108 3606
rect 13072 3534 13108 3568
rect 13038 3496 13108 3534
rect 13072 3462 13108 3496
rect 13038 3424 13108 3462
rect 13072 3390 13108 3424
rect 13038 3352 13108 3390
rect 13072 3318 13108 3352
rect 13038 3280 13108 3318
rect 13072 3246 13108 3280
rect 13038 3222 13108 3246
rect 13612 3559 13646 3593
rect 13612 3491 13646 3525
rect 13612 3423 13646 3457
rect 13612 3355 13646 3389
rect 13612 3287 13646 3321
rect 12888 3180 12944 3214
rect 12978 3180 12994 3214
rect 13612 3219 13646 3253
rect 12816 3082 12850 3117
rect 13612 3151 13646 3185
rect 13710 3590 13744 3624
rect 13710 3522 13744 3556
rect 13710 3454 13744 3488
rect 13710 3386 13744 3420
rect 13710 3318 13744 3352
rect 13710 3250 13744 3284
rect 13710 3182 13744 3216
rect 13710 3132 13744 3148
rect 13866 4066 13900 4082
rect 13866 3998 13900 4032
rect 13866 3930 13900 3964
rect 13866 3862 13900 3896
rect 13866 3816 13900 3828
rect 13866 3744 13900 3760
rect 13866 3672 13900 3692
rect 13866 3590 13900 3624
rect 13866 3522 13900 3556
rect 13866 3454 13900 3488
rect 13866 3386 13900 3420
rect 13866 3318 13900 3352
rect 13866 3250 13900 3284
rect 13866 3182 13900 3216
rect 13866 3132 13900 3148
rect 14022 4066 14056 4082
rect 14022 3998 14056 4032
rect 14022 3930 14056 3964
rect 14022 3862 14056 3896
rect 14022 3794 14056 3828
rect 14022 3726 14056 3760
rect 14022 3658 14056 3692
rect 14022 3590 14056 3624
rect 14022 3522 14056 3556
rect 14022 3454 14056 3488
rect 14022 3386 14056 3420
rect 14022 3318 14056 3352
rect 14022 3250 14056 3284
rect 14022 3182 14056 3216
rect 13612 3082 13646 3117
rect 14022 3066 14056 3148
rect 14178 4066 14212 4082
rect 14178 3998 14212 4032
rect 14178 3930 14212 3964
rect 14178 3862 14212 3896
rect 14178 3816 14212 3828
rect 14178 3744 14212 3760
rect 14178 3672 14212 3692
rect 14178 3590 14212 3624
rect 14178 3522 14212 3556
rect 14178 3454 14212 3488
rect 14178 3386 14212 3420
rect 14178 3318 14212 3352
rect 14178 3250 14212 3284
rect 14178 3182 14212 3216
rect 14178 3132 14212 3148
rect 14334 4066 14368 4082
rect 14334 3998 14368 4032
rect 14334 3930 14368 3964
rect 14334 3862 14368 3896
rect 14334 3794 14368 3828
rect 14334 3726 14368 3760
rect 14334 3658 14368 3692
rect 14334 3590 14368 3624
rect 14334 3522 14368 3556
rect 14334 3454 14368 3488
rect 14334 3386 14368 3420
rect 14334 3318 14368 3352
rect 14334 3250 14368 3284
rect 14334 3182 14368 3216
rect 14334 3066 14368 3148
rect 14490 4066 14524 4082
rect 14490 3998 14524 4032
rect 14490 3930 14524 3964
rect 14490 3862 14524 3896
rect 14490 3816 14524 3828
rect 14490 3744 14524 3760
rect 14490 3672 14524 3692
rect 14490 3590 14524 3624
rect 14490 3522 14524 3556
rect 14490 3454 14524 3488
rect 14490 3386 14524 3420
rect 14490 3318 14524 3352
rect 14490 3250 14524 3284
rect 14490 3182 14524 3216
rect 14490 3132 14524 3148
rect 14646 4066 14680 4082
rect 14646 3998 14680 4032
rect 14646 3930 14680 3964
rect 14646 3862 14680 3896
rect 14646 3794 14680 3828
rect 14646 3726 14680 3760
rect 14646 3658 14680 3692
rect 14646 3590 14680 3624
rect 14646 3522 14680 3556
rect 14646 3454 14680 3488
rect 14646 3386 14680 3420
rect 14646 3318 14680 3352
rect 14646 3250 14680 3284
rect 14646 3182 14680 3216
rect 14646 3066 14680 3148
rect 14802 4066 14836 4082
rect 14802 3998 14836 4032
rect 14802 3930 14836 3964
rect 14802 3862 14836 3896
rect 14802 3816 14836 3828
rect 14802 3744 14836 3760
rect 14802 3672 14836 3692
rect 14802 3590 14836 3624
rect 14802 3522 14836 3556
rect 14802 3454 14836 3488
rect 14802 3386 14836 3420
rect 14802 3318 14836 3352
rect 14802 3250 14836 3284
rect 14802 3182 14836 3216
rect 14802 3132 14836 3148
rect 14958 4066 14992 4082
rect 14958 3998 14992 4032
rect 14958 3930 14992 3964
rect 14958 3862 14992 3896
rect 14958 3794 14992 3828
rect 15114 4066 15148 4082
rect 15114 3998 15148 4032
rect 15114 3930 15148 3964
rect 15114 3862 15148 3896
rect 15114 3816 15148 3828
rect 15212 4035 15246 4070
rect 16656 4035 16690 4070
rect 15310 4024 15344 4032
rect 15212 3967 15246 4001
rect 15212 3899 15246 3933
rect 15212 3831 15246 3865
rect 14958 3726 14992 3760
rect 14958 3658 14992 3692
rect 14958 3590 14992 3624
rect 14958 3522 14992 3556
rect 14958 3454 14992 3488
rect 14958 3386 14992 3420
rect 14958 3318 14992 3352
rect 14958 3250 14992 3284
rect 14958 3182 14992 3216
rect 14958 3066 14992 3148
rect 15114 3590 15148 3624
rect 15114 3522 15148 3556
rect 15114 3454 15148 3488
rect 15114 3386 15148 3420
rect 15114 3318 15148 3352
rect 15114 3250 15148 3284
rect 15114 3182 15148 3216
rect 15114 3132 15148 3148
rect 15212 3627 15246 3638
rect 15212 3559 15246 3593
rect 15212 3491 15246 3525
rect 15212 3423 15246 3457
rect 15212 3355 15246 3389
rect 15212 3287 15246 3321
rect 15212 3219 15246 3253
rect 15212 3151 15246 3185
rect 15212 3082 15246 3117
rect 15305 4016 15344 4024
rect 15305 3982 15310 4016
rect 15305 3948 15344 3982
rect 15305 3914 15310 3948
rect 15305 3880 15344 3914
rect 15466 4016 15500 4032
rect 15466 3948 15500 3982
rect 15466 3896 15500 3914
rect 15622 4016 15656 4032
rect 15622 3948 15656 3982
rect 15305 3846 15310 3880
rect 15466 3880 15504 3896
rect 15305 3812 15344 3846
rect 15305 3778 15310 3812
rect 15305 3744 15344 3778
rect 15305 3710 15310 3744
rect 15305 3676 15344 3710
rect 15305 3642 15310 3676
rect 15305 3608 15344 3642
rect 15305 3574 15310 3608
rect 15500 3862 15504 3880
rect 15622 3880 15656 3914
rect 15778 4016 15812 4032
rect 15778 3948 15812 3982
rect 15778 3896 15812 3914
rect 15934 4016 15968 4032
rect 15934 3948 15968 3982
rect 15466 3812 15500 3846
rect 15466 3744 15500 3778
rect 15466 3676 15500 3710
rect 15466 3608 15500 3642
rect 15305 3558 15311 3574
rect 15345 3558 15383 3592
rect 15778 3880 15816 3896
rect 15622 3812 15656 3846
rect 15622 3744 15656 3778
rect 15622 3676 15656 3710
rect 15622 3608 15656 3642
rect 15812 3862 15816 3880
rect 15934 3880 15968 3914
rect 16090 4016 16124 4032
rect 16090 3948 16124 3982
rect 16090 3896 16124 3914
rect 16246 4016 16280 4032
rect 16246 3948 16280 3982
rect 15778 3812 15812 3846
rect 15778 3744 15812 3778
rect 15778 3676 15812 3710
rect 15778 3608 15812 3642
rect 15305 3540 15344 3558
rect 15305 3506 15310 3540
rect 15305 3472 15344 3506
rect 15305 3438 15310 3472
rect 15305 3404 15344 3438
rect 15305 3370 15310 3404
rect 15305 3336 15344 3370
rect 15305 3302 15310 3336
rect 15305 3268 15344 3302
rect 15305 3234 15310 3268
rect 15305 3200 15344 3234
rect 15305 3166 15310 3200
rect 15305 3132 15344 3166
rect 15305 3098 15310 3132
rect 15305 3082 15344 3098
rect 15466 3540 15500 3574
rect 15656 3574 15661 3592
rect 15623 3558 15661 3574
rect 16090 3880 16128 3896
rect 15934 3812 15968 3846
rect 15934 3744 15968 3778
rect 15934 3676 15968 3710
rect 15934 3608 15968 3642
rect 16124 3862 16128 3880
rect 16246 3880 16280 3914
rect 16402 4016 16436 4032
rect 16402 3948 16436 3982
rect 16402 3896 16436 3914
rect 16558 4016 16592 4032
rect 16558 3948 16592 3982
rect 16090 3812 16124 3846
rect 16090 3744 16124 3778
rect 16090 3676 16124 3710
rect 16090 3608 16124 3642
rect 15466 3472 15500 3506
rect 15466 3404 15500 3438
rect 15466 3336 15500 3370
rect 15466 3268 15500 3302
rect 15466 3200 15500 3234
rect 15466 3132 15500 3166
rect 7943 3022 7987 3056
rect 8021 3022 8049 3056
rect 7943 3006 8049 3022
rect 13721 3030 13855 3066
rect 13721 2996 13737 3030
rect 13771 2996 13805 3030
rect 13839 2996 13855 3030
rect 13928 3032 13951 3066
rect 13985 3032 14023 3066
rect 14057 3032 14095 3066
rect 14129 3032 14167 3066
rect 14201 3032 14239 3066
rect 14273 3032 14311 3066
rect 14345 3032 14383 3066
rect 14417 3032 14455 3066
rect 14489 3032 14527 3066
rect 14561 3032 14599 3066
rect 14633 3032 14671 3066
rect 14705 3032 14743 3066
rect 14777 3032 14815 3066
rect 14849 3032 14887 3066
rect 14921 3032 14959 3066
rect 14993 3032 15031 3066
rect 15065 3032 15082 3066
rect 15305 3032 15339 3082
rect 13928 3030 15339 3032
rect 13928 2996 13944 3030
rect 13978 2996 14012 3030
rect 14046 2996 14080 3030
rect 14114 2996 14148 3030
rect 14182 2996 14216 3030
rect 14250 2996 14284 3030
rect 14318 2996 14352 3030
rect 14386 2996 14420 3030
rect 14454 2996 14488 3030
rect 14522 2996 14556 3030
rect 14590 2996 14624 3030
rect 14658 2996 14692 3030
rect 14726 2996 14760 3030
rect 14794 2996 14828 3030
rect 14862 2996 14896 3030
rect 14930 2996 14964 3030
rect 14998 2996 15032 3030
rect 15066 2996 15339 3030
rect 15466 3016 15500 3098
rect 15622 3540 15656 3558
rect 15622 3472 15656 3506
rect 15622 3404 15656 3438
rect 15622 3336 15656 3370
rect 15622 3268 15656 3302
rect 15622 3200 15656 3234
rect 15622 3132 15656 3166
rect 15622 3082 15656 3098
rect 15778 3540 15812 3574
rect 15968 3574 15973 3592
rect 15935 3558 15973 3574
rect 16402 3880 16440 3896
rect 16246 3812 16280 3846
rect 16246 3744 16280 3778
rect 16246 3676 16280 3710
rect 16246 3608 16280 3642
rect 16436 3862 16440 3880
rect 16558 3880 16592 3914
rect 16402 3812 16436 3846
rect 16402 3744 16436 3778
rect 16402 3676 16436 3710
rect 16402 3608 16436 3642
rect 15778 3472 15812 3506
rect 15778 3404 15812 3438
rect 15778 3336 15812 3370
rect 15778 3268 15812 3302
rect 15778 3200 15812 3234
rect 15778 3132 15812 3166
rect 15778 3016 15812 3098
rect 15934 3540 15968 3558
rect 15934 3472 15968 3506
rect 15934 3404 15968 3438
rect 15934 3336 15968 3370
rect 15934 3268 15968 3302
rect 15934 3200 15968 3234
rect 15934 3132 15968 3166
rect 15934 3082 15968 3098
rect 16090 3540 16124 3574
rect 16280 3574 16285 3592
rect 16247 3558 16285 3574
rect 16558 3812 16592 3846
rect 16558 3744 16592 3778
rect 16558 3676 16592 3710
rect 16558 3608 16592 3642
rect 16656 3967 16690 4001
rect 16656 3899 16690 3933
rect 16656 3831 16690 3865
rect 16754 4066 16788 4082
rect 16754 3998 16788 4032
rect 16754 3930 16788 3964
rect 16754 3862 16788 3896
rect 16754 3816 16788 3828
rect 16910 4066 16944 4082
rect 16910 3998 16944 4032
rect 16910 3930 16944 3964
rect 16910 3862 16944 3896
rect 16656 3763 16657 3797
rect 16656 3695 16657 3729
rect 16656 3638 16657 3661
rect 16910 3794 16944 3828
rect 16910 3726 16944 3760
rect 16910 3658 16944 3692
rect 16656 3627 16690 3638
rect 16090 3472 16124 3506
rect 16090 3404 16124 3438
rect 16090 3336 16124 3370
rect 16090 3268 16124 3302
rect 16090 3200 16124 3234
rect 16090 3132 16124 3166
rect 16090 3016 16124 3098
rect 16246 3540 16280 3558
rect 16246 3472 16280 3506
rect 16246 3404 16280 3438
rect 16246 3336 16280 3370
rect 16246 3268 16280 3302
rect 16246 3200 16280 3234
rect 16246 3132 16280 3166
rect 16246 3082 16280 3098
rect 16402 3540 16436 3574
rect 16521 3574 16558 3592
rect 16521 3558 16559 3574
rect 16656 3559 16690 3593
rect 16402 3472 16436 3506
rect 16402 3404 16436 3438
rect 16402 3336 16436 3370
rect 16402 3268 16436 3302
rect 16402 3200 16436 3234
rect 16402 3132 16436 3166
rect 16402 3016 16436 3098
rect 16558 3540 16592 3558
rect 16558 3472 16592 3506
rect 16558 3404 16592 3438
rect 16558 3336 16592 3370
rect 16558 3268 16592 3302
rect 16558 3200 16592 3234
rect 16558 3132 16592 3166
rect 16558 3082 16592 3098
rect 16656 3491 16690 3525
rect 16656 3423 16690 3457
rect 16656 3355 16690 3389
rect 16656 3287 16690 3321
rect 16656 3219 16690 3253
rect 16656 3151 16690 3185
rect 16754 3590 16788 3624
rect 16910 3592 16944 3624
rect 17066 4066 17100 4082
rect 17066 3998 17100 4032
rect 17066 3930 17100 3964
rect 17066 3862 17100 3896
rect 17066 3816 17100 3828
rect 17066 3744 17100 3760
rect 17066 3672 17100 3692
rect 16911 3590 16949 3592
rect 16944 3558 16949 3590
rect 17066 3590 17100 3624
rect 17222 4066 17256 4082
rect 17222 3998 17256 4032
rect 17222 3930 17256 3964
rect 17222 3862 17256 3896
rect 17222 3794 17256 3828
rect 17222 3726 17256 3760
rect 17222 3658 17256 3692
rect 17222 3592 17256 3624
rect 17378 4066 17412 4082
rect 17378 3998 17412 4032
rect 17378 3930 17412 3964
rect 17378 3862 17412 3896
rect 17378 3816 17412 3828
rect 17378 3744 17412 3760
rect 17378 3672 17412 3692
rect 16754 3522 16788 3556
rect 16754 3454 16788 3488
rect 16754 3386 16788 3420
rect 16754 3318 16788 3352
rect 16754 3250 16788 3284
rect 16754 3182 16788 3216
rect 16754 3132 16788 3148
rect 16910 3522 16944 3556
rect 16910 3454 16944 3488
rect 16910 3386 16944 3420
rect 16910 3318 16944 3352
rect 16910 3250 16944 3284
rect 16910 3182 16944 3216
rect 16910 3132 16944 3148
rect 17222 3590 17260 3592
rect 17066 3522 17100 3556
rect 17066 3454 17100 3488
rect 17066 3386 17100 3420
rect 17066 3318 17100 3352
rect 17066 3250 17100 3284
rect 17066 3182 17100 3216
rect 17066 3132 17100 3148
rect 17256 3558 17260 3590
rect 17378 3590 17412 3624
rect 17534 4066 17568 4082
rect 17534 3998 17568 4032
rect 17534 3930 17568 3964
rect 17534 3862 17568 3896
rect 17534 3794 17568 3828
rect 17534 3726 17568 3760
rect 17534 3658 17568 3692
rect 17534 3592 17568 3624
rect 17634 4066 17724 4210
rect 19290 4244 19324 4260
rect 17634 4032 17690 4066
rect 17634 3998 17724 4032
rect 17634 3964 17690 3998
rect 17634 3930 17724 3964
rect 17634 3896 17690 3930
rect 17634 3862 17724 3896
rect 17634 3828 17690 3862
rect 17634 3816 17724 3828
rect 17846 4066 17880 4082
rect 17846 3998 17880 4032
rect 17846 3930 17880 3964
rect 17846 3862 17880 3896
rect 17634 3638 17640 3816
rect 17846 3794 17880 3828
rect 18002 4066 18036 4082
rect 18002 3998 18036 4032
rect 18002 3930 18036 3964
rect 18002 3862 18036 3896
rect 18002 3816 18036 3828
rect 18100 4035 18134 4070
rect 18100 3967 18134 4001
rect 18100 3899 18134 3933
rect 18100 3831 18134 3865
rect 17846 3726 17880 3760
rect 17846 3658 17880 3692
rect 17634 3624 17690 3638
rect 17222 3522 17256 3556
rect 17222 3454 17256 3488
rect 17222 3386 17256 3420
rect 17222 3318 17256 3352
rect 17222 3250 17256 3284
rect 17222 3182 17256 3216
rect 17222 3132 17256 3148
rect 17528 3590 17566 3592
rect 17528 3558 17534 3590
rect 17634 3590 17724 3624
rect 17846 3592 17880 3624
rect 17378 3522 17412 3556
rect 17378 3454 17412 3488
rect 17378 3386 17412 3420
rect 17378 3318 17412 3352
rect 17378 3250 17412 3284
rect 17378 3182 17412 3216
rect 17378 3132 17412 3148
rect 17534 3522 17568 3556
rect 17534 3454 17568 3488
rect 17534 3386 17568 3420
rect 17534 3318 17568 3352
rect 17534 3250 17568 3284
rect 17534 3182 17568 3216
rect 17534 3132 17568 3148
rect 17634 3556 17690 3590
rect 17846 3590 17884 3592
rect 17634 3522 17724 3556
rect 17634 3488 17690 3522
rect 17634 3454 17724 3488
rect 17634 3420 17690 3454
rect 17634 3386 17724 3420
rect 17634 3352 17690 3386
rect 17634 3318 17724 3352
rect 17634 3284 17690 3318
rect 17634 3250 17724 3284
rect 17634 3216 17690 3250
rect 17634 3182 17724 3216
rect 17634 3148 17690 3182
rect 17634 3132 17724 3148
rect 17880 3558 17884 3590
rect 18002 3590 18036 3624
rect 17846 3522 17880 3556
rect 17846 3454 17880 3488
rect 17846 3386 17880 3420
rect 17846 3318 17880 3352
rect 17846 3250 17880 3284
rect 17846 3182 17880 3216
rect 17846 3132 17880 3148
rect 18002 3522 18036 3556
rect 18002 3454 18036 3488
rect 18002 3386 18036 3420
rect 18002 3318 18036 3352
rect 18002 3250 18036 3284
rect 18002 3182 18036 3216
rect 18002 3132 18036 3148
rect 18100 3627 18134 3638
rect 18100 3559 18134 3593
rect 18100 3491 18134 3525
rect 18100 3423 18134 3457
rect 18100 3355 18134 3389
rect 18100 3287 18134 3321
rect 18100 3219 18134 3253
rect 18100 3151 18134 3185
rect 16656 3082 16690 3117
rect 18198 4066 18232 4082
rect 18198 3998 18232 4032
rect 18198 3930 18232 3964
rect 18198 3862 18232 3896
rect 18198 3794 18232 3828
rect 18198 3726 18232 3760
rect 18198 3658 18232 3692
rect 18198 3592 18232 3624
rect 18354 4066 18388 4082
rect 18354 3998 18388 4032
rect 18354 3930 18388 3964
rect 18354 3862 18388 3896
rect 18354 3794 18388 3828
rect 18354 3726 18388 3760
rect 18354 3658 18388 3692
rect 18232 3558 18270 3592
rect 18354 3590 18388 3624
rect 18510 4066 18544 4082
rect 18510 3998 18544 4032
rect 18510 3930 18544 3964
rect 18510 3862 18544 3896
rect 18510 3794 18544 3828
rect 18510 3726 18544 3760
rect 18510 3658 18544 3692
rect 18510 3592 18544 3624
rect 18666 4066 18700 4082
rect 18666 3998 18700 4032
rect 18666 3930 18700 3964
rect 18666 3862 18700 3896
rect 18666 3794 18700 3828
rect 18666 3726 18700 3760
rect 18666 3658 18700 3692
rect 18198 3522 18232 3556
rect 18198 3454 18232 3488
rect 18510 3590 18548 3592
rect 18354 3522 18388 3556
rect 18354 3456 18388 3488
rect 18544 3558 18548 3590
rect 18666 3590 18700 3624
rect 18822 4066 18856 4082
rect 18822 4024 18856 4032
rect 18978 4066 19012 4082
rect 18822 3998 18867 4024
rect 18856 3964 18867 3998
rect 18822 3930 18867 3964
rect 18856 3896 18867 3930
rect 18822 3862 18867 3896
rect 18856 3828 18867 3862
rect 18822 3794 18867 3828
rect 18856 3760 18867 3794
rect 18822 3726 18867 3760
rect 18856 3692 18867 3726
rect 18822 3658 18867 3692
rect 18856 3624 18867 3658
rect 18822 3592 18867 3624
rect 18978 3998 19012 4032
rect 18978 3930 19012 3964
rect 18978 3862 19012 3896
rect 18978 3794 19012 3828
rect 18978 3726 19012 3760
rect 18978 3658 19012 3692
rect 18510 3522 18544 3556
rect 18354 3454 18392 3456
rect 18198 3386 18232 3420
rect 18198 3318 18232 3352
rect 18198 3250 18232 3284
rect 18198 3182 18232 3216
rect 18198 3132 18232 3148
rect 18388 3422 18392 3454
rect 18510 3454 18544 3488
rect 18822 3590 18860 3592
rect 18666 3522 18700 3556
rect 18666 3456 18700 3488
rect 18856 3558 18860 3590
rect 18978 3590 19012 3624
rect 19134 4066 19168 4082
rect 19134 3998 19168 4032
rect 19134 3930 19168 3964
rect 19134 3862 19168 3896
rect 19134 3794 19168 3828
rect 19134 3726 19168 3760
rect 19134 3658 19168 3692
rect 19134 3592 19168 3624
rect 19290 4066 19324 4210
rect 19583 4155 19591 4189
rect 19625 4160 19663 4189
rect 19697 4160 19735 4189
rect 19769 4160 19807 4189
rect 19633 4155 19663 4160
rect 19583 4126 19599 4155
rect 19633 4126 19667 4155
rect 19701 4126 19735 4160
rect 19769 4126 19803 4160
rect 19841 4155 19853 4189
rect 19837 4126 19853 4155
rect 19290 3998 19324 4032
rect 19290 3930 19324 3964
rect 19290 3862 19324 3896
rect 19290 3794 19324 3828
rect 19290 3726 19324 3760
rect 19290 3658 19324 3692
rect 18856 3556 18867 3558
rect 18822 3522 18867 3556
rect 18856 3488 18867 3522
rect 18354 3386 18388 3420
rect 18354 3318 18388 3352
rect 18354 3250 18388 3284
rect 18354 3182 18388 3216
rect 18100 3082 18134 3117
rect 16817 3026 16830 3060
rect 16864 3030 16902 3060
rect 16936 3030 16974 3060
rect 17008 3030 17046 3060
rect 17080 3030 17118 3060
rect 17152 3030 17190 3060
rect 17224 3030 17262 3060
rect 17296 3030 17334 3060
rect 17368 3030 17406 3060
rect 17440 3030 17478 3060
rect 17512 3030 17550 3060
rect 17584 3030 17622 3060
rect 17656 3030 17694 3060
rect 17728 3030 17766 3060
rect 17800 3030 17838 3060
rect 17872 3030 17910 3060
rect 17944 3030 17971 3060
rect 18354 3030 18388 3148
rect 18665 3454 18703 3456
rect 18665 3422 18666 3454
rect 18510 3386 18544 3420
rect 18510 3318 18544 3352
rect 18510 3250 18544 3284
rect 18510 3182 18544 3216
rect 18510 3132 18544 3148
rect 18700 3422 18703 3454
rect 18822 3454 18867 3488
rect 18666 3386 18700 3420
rect 18666 3318 18700 3352
rect 18666 3250 18700 3284
rect 18666 3182 18700 3216
rect 18666 3030 18700 3148
rect 18856 3420 18867 3454
rect 18822 3386 18867 3420
rect 18856 3352 18867 3386
rect 19134 3590 19172 3592
rect 18978 3522 19012 3556
rect 18978 3454 19012 3488
rect 18978 3386 19012 3420
rect 18822 3318 18867 3352
rect 19168 3558 19172 3590
rect 19290 3590 19324 3624
rect 19446 4066 19480 4082
rect 19446 3998 19480 4032
rect 19446 3930 19480 3964
rect 19446 3862 19480 3896
rect 19446 3794 19480 3828
rect 19446 3726 19480 3760
rect 19446 3658 19480 3692
rect 19446 3592 19480 3624
rect 19134 3522 19168 3556
rect 19134 3454 19168 3488
rect 19134 3386 19168 3420
rect 19012 3352 19016 3370
rect 18978 3336 19016 3352
rect 19408 3558 19446 3592
rect 19290 3522 19324 3556
rect 19290 3454 19324 3488
rect 19290 3386 19324 3420
rect 18856 3284 18867 3318
rect 18822 3250 18867 3284
rect 18856 3216 18867 3250
rect 18822 3182 18867 3216
rect 18856 3148 18867 3182
rect 18822 3132 18867 3148
rect 18978 3318 19012 3336
rect 18978 3250 19012 3284
rect 18978 3182 19012 3216
rect 18978 3132 19012 3148
rect 19134 3318 19168 3352
rect 19289 3352 19290 3370
rect 19446 3522 19480 3556
rect 19446 3454 19480 3488
rect 19446 3386 19480 3420
rect 19324 3352 19327 3370
rect 19289 3336 19327 3352
rect 19134 3250 19168 3284
rect 19134 3182 19168 3216
rect 18833 3030 18867 3132
rect 19134 3030 19168 3148
rect 19290 3318 19324 3336
rect 19290 3250 19324 3284
rect 19290 3182 19324 3216
rect 19290 3132 19324 3148
rect 19446 3318 19480 3352
rect 19446 3250 19480 3284
rect 19446 3182 19480 3216
rect 19446 3030 19480 3148
rect 19556 4066 19590 4082
rect 19556 3998 19590 4032
rect 19556 3930 19590 3964
rect 19556 3862 19590 3896
rect 19556 3794 19590 3828
rect 19556 3726 19590 3760
rect 19556 3658 19590 3692
rect 19556 3590 19590 3624
rect 19556 3522 19590 3556
rect 19556 3454 19590 3488
rect 19556 3386 19590 3420
rect 19712 4066 19746 4082
rect 19712 3998 19746 4032
rect 19712 3930 19746 3964
rect 19868 4066 19902 4082
rect 19868 3998 19902 4032
rect 19868 3930 19902 3964
rect 19712 3862 19746 3896
rect 19830 3862 19868 3896
rect 19712 3816 19746 3828
rect 19712 3744 19746 3760
rect 19712 3672 19746 3692
rect 19712 3590 19746 3624
rect 19712 3522 19746 3556
rect 19712 3454 19746 3488
rect 19712 3386 19746 3420
rect 19590 3336 19628 3370
rect 19556 3318 19590 3336
rect 19556 3250 19590 3284
rect 19556 3182 19590 3216
rect 19556 3132 19590 3148
rect 19712 3318 19746 3352
rect 19712 3250 19746 3284
rect 19712 3182 19746 3216
rect 19712 3132 19746 3148
rect 19868 3794 19902 3828
rect 19868 3726 19902 3760
rect 19868 3658 19902 3692
rect 19868 3590 19902 3624
rect 19868 3522 19902 3556
rect 19868 3454 19902 3488
rect 19868 3386 19902 3420
rect 19868 3318 19902 3352
rect 19868 3250 19902 3284
rect 19868 3182 19902 3216
rect 19868 3132 19902 3148
rect 19966 3287 20071 3344
rect 20000 3253 20071 3287
rect 19966 3219 20071 3253
rect 20000 3185 20071 3219
rect 19966 3151 20071 3185
rect 15373 2982 16527 3016
rect 16817 2996 16833 3026
rect 16867 2996 16901 3030
rect 16936 3026 16969 3030
rect 17008 3026 17037 3030
rect 17080 3026 17105 3030
rect 17152 3026 17173 3030
rect 17224 3026 17241 3030
rect 17296 3026 17309 3030
rect 17368 3026 17377 3030
rect 17440 3026 17445 3030
rect 17512 3026 17513 3030
rect 16935 2996 16969 3026
rect 17003 2996 17037 3026
rect 17071 2996 17105 3026
rect 17139 2996 17173 3026
rect 17207 2996 17241 3026
rect 17275 2996 17309 3026
rect 17343 2996 17377 3026
rect 17411 2996 17445 3026
rect 17479 2996 17513 3026
rect 17547 3026 17550 3030
rect 17615 3026 17622 3030
rect 17683 3026 17694 3030
rect 17751 3026 17766 3030
rect 17819 3026 17838 3030
rect 17887 3026 17910 3030
rect 17547 2996 17581 3026
rect 17615 2996 17649 3026
rect 17683 2996 17717 3026
rect 17751 2996 17785 3026
rect 17819 2996 17853 3026
rect 17887 2996 17921 3026
rect 17955 2996 17971 3030
rect 18257 2996 18273 3030
rect 18307 2996 18341 3030
rect 18375 2996 18409 3030
rect 18443 2996 18477 3030
rect 18511 2996 18545 3030
rect 18579 2996 18613 3030
rect 18647 2996 18681 3030
rect 18715 2996 18749 3030
rect 18783 2996 18799 3030
rect 18833 2996 18897 3030
rect 18931 2996 18965 3030
rect 18999 2996 19033 3030
rect 19067 2996 19101 3030
rect 19135 2996 19169 3030
rect 19203 2996 19237 3030
rect 19271 2996 19305 3030
rect 19339 2996 19373 3030
rect 19407 2996 19480 3030
rect 20000 3117 20071 3151
rect 19966 3083 20071 3117
rect 20000 3049 20071 3083
rect 19966 3015 20071 3049
rect 20000 3012 20071 3015
rect 15373 2980 15401 2982
rect 15435 2980 15473 2982
rect 15507 2980 15545 2982
rect 15579 2980 15617 2982
rect 15651 2980 15689 2982
rect 15723 2980 15761 2982
rect 15795 2980 15833 2982
rect 15867 2980 15905 2982
rect 15939 2980 15977 2982
rect 16011 2980 16049 2982
rect 16083 2980 16121 2982
rect 16155 2980 16193 2982
rect 16227 2980 16265 2982
rect 16299 2980 16337 2982
rect 16371 2980 16409 2982
rect 16443 2980 16481 2982
rect 15373 2946 15389 2980
rect 15435 2948 15457 2980
rect 15507 2948 15525 2980
rect 15579 2948 15593 2980
rect 15651 2948 15661 2980
rect 15723 2948 15729 2980
rect 15795 2948 15797 2980
rect 15423 2946 15457 2948
rect 15491 2946 15525 2948
rect 15559 2946 15593 2948
rect 15627 2946 15661 2948
rect 15695 2946 15729 2948
rect 15763 2946 15797 2948
rect 15831 2948 15833 2980
rect 15899 2948 15905 2980
rect 15967 2948 15977 2980
rect 16035 2948 16049 2980
rect 16103 2948 16121 2980
rect 16171 2948 16193 2980
rect 16239 2948 16265 2980
rect 16307 2948 16337 2980
rect 15831 2946 15865 2948
rect 15899 2946 15933 2948
rect 15967 2946 16001 2948
rect 16035 2946 16069 2948
rect 16103 2946 16137 2948
rect 16171 2946 16205 2948
rect 16239 2946 16273 2948
rect 16307 2946 16341 2948
rect 16375 2946 16409 2980
rect 16443 2946 16477 2980
rect 16515 2948 16527 2982
rect 16511 2946 16527 2948
rect 19966 2882 20071 3012
<< viali >>
rect 7369 6383 7403 6416
rect 7369 6382 7403 6383
rect 7369 6315 7403 6344
rect 7369 6310 7403 6315
rect 7369 6247 7403 6272
rect 7369 6238 7403 6247
rect 7525 5567 7559 5580
rect 7525 5546 7559 5567
rect 7525 5499 7559 5504
rect 7525 5470 7559 5499
rect 7525 5397 7559 5428
rect 7525 5394 7559 5397
rect 7525 5329 7559 5351
rect 7525 5317 7559 5329
rect 7525 5261 7559 5274
rect 7525 5240 7559 5261
rect 7525 5193 7559 5197
rect 7525 5163 7559 5193
rect 7525 5091 7559 5120
rect 7525 5086 7559 5091
rect 7525 5023 7559 5043
rect 7525 5009 7559 5023
rect 7525 4955 7559 4966
rect 7525 4932 7559 4955
rect 7525 4887 7559 4889
rect 7525 4855 7559 4887
rect 7681 6383 7715 6416
rect 7681 6382 7715 6383
rect 7681 6315 7715 6344
rect 7681 6310 7715 6315
rect 7681 6247 7715 6272
rect 7681 6238 7715 6247
rect 7837 5941 7871 5967
rect 7837 5933 7871 5941
rect 7837 5873 7871 5895
rect 7837 5861 7871 5873
rect 7837 5805 7871 5823
rect 7837 5789 7871 5805
rect 7757 5163 7791 5197
rect 7757 5091 7791 5125
rect 7993 6383 8027 6416
rect 7993 6382 8027 6383
rect 7993 6315 8027 6344
rect 7993 6310 8027 6315
rect 7993 6247 8027 6272
rect 7993 6238 8027 6247
rect 7913 5163 7947 5197
rect 7913 5091 7947 5125
rect 12304 5435 12338 5441
rect 12304 5407 12338 5435
rect 12304 5367 12338 5369
rect 12304 5335 12338 5367
rect 12304 5265 12338 5297
rect 12304 5263 12338 5265
rect 11538 4795 11572 4805
rect 11610 4795 11640 4805
rect 11640 4795 11644 4805
rect 11682 4795 11708 4805
rect 11708 4795 11716 4805
rect 11754 4795 11776 4805
rect 11776 4795 11788 4805
rect 11826 4795 11844 4805
rect 11844 4795 11860 4805
rect 11898 4795 11912 4805
rect 11912 4795 11932 4805
rect 11970 4795 11980 4805
rect 11980 4795 12004 4805
rect 11538 4771 11572 4795
rect 11610 4771 11644 4795
rect 11682 4771 11716 4795
rect 11754 4771 11788 4795
rect 11826 4771 11860 4795
rect 11898 4771 11932 4795
rect 11970 4771 12004 4795
rect 12296 4925 12304 4957
rect 12304 4925 12338 4957
rect 12338 4925 12402 4957
rect 12296 4891 12402 4925
rect 12296 4857 12304 4891
rect 12304 4857 12338 4891
rect 12338 4857 12402 4891
rect 12296 4851 12402 4857
rect 12841 4849 12875 4879
rect 12913 4849 12947 4879
rect 12985 4849 13019 4879
rect 7438 4691 7464 4725
rect 7464 4691 7472 4725
rect 7530 4691 7559 4725
rect 7559 4691 7564 4725
rect 7623 4691 7654 4725
rect 7654 4691 7657 4725
rect 11538 4639 11572 4663
rect 11610 4639 11640 4663
rect 11640 4639 11644 4663
rect 11682 4639 11708 4663
rect 11708 4639 11716 4663
rect 11754 4639 11776 4663
rect 11776 4639 11788 4663
rect 11826 4639 11844 4663
rect 11844 4639 11860 4663
rect 11898 4639 11912 4663
rect 11912 4639 11932 4663
rect 11970 4639 11980 4663
rect 11980 4639 12004 4663
rect 11538 4629 11572 4639
rect 11610 4629 11644 4639
rect 11682 4629 11716 4639
rect 11754 4629 11788 4639
rect 11826 4629 11860 4639
rect 11898 4629 11932 4639
rect 11970 4629 12004 4639
rect 12056 4553 12090 4587
rect 12128 4585 12162 4587
rect 12128 4553 12162 4585
rect 12841 4845 12860 4849
rect 12860 4845 12875 4849
rect 12913 4845 12928 4849
rect 12928 4845 12947 4849
rect 12985 4845 12996 4849
rect 12996 4845 13019 4849
rect 13386 4771 13420 4805
rect 13458 4788 13492 4805
rect 13458 4771 13488 4788
rect 13488 4771 13492 4788
rect 7584 4492 7618 4508
rect 7671 4492 7705 4508
rect 7758 4492 7792 4508
rect 7846 4492 7880 4508
rect 7934 4492 7968 4508
rect 7584 4474 7614 4492
rect 7614 4474 7618 4492
rect 7671 4474 7683 4492
rect 7683 4474 7705 4492
rect 7758 4474 7787 4492
rect 7787 4474 7792 4492
rect 7846 4474 7856 4492
rect 7856 4474 7880 4492
rect 7934 4474 7960 4492
rect 7960 4474 7968 4492
rect 7675 4387 7709 4421
rect 7519 4144 7553 4174
rect 7519 4140 7553 4144
rect 7519 4008 7553 4033
rect 7519 3999 7553 4008
rect 7943 4388 7977 4422
rect 8015 4388 8049 4422
rect 7675 4348 7709 4349
rect 7675 4315 7709 4348
rect 7831 4144 7865 4174
rect 7831 4140 7865 4144
rect 7831 4008 7865 4033
rect 7831 3999 7865 4008
rect 11718 4391 11752 4425
rect 11790 4391 11792 4425
rect 11792 4391 11824 4425
rect 11548 4323 11570 4347
rect 11570 4323 11582 4347
rect 11548 4313 11582 4323
rect 11620 4313 11654 4347
rect 12232 4387 12266 4421
rect 12304 4391 12338 4421
rect 12304 4387 12338 4391
rect 12014 4313 12048 4347
rect 12086 4313 12120 4347
rect 12630 4571 12664 4605
rect 12702 4571 12736 4605
rect 12788 4559 12820 4593
rect 12820 4559 12822 4593
rect 12860 4559 12888 4593
rect 12888 4559 12894 4593
rect 13154 4593 13188 4602
rect 13226 4593 13260 4602
rect 13154 4568 13172 4593
rect 13172 4568 13188 4593
rect 13226 4568 13240 4593
rect 13240 4568 13260 4593
rect 13298 4568 13332 4602
rect 11623 4155 11657 4189
rect 11695 4155 11729 4189
rect 11767 4155 11801 4189
rect 11839 4155 11873 4189
rect 11911 4155 11945 4189
rect 11983 4155 12017 4189
rect 12055 4155 12089 4189
rect 12127 4155 12161 4189
rect 12199 4155 12233 4189
rect 12271 4155 12305 4189
rect 12343 4155 12377 4189
rect 12488 4307 12522 4341
rect 12560 4323 12594 4341
rect 12560 4307 12594 4323
rect 12840 4313 12874 4347
rect 12912 4323 12946 4347
rect 12912 4313 12946 4323
rect 13230 4313 13264 4347
rect 13302 4313 13336 4347
rect 17719 4304 17753 4338
rect 17791 4304 17821 4338
rect 17821 4304 17825 4338
rect 17863 4304 17889 4338
rect 17889 4304 17897 4338
rect 17935 4304 17957 4338
rect 17957 4304 17969 4338
rect 18007 4304 18025 4338
rect 18025 4304 18041 4338
rect 18079 4304 18093 4338
rect 18093 4304 18113 4338
rect 18151 4304 18161 4338
rect 18161 4304 18185 4338
rect 18223 4304 18229 4338
rect 18229 4304 18257 4338
rect 18295 4304 18297 4338
rect 18297 4304 18329 4338
rect 18367 4304 18399 4338
rect 18399 4304 18401 4338
rect 18439 4304 18467 4338
rect 18467 4304 18473 4338
rect 18511 4304 18535 4338
rect 18535 4304 18545 4338
rect 18583 4304 18603 4338
rect 18603 4304 18617 4338
rect 18655 4304 18671 4338
rect 18671 4304 18689 4338
rect 18727 4304 18739 4338
rect 18739 4304 18761 4338
rect 18799 4304 18807 4338
rect 18807 4304 18833 4338
rect 18871 4304 18875 4338
rect 18875 4304 18905 4338
rect 18943 4304 18977 4338
rect 19015 4304 19045 4338
rect 19045 4304 19049 4338
rect 19087 4304 19113 4338
rect 19113 4304 19121 4338
rect 19159 4304 19181 4338
rect 19181 4304 19193 4338
rect 19231 4304 19249 4338
rect 19249 4304 19265 4338
rect 12990 4155 13024 4189
rect 13062 4155 13096 4189
rect 12568 4036 12602 4070
rect 12640 4036 12650 4070
rect 12650 4036 12674 4070
rect 12884 3979 12918 4013
rect 12956 3979 12990 4013
rect 13148 4155 13182 4189
rect 13220 4155 13254 4189
rect 13475 4155 13509 4189
rect 13547 4155 13581 4189
rect 12816 3797 12850 3816
rect 12850 3797 12994 3816
rect 12816 3763 12994 3797
rect 12816 3729 12850 3763
rect 12850 3729 12994 3763
rect 12816 3695 12994 3729
rect 12816 3661 12850 3695
rect 12850 3661 12994 3695
rect 12816 3638 12994 3661
rect 12299 3395 12333 3429
rect 12371 3404 12386 3429
rect 12386 3404 12405 3429
rect 12371 3395 12405 3404
rect 13286 3942 13320 3976
rect 13358 3959 13392 3976
rect 13358 3942 13392 3959
rect 13710 3964 13744 3974
rect 13710 3940 13744 3964
rect 13710 3896 13744 3902
rect 13710 3868 13744 3896
rect 13192 3782 13226 3816
rect 13192 3710 13226 3744
rect 13192 3638 13226 3672
rect 13498 3797 13612 3816
rect 13612 3797 13646 3816
rect 13646 3797 13676 3816
rect 13498 3763 13676 3797
rect 13498 3729 13612 3763
rect 13612 3729 13646 3763
rect 13646 3729 13676 3763
rect 13498 3695 13676 3729
rect 13498 3661 13612 3695
rect 13612 3661 13646 3695
rect 13646 3661 13676 3695
rect 13498 3638 13676 3661
rect 13866 3794 13900 3816
rect 13866 3782 13900 3794
rect 13866 3726 13900 3744
rect 13866 3710 13900 3726
rect 13866 3658 13900 3672
rect 13866 3638 13900 3658
rect 14178 3794 14212 3816
rect 14178 3782 14212 3794
rect 14178 3726 14212 3744
rect 14178 3710 14212 3726
rect 14178 3658 14212 3672
rect 14178 3638 14212 3658
rect 14490 3794 14524 3816
rect 14490 3782 14524 3794
rect 14490 3726 14524 3744
rect 14490 3710 14524 3726
rect 14490 3658 14524 3672
rect 14490 3638 14524 3658
rect 14802 3794 14836 3816
rect 14802 3782 14836 3794
rect 14802 3726 14836 3744
rect 14802 3710 14836 3726
rect 14802 3658 14836 3672
rect 14802 3638 14836 3658
rect 15068 3797 15212 3816
rect 15212 3797 15246 3816
rect 15068 3794 15246 3797
rect 15068 3760 15114 3794
rect 15114 3760 15148 3794
rect 15148 3763 15246 3794
rect 15148 3760 15212 3763
rect 15068 3729 15212 3760
rect 15212 3729 15246 3763
rect 15068 3726 15246 3729
rect 15068 3692 15114 3726
rect 15114 3692 15148 3726
rect 15148 3695 15246 3726
rect 15148 3692 15212 3695
rect 15068 3661 15212 3692
rect 15212 3661 15246 3695
rect 15068 3658 15246 3661
rect 15068 3638 15114 3658
rect 15114 3638 15148 3658
rect 15148 3638 15246 3658
rect 15432 3862 15466 3896
rect 15504 3862 15538 3896
rect 15311 3574 15344 3592
rect 15344 3574 15345 3592
rect 15311 3558 15345 3574
rect 15383 3558 15417 3592
rect 15744 3862 15778 3896
rect 15816 3862 15850 3896
rect 15589 3574 15622 3592
rect 15622 3574 15623 3592
rect 15589 3558 15623 3574
rect 15661 3558 15695 3592
rect 16056 3862 16090 3896
rect 16128 3862 16162 3896
rect 13951 3032 13985 3066
rect 14023 3032 14057 3066
rect 14095 3032 14129 3066
rect 14167 3032 14201 3066
rect 14239 3032 14273 3066
rect 14311 3032 14345 3066
rect 14383 3032 14417 3066
rect 14455 3032 14489 3066
rect 14527 3032 14561 3066
rect 14599 3032 14633 3066
rect 14671 3032 14705 3066
rect 14743 3032 14777 3066
rect 14815 3032 14849 3066
rect 14887 3032 14921 3066
rect 14959 3032 14993 3066
rect 15031 3032 15065 3066
rect 15901 3574 15934 3592
rect 15934 3574 15935 3592
rect 15901 3558 15935 3574
rect 15973 3558 16007 3592
rect 16368 3862 16402 3896
rect 16440 3862 16474 3896
rect 16213 3574 16246 3592
rect 16246 3574 16247 3592
rect 16213 3558 16247 3574
rect 16285 3558 16319 3592
rect 16657 3797 16690 3816
rect 16690 3797 16835 3816
rect 16657 3794 16835 3797
rect 16657 3763 16754 3794
rect 16657 3729 16690 3763
rect 16690 3760 16754 3763
rect 16754 3760 16788 3794
rect 16788 3760 16835 3794
rect 16690 3729 16835 3760
rect 16657 3726 16835 3729
rect 16657 3695 16754 3726
rect 16657 3661 16690 3695
rect 16690 3692 16754 3695
rect 16754 3692 16788 3726
rect 16788 3692 16835 3726
rect 16690 3661 16835 3692
rect 16657 3658 16835 3661
rect 16657 3638 16754 3658
rect 16754 3638 16788 3658
rect 16788 3638 16835 3658
rect 16487 3558 16521 3592
rect 16559 3574 16592 3592
rect 16592 3574 16593 3592
rect 16559 3558 16593 3574
rect 17066 3794 17100 3816
rect 17066 3782 17100 3794
rect 17066 3726 17100 3744
rect 17066 3710 17100 3726
rect 17066 3658 17100 3672
rect 17066 3638 17100 3658
rect 16877 3590 16911 3592
rect 16877 3558 16910 3590
rect 16910 3558 16911 3590
rect 16949 3558 16983 3592
rect 17378 3794 17412 3816
rect 17378 3782 17412 3794
rect 17378 3726 17412 3744
rect 17378 3710 17412 3726
rect 17378 3658 17412 3672
rect 17378 3638 17412 3658
rect 17188 3558 17222 3592
rect 17260 3558 17294 3592
rect 17640 3794 17746 3816
rect 17640 3760 17690 3794
rect 17690 3760 17724 3794
rect 17724 3760 17746 3794
rect 17640 3726 17746 3760
rect 17640 3692 17690 3726
rect 17690 3692 17724 3726
rect 17724 3692 17746 3726
rect 17640 3658 17746 3692
rect 17640 3638 17690 3658
rect 17690 3638 17724 3658
rect 17724 3638 17746 3658
rect 17494 3558 17528 3592
rect 17566 3590 17600 3592
rect 17566 3558 17568 3590
rect 17568 3558 17600 3590
rect 17956 3797 18100 3816
rect 18100 3797 18134 3816
rect 17956 3794 18134 3797
rect 17956 3760 18002 3794
rect 18002 3760 18036 3794
rect 18036 3763 18134 3794
rect 18036 3760 18100 3763
rect 17956 3729 18100 3760
rect 18100 3729 18134 3763
rect 17956 3726 18134 3729
rect 17956 3692 18002 3726
rect 18002 3692 18036 3726
rect 18036 3695 18134 3726
rect 18036 3692 18100 3695
rect 17956 3661 18100 3692
rect 18100 3661 18134 3695
rect 17956 3658 18134 3661
rect 17956 3638 18002 3658
rect 18002 3638 18036 3658
rect 18036 3638 18134 3658
rect 17812 3558 17846 3592
rect 17884 3558 17918 3592
rect 18198 3590 18232 3592
rect 18198 3558 18232 3590
rect 18270 3558 18304 3592
rect 18476 3558 18510 3592
rect 18548 3558 18582 3592
rect 18320 3422 18354 3456
rect 18392 3422 18426 3456
rect 18788 3558 18822 3592
rect 18860 3558 18894 3592
rect 19591 4160 19625 4189
rect 19663 4160 19697 4189
rect 19735 4160 19769 4189
rect 19807 4160 19841 4189
rect 19591 4155 19599 4160
rect 19599 4155 19625 4160
rect 19663 4155 19667 4160
rect 19667 4155 19697 4160
rect 19735 4155 19769 4160
rect 19807 4155 19837 4160
rect 19837 4155 19841 4160
rect 16830 3030 16864 3060
rect 16902 3030 16936 3060
rect 16974 3030 17008 3060
rect 17046 3030 17080 3060
rect 17118 3030 17152 3060
rect 17190 3030 17224 3060
rect 17262 3030 17296 3060
rect 17334 3030 17368 3060
rect 17406 3030 17440 3060
rect 17478 3030 17512 3060
rect 17550 3030 17584 3060
rect 17622 3030 17656 3060
rect 17694 3030 17728 3060
rect 17766 3030 17800 3060
rect 17838 3030 17872 3060
rect 17910 3030 17944 3060
rect 18631 3422 18665 3456
rect 18703 3422 18737 3456
rect 19100 3558 19134 3592
rect 18944 3336 18978 3370
rect 19172 3558 19206 3592
rect 19016 3336 19050 3370
rect 19374 3558 19408 3592
rect 19446 3590 19480 3592
rect 19446 3558 19480 3590
rect 19255 3336 19289 3370
rect 19327 3336 19361 3370
rect 19796 3862 19830 3896
rect 19868 3862 19902 3896
rect 19712 3794 19746 3816
rect 19712 3782 19746 3794
rect 19712 3726 19746 3744
rect 19712 3710 19746 3726
rect 19712 3658 19746 3672
rect 19712 3638 19746 3658
rect 19556 3352 19590 3370
rect 19556 3336 19590 3352
rect 19628 3336 19662 3370
rect 16830 3026 16833 3030
rect 16833 3026 16864 3030
rect 16902 3026 16935 3030
rect 16935 3026 16936 3030
rect 16974 3026 17003 3030
rect 17003 3026 17008 3030
rect 17046 3026 17071 3030
rect 17071 3026 17080 3030
rect 17118 3026 17139 3030
rect 17139 3026 17152 3030
rect 17190 3026 17207 3030
rect 17207 3026 17224 3030
rect 17262 3026 17275 3030
rect 17275 3026 17296 3030
rect 17334 3026 17343 3030
rect 17343 3026 17368 3030
rect 17406 3026 17411 3030
rect 17411 3026 17440 3030
rect 17478 3026 17479 3030
rect 17479 3026 17512 3030
rect 17550 3026 17581 3030
rect 17581 3026 17584 3030
rect 17622 3026 17649 3030
rect 17649 3026 17656 3030
rect 17694 3026 17717 3030
rect 17717 3026 17728 3030
rect 17766 3026 17785 3030
rect 17785 3026 17800 3030
rect 17838 3026 17853 3030
rect 17853 3026 17872 3030
rect 17910 3026 17921 3030
rect 17921 3026 17944 3030
rect 15401 2980 15435 2982
rect 15473 2980 15507 2982
rect 15545 2980 15579 2982
rect 15617 2980 15651 2982
rect 15689 2980 15723 2982
rect 15761 2980 15795 2982
rect 15833 2980 15867 2982
rect 15905 2980 15939 2982
rect 15977 2980 16011 2982
rect 16049 2980 16083 2982
rect 16121 2980 16155 2982
rect 16193 2980 16227 2982
rect 16265 2980 16299 2982
rect 16337 2980 16371 2982
rect 16409 2980 16443 2982
rect 16481 2980 16515 2982
rect 15401 2948 15423 2980
rect 15423 2948 15435 2980
rect 15473 2948 15491 2980
rect 15491 2948 15507 2980
rect 15545 2948 15559 2980
rect 15559 2948 15579 2980
rect 15617 2948 15627 2980
rect 15627 2948 15651 2980
rect 15689 2948 15695 2980
rect 15695 2948 15723 2980
rect 15761 2948 15763 2980
rect 15763 2948 15795 2980
rect 15833 2948 15865 2980
rect 15865 2948 15867 2980
rect 15905 2948 15933 2980
rect 15933 2948 15939 2980
rect 15977 2948 16001 2980
rect 16001 2948 16011 2980
rect 16049 2948 16069 2980
rect 16069 2948 16083 2980
rect 16121 2948 16137 2980
rect 16137 2948 16155 2980
rect 16193 2948 16205 2980
rect 16205 2948 16227 2980
rect 16265 2948 16273 2980
rect 16273 2948 16299 2980
rect 16337 2948 16341 2980
rect 16341 2948 16371 2980
rect 16409 2948 16443 2980
rect 16481 2948 16511 2980
rect 16511 2948 16515 2980
<< metal1 >>
rect 7363 6416 8033 6428
rect 7363 6382 7369 6416
rect 7403 6382 7681 6416
rect 7715 6382 7993 6416
rect 8027 6382 8033 6416
rect 7363 6344 8033 6382
rect 7363 6310 7369 6344
rect 7403 6310 7681 6344
rect 7715 6310 7993 6344
rect 8027 6310 8033 6344
rect 7363 6272 8033 6310
rect 7363 6238 7369 6272
rect 7403 6238 7681 6272
rect 7715 6238 7993 6272
rect 8027 6238 8033 6272
rect 7363 6226 8033 6238
rect 7831 5967 7877 5979
rect 7831 5933 7837 5967
rect 7871 5933 7877 5967
rect 7831 5895 7877 5933
rect 7831 5861 7837 5895
rect 7871 5861 7877 5895
rect 7831 5823 7877 5861
rect 7831 5789 7837 5823
rect 7871 5789 7877 5823
rect 7831 5777 7877 5789
rect 7519 5580 7565 5592
rect 7519 5546 7525 5580
rect 7559 5546 7565 5580
rect 7519 5504 7565 5546
rect 7519 5470 7525 5504
rect 7559 5470 7565 5504
rect 7519 5428 7565 5470
rect 7519 5394 7525 5428
rect 7559 5394 7565 5428
rect 7519 5351 7565 5394
rect 7519 5317 7525 5351
rect 7559 5317 7565 5351
rect 7519 5274 7565 5317
rect 7519 5240 7525 5274
rect 7559 5240 7565 5274
rect 11364 5441 13508 5453
rect 11364 5407 12304 5441
rect 12338 5407 13508 5441
rect 11364 5369 13508 5407
rect 11364 5335 12304 5369
rect 12338 5335 13508 5369
rect 11364 5297 13508 5335
rect 11364 5263 12304 5297
rect 12338 5263 13508 5297
rect 11364 5251 13508 5263
rect 7519 5197 7565 5240
rect 7519 5163 7525 5197
rect 7559 5163 7565 5197
rect 7519 5120 7565 5163
rect 7519 5086 7525 5120
rect 7559 5086 7565 5120
tri 7516 5052 7519 5055 se
rect 7519 5052 7565 5086
rect 7751 5197 10441 5212
tri 10441 5197 10456 5212 sw
rect 7751 5163 7757 5197
rect 7791 5163 7913 5197
rect 7947 5163 10456 5197
rect 7751 5160 10456 5163
rect 7751 5125 7797 5160
rect 7751 5091 7757 5125
rect 7791 5091 7797 5125
rect 7751 5079 7797 5091
rect 7907 5125 7953 5160
tri 10419 5132 10447 5160 ne
rect 10447 5132 10456 5160
rect 7907 5091 7913 5125
rect 7947 5091 7953 5125
rect 7907 5079 7953 5091
rect 9831 5080 9837 5132
rect 9889 5080 9901 5132
rect 9953 5123 10316 5132
tri 10316 5123 10325 5132 sw
tri 10447 5123 10456 5132 ne
tri 10456 5123 10530 5197 sw
rect 9953 5105 10325 5123
tri 10325 5105 10343 5123 sw
tri 10456 5105 10474 5123 ne
rect 10474 5105 10595 5123
rect 9953 5080 10343 5105
tri 10306 5079 10307 5080 ne
rect 10307 5079 10343 5080
tri 10343 5079 10369 5105 sw
tri 10474 5079 10500 5105 ne
rect 10500 5079 10595 5105
tri 10307 5055 10331 5079 ne
rect 10331 5071 10369 5079
tri 10369 5071 10377 5079 sw
tri 10500 5071 10508 5079 ne
rect 10508 5071 10595 5079
rect 10647 5071 10659 5123
rect 10711 5071 10717 5123
rect 10331 5055 10377 5071
tri 7565 5052 7568 5055 sw
rect 7516 5046 7568 5052
tri 10331 5043 10343 5055 ne
rect 10343 5050 10377 5055
tri 10377 5050 10398 5071 sw
rect 10343 5043 10398 5050
tri 10398 5043 10405 5050 sw
tri 13053 5043 13060 5050 se
rect 13060 5043 13066 5050
tri 10343 4998 10388 5043 ne
rect 10388 4998 13066 5043
rect 13118 4998 13130 5050
rect 13182 4998 13188 5050
rect 7516 4972 7568 4994
rect 7516 4898 7568 4920
rect 7516 4840 7568 4846
rect 11364 4957 13508 4969
rect 11364 4851 12296 4957
rect 12402 4879 13508 4957
rect 12402 4851 12841 4879
rect 11364 4845 12841 4851
rect 12875 4845 12913 4879
rect 12947 4845 12985 4879
rect 13019 4845 13508 4879
rect 11364 4839 13508 4845
rect 11523 4805 13504 4811
rect 11523 4771 11538 4805
rect 11572 4771 11610 4805
rect 11644 4771 11682 4805
rect 11716 4771 11754 4805
rect 11788 4771 11826 4805
rect 11860 4771 11898 4805
rect 11932 4771 11970 4805
rect 12004 4771 13386 4805
rect 13420 4771 13458 4805
rect 13492 4771 13504 4805
rect 11523 4765 13504 4771
tri 9157 4735 9182 4760 se
rect 9182 4735 9837 4760
rect 7420 4725 8769 4735
rect 7420 4691 7438 4725
rect 7472 4691 7530 4725
rect 7564 4691 7623 4725
rect 7657 4691 8769 4725
rect 7420 4683 8769 4691
rect 8821 4683 8833 4735
rect 8885 4683 8891 4735
tri 9130 4708 9157 4735 se
rect 9157 4708 9837 4735
rect 9889 4708 9901 4760
rect 9953 4708 9959 4760
rect 11523 4740 12023 4765
tri 12023 4740 12048 4765 nw
tri 12593 4740 12618 4765 ne
rect 11524 4738 12022 4739
tri 9122 4700 9130 4708 se
rect 9130 4700 9196 4708
tri 9196 4700 9204 4708 nw
rect 11524 4701 12022 4702
tri 9108 4686 9122 4700 se
rect 9122 4686 9182 4700
tri 9182 4686 9196 4700 nw
tri 9105 4683 9108 4686 se
rect 9108 4683 9171 4686
tri 9097 4675 9105 4683 se
rect 9105 4675 9171 4683
tri 9171 4675 9182 4686 nw
rect 11523 4675 12023 4700
tri 12023 4675 12048 4700 sw
tri 9085 4663 9097 4675 se
rect 9097 4663 9159 4675
tri 9159 4663 9171 4675 nw
tri 9051 4629 9085 4663 se
rect 9085 4629 9125 4663
tri 9125 4629 9159 4663 nw
tri 9045 4623 9051 4629 se
rect 9051 4623 9119 4629
tri 9119 4623 9125 4629 nw
rect 11523 4623 11529 4675
rect 11581 4623 11593 4675
rect 11645 4663 12258 4675
rect 11645 4629 11682 4663
rect 11716 4629 11754 4663
rect 11788 4629 11826 4663
rect 11860 4629 11898 4663
rect 11932 4629 11970 4663
rect 12004 4629 12258 4663
rect 11645 4623 12258 4629
tri 9034 4612 9045 4623 se
rect 9045 4612 9108 4623
tri 9108 4612 9119 4623 nw
tri 9033 4611 9034 4612 se
rect 9034 4611 9107 4612
tri 9107 4611 9108 4612 nw
tri 9027 4605 9033 4611 se
rect 9033 4605 9101 4611
tri 9101 4605 9107 4611 nw
rect 12618 4605 12748 4765
tri 12748 4740 12773 4765 nw
tri 9021 4599 9027 4605 se
rect 9027 4599 9095 4605
tri 9095 4599 9101 4605 nw
tri 9017 4595 9021 4599 se
rect 9021 4595 9091 4599
tri 9091 4595 9095 4599 nw
tri 9009 4587 9017 4595 se
rect 9017 4587 9083 4595
tri 9083 4587 9091 4595 nw
tri 8975 4553 9009 4587 se
rect 9009 4553 9049 4587
tri 9049 4553 9083 4587 nw
tri 8965 4543 8975 4553 se
rect 8975 4543 9039 4553
tri 9039 4543 9049 4553 nw
rect 11612 4543 11618 4595
rect 11670 4543 11682 4595
rect 11734 4587 12174 4595
rect 11734 4553 12056 4587
rect 12090 4553 12128 4587
rect 12162 4553 12174 4587
rect 12618 4571 12630 4605
rect 12664 4571 12702 4605
rect 12736 4571 12748 4605
rect 12618 4565 12748 4571
rect 12776 4636 13508 4682
rect 12776 4593 12906 4636
tri 12906 4611 12931 4636 nw
tri 13052 4602 13058 4608 se
rect 13058 4602 13222 4608
tri 13049 4599 13052 4602 se
rect 13052 4599 13154 4602
tri 13045 4595 13049 4599 se
rect 13049 4595 13154 4599
rect 12776 4559 12788 4593
rect 12822 4559 12860 4593
rect 12894 4559 12906 4593
tri 13018 4568 13045 4595 se
rect 13045 4568 13154 4595
rect 13188 4568 13222 4602
rect 12776 4553 12906 4559
tri 13006 4556 13018 4568 se
rect 13018 4556 13222 4568
rect 13274 4556 13286 4608
rect 13338 4556 13348 4608
tri 13003 4553 13006 4556 se
rect 13006 4553 13067 4556
rect 11734 4543 12174 4553
tri 12993 4543 13003 4553 se
rect 13003 4543 13067 4553
tri 13067 4543 13080 4556 nw
tri 8960 4538 8965 4543 se
rect 8965 4538 9034 4543
tri 9034 4538 9039 4543 nw
tri 12988 4538 12993 4543 se
rect 12993 4538 13062 4543
tri 13062 4538 13067 4543 nw
tri 8937 4515 8960 4538 se
rect 8960 4515 9011 4538
tri 9011 4515 9034 4538 nw
tri 12985 4535 12988 4538 se
rect 12988 4535 13059 4538
tri 13059 4535 13062 4538 nw
tri 12965 4515 12985 4535 se
rect 12985 4515 13039 4535
tri 13039 4515 13059 4535 nw
rect 7564 4513 9009 4515
tri 9009 4513 9011 4515 nw
tri 12963 4513 12965 4515 se
rect 12965 4513 13037 4515
tri 13037 4513 13039 4515 nw
rect 7564 4508 8959 4513
rect 7564 4474 7584 4508
rect 7618 4474 7671 4508
rect 7705 4474 7758 4508
rect 7792 4474 7846 4508
rect 7880 4474 7934 4508
rect 7968 4474 8959 4508
rect 7564 4463 8959 4474
tri 8959 4463 9009 4513 nw
rect 10589 4461 10595 4513
rect 10647 4461 10659 4513
rect 10711 4461 12985 4513
tri 12985 4461 13037 4513 nw
rect 7669 4422 10278 4433
rect 7669 4421 7943 4422
rect 7669 4387 7675 4421
rect 7709 4388 7943 4421
rect 7977 4388 8015 4422
rect 8049 4388 10278 4422
rect 7709 4387 10278 4388
rect 7669 4381 10278 4387
rect 10330 4381 10342 4433
rect 10394 4381 10400 4433
rect 11706 4425 11839 4433
rect 11841 4432 11877 4433
rect 11706 4391 11718 4425
rect 11752 4391 11790 4425
rect 11824 4391 11839 4425
rect 11706 4381 11839 4391
rect 11840 4382 11878 4432
rect 11879 4421 12478 4433
rect 11879 4387 12232 4421
rect 12266 4387 12304 4421
rect 12338 4387 12478 4421
rect 11841 4381 11877 4382
rect 11879 4381 12478 4387
rect 12530 4381 12542 4433
rect 12594 4381 12600 4433
rect 7669 4349 7715 4381
rect 16384 4353 18188 4459
rect 7669 4315 7675 4349
rect 7709 4315 7715 4349
rect 7669 4303 7715 4315
rect 11364 4347 16355 4353
rect 11364 4313 11548 4347
rect 11582 4313 11620 4347
rect 11654 4313 12014 4347
rect 12048 4313 12086 4347
rect 12120 4341 12840 4347
rect 12120 4313 12488 4341
rect 11364 4307 12488 4313
rect 12522 4307 12560 4341
rect 12594 4313 12840 4341
rect 12874 4313 12912 4347
rect 12946 4313 13230 4347
rect 13264 4313 13302 4347
rect 13336 4313 16355 4347
rect 16384 4338 20028 4353
rect 16384 4329 17719 4338
rect 12594 4307 16355 4313
rect 11364 4223 16355 4307
rect 17701 4304 17719 4329
rect 17753 4304 17791 4338
rect 17825 4304 17863 4338
rect 17897 4304 17935 4338
rect 17969 4304 18007 4338
rect 18041 4304 18079 4338
rect 18113 4304 18151 4338
rect 18185 4304 18223 4338
rect 18257 4304 18295 4338
rect 18329 4304 18367 4338
rect 18401 4304 18439 4338
rect 18473 4304 18511 4338
rect 18545 4304 18583 4338
rect 18617 4304 18655 4338
rect 18689 4304 18727 4338
rect 18761 4304 18799 4338
rect 18833 4304 18871 4338
rect 18905 4304 18943 4338
rect 18977 4304 19015 4338
rect 19049 4304 19087 4338
rect 19121 4304 19159 4338
rect 19193 4304 19231 4338
rect 19265 4304 20028 4338
rect 17701 4223 20028 4304
rect 7513 4180 7871 4186
rect 7513 4128 7516 4180
rect 7568 4174 7871 4180
rect 7568 4140 7831 4174
rect 7865 4140 7871 4174
rect 10272 4143 10278 4195
rect 10330 4143 10342 4195
rect 10394 4160 11401 4195
rect 11589 4189 13108 4195
rect 10394 4155 10412 4160
tri 10412 4155 10417 4160 nw
rect 11589 4155 11623 4189
rect 11657 4155 11695 4189
rect 11729 4155 11767 4189
rect 11801 4155 11839 4189
rect 11873 4155 11911 4189
rect 11945 4155 11983 4189
rect 12017 4155 12055 4189
rect 12089 4155 12127 4189
rect 12161 4155 12199 4189
rect 12233 4155 12271 4189
rect 12305 4155 12343 4189
rect 12377 4155 12990 4189
rect 13024 4155 13062 4189
rect 13096 4155 13108 4189
rect 10394 4143 10400 4155
tri 10400 4143 10412 4155 nw
rect 11589 4149 13108 4155
tri 12531 4143 12537 4149 ne
rect 12537 4143 12705 4149
tri 12705 4143 12711 4149 nw
rect 13136 4143 13142 4195
rect 13194 4143 13206 4195
rect 13258 4143 13266 4195
rect 13463 4189 19854 4195
rect 13463 4155 13475 4189
rect 13509 4155 13547 4189
rect 13581 4155 19591 4189
rect 19625 4155 19663 4189
rect 19697 4155 19735 4189
rect 19769 4155 19807 4189
rect 19841 4155 19854 4189
rect 13463 4149 19854 4155
rect 7568 4128 7871 4140
rect 7513 4114 7871 4128
tri 12537 4124 12556 4143 ne
rect 12556 4124 12686 4143
tri 12686 4124 12705 4143 nw
rect 7513 4062 7516 4114
rect 7568 4062 7871 4114
rect 7513 4047 7871 4062
rect 7513 3995 7516 4047
rect 7568 4033 7871 4047
rect 7568 3999 7831 4033
rect 7865 3999 7871 4033
rect 12557 4122 12685 4123
rect 12556 4086 12686 4122
rect 12557 4085 12685 4086
rect 12556 4070 12686 4084
rect 12556 4036 12568 4070
rect 12602 4036 12640 4070
rect 12674 4036 12686 4070
rect 12556 4030 12686 4036
rect 7568 3995 7871 3999
rect 7513 3987 7871 3995
rect 12872 4013 13002 4025
rect 12872 3979 12884 4013
rect 12918 3979 12956 4013
rect 12990 3979 13002 4013
rect 12872 3973 13002 3979
rect 12873 3971 13001 3972
rect 12872 3935 13002 3971
rect 13274 3976 13404 3982
rect 13274 3942 13286 3976
rect 13320 3942 13358 3976
rect 13392 3942 13404 3976
rect 13274 3936 13404 3942
rect 13704 3974 13750 3986
rect 13704 3940 13710 3974
rect 13744 3940 13750 3974
rect 12873 3934 13001 3935
tri 12847 3908 12872 3933 se
rect 12872 3908 13002 3933
tri 13002 3908 13027 3933 sw
tri 13679 3908 13704 3933 se
rect 13704 3908 13750 3940
tri 13750 3908 13775 3933 sw
rect 11428 3856 12478 3908
rect 12530 3856 12542 3908
rect 12594 3902 19963 3908
rect 12594 3868 13710 3902
rect 13744 3896 19963 3902
rect 13744 3868 15432 3896
rect 12594 3862 15432 3868
rect 15466 3862 15504 3896
rect 15538 3862 15744 3896
rect 15778 3862 15816 3896
rect 15850 3862 16056 3896
rect 16090 3862 16128 3896
rect 16162 3862 16368 3896
rect 16402 3862 16440 3896
rect 16474 3862 19796 3896
rect 19830 3862 19868 3896
rect 19902 3862 19963 3896
rect 12594 3856 19963 3862
rect 11364 3816 19985 3828
rect 11364 3638 12816 3816
rect 12994 3782 13192 3816
rect 13226 3782 13498 3816
rect 12994 3744 13498 3782
rect 12994 3710 13192 3744
rect 13226 3710 13498 3744
rect 12994 3672 13498 3710
rect 12994 3638 13192 3672
rect 13226 3638 13498 3672
rect 13676 3782 13866 3816
rect 13900 3782 14178 3816
rect 14212 3782 14490 3816
rect 14524 3782 14802 3816
rect 14836 3782 15068 3816
rect 13676 3744 15068 3782
rect 13676 3710 13866 3744
rect 13900 3710 14178 3744
rect 14212 3710 14490 3744
rect 14524 3710 14802 3744
rect 14836 3710 15068 3744
rect 13676 3672 15068 3710
rect 13676 3638 13866 3672
rect 13900 3638 14178 3672
rect 14212 3638 14490 3672
rect 14524 3638 14802 3672
rect 14836 3638 15068 3672
rect 15246 3638 16657 3816
rect 16835 3782 17066 3816
rect 17100 3782 17378 3816
rect 17412 3782 17640 3816
rect 16835 3744 17640 3782
rect 16835 3710 17066 3744
rect 17100 3710 17378 3744
rect 17412 3710 17640 3744
rect 16835 3672 17640 3710
rect 16835 3638 17066 3672
rect 17100 3638 17378 3672
rect 17412 3638 17640 3672
rect 17746 3638 17956 3816
rect 18134 3782 19712 3816
rect 19746 3782 19985 3816
rect 18134 3744 19985 3782
rect 18134 3710 19712 3744
rect 19746 3710 19985 3744
rect 18134 3672 19985 3710
rect 18134 3638 19712 3672
rect 19746 3638 19985 3672
rect 11364 3626 19985 3638
rect 8763 3546 8769 3598
rect 8821 3546 8833 3598
rect 8885 3592 10630 3598
tri 10630 3592 10636 3598 sw
rect 8885 3564 10636 3592
rect 8885 3558 8903 3564
tri 8903 3558 8909 3564 nw
tri 10590 3558 10596 3564 ne
rect 10596 3558 10636 3564
tri 10636 3558 10670 3592 sw
rect 8885 3555 8900 3558
tri 8900 3555 8903 3558 nw
tri 10596 3555 10599 3558 ne
rect 10599 3555 10670 3558
tri 10670 3555 10673 3558 sw
rect 8885 3546 8891 3555
tri 8891 3546 8900 3555 nw
tri 10599 3546 10608 3555 ne
rect 10608 3546 10673 3555
tri 10673 3546 10682 3555 sw
rect 11523 3546 11529 3598
rect 11581 3546 11593 3598
rect 11645 3546 13250 3598
tri 10608 3524 10630 3546 ne
rect 10630 3524 10682 3546
tri 10630 3481 10673 3524 ne
rect 10673 3518 10682 3524
tri 10682 3518 10710 3546 sw
tri 13104 3518 13132 3546 ne
rect 13132 3518 13250 3546
rect 10673 3481 10710 3518
tri 10710 3481 10747 3518 sw
tri 10673 3456 10698 3481 ne
rect 10698 3466 10962 3481
tri 10962 3466 10977 3481 sw
rect 11612 3466 11618 3518
rect 11670 3466 11682 3518
rect 11734 3516 13092 3518
tri 13092 3516 13094 3518 sw
tri 13132 3516 13134 3518 ne
rect 13134 3516 13250 3518
rect 11734 3506 13094 3516
tri 13094 3506 13104 3516 sw
tri 13134 3506 13144 3516 ne
rect 13144 3506 13250 3516
rect 11734 3470 13104 3506
tri 13104 3470 13140 3506 sw
tri 13144 3470 13180 3506 ne
rect 13180 3470 13250 3506
rect 13251 3471 13252 3597
rect 13288 3471 13289 3597
rect 13290 3592 13346 3598
rect 13290 3540 13292 3592
rect 13344 3540 13346 3592
rect 15299 3592 16796 3598
rect 16798 3597 16834 3598
rect 15299 3558 15311 3592
rect 15345 3558 15383 3592
rect 15417 3558 15589 3592
rect 15623 3558 15661 3592
rect 15695 3558 15901 3592
rect 15935 3558 15973 3592
rect 16007 3558 16213 3592
rect 16247 3558 16285 3592
rect 16319 3558 16487 3592
rect 16521 3558 16559 3592
rect 16593 3558 16796 3592
rect 15299 3552 16796 3558
rect 16797 3553 16835 3597
rect 16836 3592 17930 3598
rect 16836 3558 16877 3592
rect 16911 3558 16949 3592
rect 16983 3558 17188 3592
rect 17222 3558 17260 3592
rect 17294 3558 17494 3592
rect 17528 3558 17566 3592
rect 17600 3558 17812 3592
rect 17846 3558 17884 3592
rect 17918 3558 17930 3592
rect 16798 3552 16834 3553
rect 16836 3552 17930 3558
rect 18186 3592 19492 3598
rect 18186 3558 18198 3592
rect 18232 3558 18270 3592
rect 18304 3558 18476 3592
rect 18510 3558 18548 3592
rect 18582 3558 18788 3592
rect 18822 3558 18860 3592
rect 18894 3558 19100 3592
rect 19134 3558 19172 3592
rect 19206 3558 19374 3592
rect 19408 3558 19446 3592
rect 19480 3558 19492 3592
rect 18186 3552 19492 3558
rect 13290 3528 13346 3540
rect 13290 3476 13292 3528
rect 13344 3476 13346 3528
rect 13290 3470 13346 3476
rect 11734 3466 13140 3470
rect 10698 3456 10977 3466
tri 10977 3456 10987 3466 sw
tri 13070 3456 13080 3466 ne
rect 13080 3462 13140 3466
tri 13140 3462 13148 3470 sw
rect 13080 3456 13148 3462
tri 13148 3456 13154 3462 sw
tri 13474 3456 13480 3462 se
rect 13480 3456 18749 3462
tri 10698 3438 10716 3456 ne
rect 10716 3442 10987 3456
tri 10987 3442 11001 3456 sw
tri 13080 3442 13094 3456 ne
rect 13094 3442 13154 3456
tri 13154 3442 13168 3456 sw
tri 13460 3442 13474 3456 se
rect 13474 3442 18320 3456
rect 10716 3438 11001 3442
tri 11001 3438 11005 3442 sw
tri 13094 3438 13098 3442 ne
rect 13098 3438 18320 3442
tri 10716 3429 10725 3438 ne
rect 10725 3429 11529 3438
tri 10940 3395 10974 3429 ne
rect 10974 3395 11529 3429
tri 10974 3386 10983 3395 ne
rect 10983 3386 11529 3395
rect 11581 3386 11593 3438
rect 11645 3386 11680 3438
rect 11682 3437 11718 3438
rect 11681 3387 11719 3437
rect 11720 3429 12417 3438
rect 11720 3395 12299 3429
rect 12333 3395 12371 3429
rect 12405 3395 12417 3429
tri 13098 3422 13114 3438 ne
rect 13114 3422 18320 3438
rect 18354 3422 18392 3456
rect 18426 3422 18631 3456
rect 18665 3422 18703 3456
rect 18737 3422 18749 3456
rect 11682 3386 11718 3387
rect 11720 3386 12417 3395
tri 13114 3390 13146 3422 ne
rect 13146 3410 18749 3422
rect 13146 3390 13482 3410
tri 13482 3390 13502 3410 nw
rect 17190 3330 17196 3382
rect 17248 3330 17260 3382
rect 17312 3370 19674 3382
rect 17312 3336 18944 3370
rect 18978 3336 19016 3370
rect 19050 3336 19255 3370
rect 19289 3336 19327 3370
rect 19361 3336 19556 3370
rect 19590 3336 19628 3370
rect 19662 3336 19674 3370
rect 17312 3330 19674 3336
rect 11364 3100 19871 3302
rect 13939 3066 15140 3072
rect 13939 3032 13951 3066
rect 13985 3032 14023 3066
rect 14057 3032 14095 3066
rect 14129 3032 14167 3066
rect 14201 3032 14239 3066
rect 14273 3032 14311 3066
rect 14345 3032 14383 3066
rect 14417 3032 14455 3066
rect 14489 3032 14527 3066
rect 14561 3032 14599 3066
rect 14633 3032 14671 3066
rect 14705 3032 14743 3066
rect 14777 3032 14815 3066
rect 14849 3032 14887 3066
rect 14921 3032 14959 3066
rect 14993 3032 15031 3066
rect 15065 3032 15140 3066
rect 13939 3026 15140 3032
rect 15141 3027 15142 3071
rect 15178 3027 15179 3071
rect 15180 3060 15316 3072
tri 15316 3060 15328 3072 sw
rect 16818 3060 17196 3072
rect 15180 3026 15328 3060
tri 15328 3026 15362 3060 sw
rect 16818 3026 16830 3060
rect 16864 3026 16902 3060
rect 16936 3026 16974 3060
rect 17008 3026 17046 3060
rect 17080 3026 17118 3060
rect 17152 3026 17190 3060
tri 15296 2982 15340 3026 ne
rect 15340 2988 15362 3026
tri 15362 2988 15400 3026 sw
rect 16818 3020 17196 3026
rect 17248 3020 17260 3072
rect 17312 3060 17956 3072
rect 17312 3026 17334 3060
rect 17368 3026 17406 3060
rect 17440 3026 17478 3060
rect 17512 3026 17550 3060
rect 17584 3026 17622 3060
rect 17656 3026 17694 3060
rect 17728 3026 17766 3060
rect 17800 3026 17838 3060
rect 17872 3026 17910 3060
rect 17944 3026 17956 3060
rect 17312 3020 17956 3026
rect 15340 2982 16527 2988
tri 15340 2960 15362 2982 ne
rect 15362 2960 15401 2982
tri 15362 2948 15374 2960 ne
rect 15374 2948 15401 2960
rect 15435 2948 15473 2982
rect 15507 2948 15545 2982
rect 15579 2948 15617 2982
rect 15651 2948 15689 2982
rect 15723 2948 15761 2982
rect 15795 2948 15833 2982
rect 15867 2948 15905 2982
rect 15939 2948 15977 2982
rect 16011 2948 16049 2982
rect 16083 2948 16121 2982
rect 16155 2948 16193 2982
rect 16227 2948 16265 2982
rect 16299 2948 16337 2982
rect 16371 2948 16409 2982
rect 16443 2948 16481 2982
rect 16515 2948 16527 2982
tri 15374 2942 15380 2948 ne
rect 15380 2942 16527 2948
<< rmetal1 >>
rect 11523 4739 12023 4740
rect 11523 4738 11524 4739
rect 12022 4738 12023 4739
rect 11523 4701 11524 4702
rect 12022 4701 12023 4702
rect 11523 4700 12023 4701
rect 11839 4432 11841 4433
rect 11877 4432 11879 4433
rect 11839 4382 11840 4432
rect 11878 4382 11879 4432
rect 11839 4381 11841 4382
rect 11877 4381 11879 4382
rect 12556 4123 12686 4124
rect 12556 4122 12557 4123
rect 12685 4122 12686 4123
rect 12556 4085 12557 4086
rect 12685 4085 12686 4086
rect 12556 4084 12686 4085
rect 12872 3972 13002 3973
rect 12872 3971 12873 3972
rect 13001 3971 13002 3972
rect 12872 3934 12873 3935
rect 13001 3934 13002 3935
rect 12872 3933 13002 3934
rect 13250 3597 13252 3598
rect 13250 3471 13251 3597
rect 13250 3470 13252 3471
rect 13288 3597 13290 3598
rect 13289 3471 13290 3597
rect 16796 3597 16798 3598
rect 16834 3597 16836 3598
rect 16796 3553 16797 3597
rect 16835 3553 16836 3597
rect 16796 3552 16798 3553
rect 16834 3552 16836 3553
rect 13288 3470 13290 3471
rect 11680 3437 11682 3438
rect 11718 3437 11720 3438
rect 11680 3387 11681 3437
rect 11719 3387 11720 3437
rect 11680 3386 11682 3387
rect 11718 3386 11720 3387
rect 15140 3071 15142 3072
rect 15140 3027 15141 3071
rect 15140 3026 15142 3027
rect 15178 3071 15180 3072
rect 15179 3027 15180 3071
rect 15178 3026 15180 3027
<< via1 >>
rect 9837 5080 9889 5132
rect 9901 5080 9953 5132
rect 10595 5071 10647 5123
rect 10659 5071 10711 5123
rect 7516 5043 7568 5046
rect 7516 5009 7525 5043
rect 7525 5009 7559 5043
rect 7559 5009 7568 5043
rect 7516 4994 7568 5009
rect 13066 4998 13118 5050
rect 13130 4998 13182 5050
rect 7516 4966 7568 4972
rect 7516 4932 7525 4966
rect 7525 4932 7559 4966
rect 7559 4932 7568 4966
rect 7516 4920 7568 4932
rect 7516 4889 7568 4898
rect 7516 4855 7525 4889
rect 7525 4855 7559 4889
rect 7559 4855 7568 4889
rect 7516 4846 7568 4855
rect 8769 4683 8821 4735
rect 8833 4683 8885 4735
rect 9837 4708 9889 4760
rect 9901 4708 9953 4760
rect 11529 4663 11581 4675
rect 11529 4629 11538 4663
rect 11538 4629 11572 4663
rect 11572 4629 11581 4663
rect 11529 4623 11581 4629
rect 11593 4663 11645 4675
rect 11593 4629 11610 4663
rect 11610 4629 11644 4663
rect 11644 4629 11645 4663
rect 11593 4623 11645 4629
rect 11618 4543 11670 4595
rect 11682 4543 11734 4595
rect 13222 4602 13274 4608
rect 13222 4568 13226 4602
rect 13226 4568 13260 4602
rect 13260 4568 13274 4602
rect 13222 4556 13274 4568
rect 13286 4602 13338 4608
rect 13286 4568 13298 4602
rect 13298 4568 13332 4602
rect 13332 4568 13338 4602
rect 13286 4556 13338 4568
rect 10595 4461 10647 4513
rect 10659 4461 10711 4513
rect 10278 4381 10330 4433
rect 10342 4381 10394 4433
rect 12478 4381 12530 4433
rect 12542 4381 12594 4433
rect 7516 4174 7568 4180
rect 7516 4140 7519 4174
rect 7519 4140 7553 4174
rect 7553 4140 7568 4174
rect 10278 4143 10330 4195
rect 10342 4143 10394 4195
rect 13142 4189 13194 4195
rect 13142 4155 13148 4189
rect 13148 4155 13182 4189
rect 13182 4155 13194 4189
rect 13142 4143 13194 4155
rect 13206 4189 13258 4195
rect 13206 4155 13220 4189
rect 13220 4155 13254 4189
rect 13254 4155 13258 4189
rect 13206 4143 13258 4155
rect 7516 4128 7568 4140
rect 7516 4062 7568 4114
rect 7516 4033 7568 4047
rect 7516 3999 7519 4033
rect 7519 3999 7553 4033
rect 7553 3999 7568 4033
rect 7516 3995 7568 3999
rect 12478 3856 12530 3908
rect 12542 3856 12594 3908
rect 8769 3546 8821 3598
rect 8833 3546 8885 3598
rect 11529 3546 11581 3598
rect 11593 3546 11645 3598
rect 11618 3466 11670 3518
rect 11682 3466 11734 3518
rect 13292 3540 13344 3592
rect 13292 3476 13344 3528
rect 11529 3386 11581 3438
rect 11593 3386 11645 3438
rect 17196 3330 17248 3382
rect 17260 3330 17312 3382
rect 17196 3060 17248 3072
rect 17196 3026 17224 3060
rect 17224 3026 17248 3060
rect 17196 3020 17248 3026
rect 17260 3060 17312 3072
rect 17260 3026 17262 3060
rect 17262 3026 17296 3060
rect 17296 3026 17312 3060
rect 17260 3020 17312 3026
<< metal2 >>
rect 9831 5080 9837 5132
rect 9889 5080 9901 5132
rect 9953 5080 9959 5132
rect 7516 5046 7568 5052
rect 7516 4972 7568 4994
rect 7516 4898 7568 4920
rect 7516 4180 7568 4846
rect 9831 4760 9959 5080
rect 7516 4114 7568 4128
rect 7516 4047 7568 4062
rect 7516 3987 7568 3995
rect 8763 4683 8769 4735
rect 8821 4683 8833 4735
rect 8885 4683 8891 4735
rect 9831 4708 9837 4760
rect 9889 4708 9901 4760
rect 9953 4708 9959 4760
rect 10589 5071 10595 5123
rect 10647 5071 10659 5123
rect 10711 5071 10717 5123
rect 8763 3598 8891 4683
rect 10589 4513 10717 5071
rect 13060 4998 13066 5050
rect 13118 4998 13130 5050
rect 13182 4998 13188 5050
tri 13060 4922 13136 4998 ne
rect 10589 4461 10595 4513
rect 10647 4461 10659 4513
rect 10711 4461 10717 4513
rect 11523 4623 11529 4675
rect 11581 4623 11593 4675
rect 11645 4623 11651 4675
rect 11523 4608 11585 4623
tri 11585 4608 11600 4623 nw
rect 10272 4381 10278 4433
rect 10330 4381 10342 4433
rect 10394 4381 10400 4433
rect 10272 4195 10400 4381
rect 10272 4143 10278 4195
rect 10330 4143 10342 4195
rect 10394 4143 10400 4195
rect 8763 3546 8769 3598
rect 8821 3546 8833 3598
rect 8885 3546 8891 3598
rect 11523 3598 11575 4608
tri 11575 4598 11585 4608 nw
rect 11612 4543 11618 4595
rect 11670 4543 11682 4595
rect 11734 4543 11740 4595
tri 11663 4518 11688 4543 ne
tri 11575 3598 11600 3623 sw
rect 11523 3546 11529 3598
rect 11581 3546 11593 3598
rect 11645 3546 11651 3598
rect 11523 3543 11597 3546
tri 11597 3543 11600 3546 nw
rect 11523 3540 11594 3543
tri 11594 3540 11597 3543 nw
tri 11685 3540 11688 3543 se
rect 11688 3540 11740 4543
rect 12472 4381 12478 4433
rect 12530 4381 12542 4433
rect 12594 4381 12600 4433
rect 12472 3908 12524 4381
tri 12524 4356 12549 4381 nw
rect 13136 4195 13188 4998
rect 13216 4556 13222 4608
rect 13274 4556 13286 4608
rect 13338 4556 13344 4608
tri 13267 4531 13292 4556 ne
tri 13188 4195 13264 4271 sw
rect 13136 4143 13142 4195
rect 13194 4143 13206 4195
rect 13258 4143 13264 4195
tri 12524 3908 12549 3933 sw
rect 12472 3856 12478 3908
rect 12530 3856 12542 3908
rect 12594 3856 12600 3908
rect 11523 3528 11582 3540
tri 11582 3528 11594 3540 nw
tri 11673 3528 11685 3540 se
rect 11685 3528 11740 3540
rect 11523 3461 11575 3528
tri 11575 3521 11582 3528 nw
tri 11666 3521 11673 3528 se
rect 11673 3521 11740 3528
tri 11663 3518 11666 3521 se
rect 11666 3518 11740 3521
rect 11612 3466 11618 3518
rect 11670 3466 11682 3518
rect 11734 3466 11740 3518
rect 13292 3592 13344 4556
rect 13292 3528 13344 3540
tri 11575 3461 11577 3463 sw
rect 13292 3461 13344 3476
rect 11523 3438 11577 3461
tri 11577 3438 11600 3461 sw
rect 11523 3386 11529 3438
rect 11581 3386 11593 3438
rect 11645 3386 11651 3438
rect 17190 3330 17196 3382
rect 17248 3330 17260 3382
rect 17312 3330 17318 3382
rect 17190 3072 17318 3330
rect 17190 3020 17196 3072
rect 17248 3020 17260 3072
rect 17312 3020 17318 3072
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_0
timestamp 1666199351
transform -1 0 15232 0 1 3026
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_55959141808327  sky130_fd_io__tk_em1o_cdns_55959141808327_0
timestamp 1666199351
transform -1 0 13342 0 1 3470
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_55959141808328  sky130_fd_io__tk_em1o_cdns_55959141808328_0
timestamp 1666199351
transform 0 -1 12023 -1 0 4792
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1666199351
transform 1 0 16744 0 1 3552
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1666199351
transform 1 0 11787 0 1 4381
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1666199351
transform 1 0 11628 0 1 3386
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_0
timestamp 1666199351
transform 0 -1 12686 1 0 4032
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_1
timestamp 1666199351
transform 0 -1 13002 1 0 3881
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808134  sky130_fd_pr__nfet_01v8__example_55959141808134_0
timestamp 1666199351
transform -1 0 12901 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808304  sky130_fd_pr__nfet_01v8__example_55959141808304_0
timestamp 1666199351
transform 0 -1 12060 -1 0 4784
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_0
timestamp 1666199351
transform 1 0 13309 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_1
timestamp 1666199351
transform -1 0 13253 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_2
timestamp 1666199351
transform 1 0 12957 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_3
timestamp 1666199351
transform 1 0 12605 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808330  sky130_fd_pr__nfet_01v8__example_55959141808330_0
timestamp 1666199351
transform -1 0 12293 0 1 4573
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808330  sky130_fd_pr__nfet_01v8__example_55959141808330_1
timestamp 1666199351
transform 0 1 12406 -1 0 4804
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808331  sky130_fd_pr__nfet_01v8__example_55959141808331_0
timestamp 1666199351
transform 1 0 11581 0 1 4311
box -1 0 457 1
use sky130_fd_pr__nfet_01v8__example_55959141808332  sky130_fd_pr__nfet_01v8__example_55959141808332_0
timestamp 1666199351
transform 1 0 12093 0 1 4311
box -1 0 457 1
use sky130_fd_pr__nfet_01v8__example_55959141808333  sky130_fd_pr__nfet_01v8__example_55959141808333_0
timestamp 1666199351
transform 0 -1 12662 1 0 3225
box -1 0 801 1
use sky130_fd_pr__nfet_01v8__example_55959141808334  sky130_fd_pr__nfet_01v8__example_55959141808334_0
timestamp 1666199351
transform 0 -1 12518 -1 0 4025
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808335  sky130_fd_pr__pfet_01v8__example_55959141808335_0
timestamp 1666199351
transform -1 0 7976 0 1 3010
box -1 0 413 1
use sky130_fd_pr__pfet_01v8__example_55959141808339  sky130_fd_pr__pfet_01v8__example_55959141808339_0
timestamp 1666199351
transform -1 0 7982 0 1 4773
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808343  sky130_fd_pr__pfet_01v8__example_55959141808343_0
timestamp 1666199351
transform -1 0 17991 0 -1 4078
box -1 0 1193 1
use sky130_fd_pr__pfet_01v8__example_55959141808343  sky130_fd_pr__pfet_01v8__example_55959141808343_1
timestamp 1666199351
transform 1 0 13911 0 -1 4078
box -1 0 1193 1
use sky130_fd_pr__pfet_01v8__example_55959141808343  sky130_fd_pr__pfet_01v8__example_55959141808343_2
timestamp 1666199351
transform 1 0 15355 0 -1 4028
box -1 0 1193 1
use sky130_fd_pr__pfet_01v8__example_55959141808344  sky130_fd_pr__pfet_01v8__example_55959141808344_0
timestamp 1666199351
transform -1 0 19701 0 -1 4078
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808344  sky130_fd_pr__pfet_01v8__example_55959141808344_1
timestamp 1666199351
transform 1 0 19757 0 -1 4078
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808344  sky130_fd_pr__pfet_01v8__example_55959141808344_2
timestamp 1666199351
transform -1 0 13855 0 -1 4078
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808345  sky130_fd_pr__pfet_01v8__example_55959141808345_0
timestamp 1666199351
transform 0 -1 12990 1 0 3225
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808346  sky130_fd_pr__pfet_01v8__example_55959141808346_0
timestamp 1666199351
transform 1 0 18867 0 -1 4078
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808346  sky130_fd_pr__pfet_01v8__example_55959141808346_1
timestamp 1666199351
transform 1 0 18243 0 -1 4078
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808347  sky130_fd_pr__pfet_01v8__example_55959141808347_0
timestamp 1666199351
transform -1 0 13503 0 -1 4073
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808348  sky130_fd_pr__pfet_01v8__example_55959141808348_0
timestamp 1666199351
transform 1 0 17679 0 -1 4256
box -1 0 1601 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1666199351
transform -1 0 13392 0 -1 3976
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1666199351
transform 1 0 12299 0 -1 3429
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1666199351
transform -1 0 12674 0 1 4036
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1666199351
transform 1 0 12990 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1666199351
transform -1 0 12736 0 1 4571
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1666199351
transform 1 0 11718 0 1 4391
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1666199351
transform 1 0 12232 0 1 4387
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1666199351
transform 1 0 16368 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1666199351
transform 1 0 16056 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1666199351
transform 1 0 15744 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1666199351
transform 1 0 15432 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1666199351
transform 1 0 19796 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1666199351
transform 0 1 13710 1 0 3868
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1666199351
transform -1 0 12990 0 -1 4013
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1666199351
transform 1 0 12056 0 1 4553
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1666199351
transform 1 0 13475 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1666199351
transform 1 0 13148 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1666199351
transform 1 0 17494 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1666199351
transform 1 0 17812 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1666199351
transform 1 0 16877 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1666199351
transform 1 0 17188 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_21
timestamp 1666199351
transform 1 0 15901 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_22
timestamp 1666199351
transform 1 0 16213 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_23
timestamp 1666199351
transform 1 0 16487 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_24
timestamp 1666199351
transform 1 0 15589 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_25
timestamp 1666199351
transform 1 0 15311 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_26
timestamp 1666199351
transform 1 0 19556 0 1 3336
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_27
timestamp 1666199351
transform 1 0 18631 0 1 3422
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_28
timestamp 1666199351
transform 1 0 18320 0 1 3422
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_29
timestamp 1666199351
transform 1 0 19255 0 1 3336
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_30
timestamp 1666199351
transform 1 0 18944 0 1 3336
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_31
timestamp 1666199351
transform 1 0 18198 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_32
timestamp 1666199351
transform 1 0 18476 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_33
timestamp 1666199351
transform 1 0 19374 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_34
timestamp 1666199351
transform 1 0 19100 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_35
timestamp 1666199351
transform 1 0 18788 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_36
timestamp 1666199351
transform -1 0 12894 0 1 4559
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_37
timestamp 1666199351
transform 1 0 12014 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_38
timestamp 1666199351
transform 1 0 11548 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_39
timestamp 1666199351
transform 1 0 12488 0 1 4307
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_40
timestamp 1666199351
transform 1 0 13230 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_41
timestamp 1666199351
transform 1 0 12840 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_42
timestamp 1666199351
transform 1 0 13386 0 -1 4805
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_0
timestamp 1666199351
transform 0 1 17640 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1666199351
transform 0 -1 12402 1 0 4851
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1666199351
transform 0 -1 13226 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1666199351
transform -1 0 13332 0 1 4568
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1666199351
transform 0 -1 12338 -1 0 5441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1666199351
transform 1 0 12841 0 1 4845
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1666199351
transform 0 -1 13900 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1666199351
transform 0 -1 14836 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1666199351
transform 0 -1 14212 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1666199351
transform 0 -1 14524 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_8
timestamp 1666199351
transform 0 -1 17100 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_9
timestamp 1666199351
transform 0 -1 17412 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_10
timestamp 1666199351
transform 0 -1 19746 1 0 3638
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1666199351
transform 1 0 19591 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808291  sky130_fd_pr__via_l1m1__example_55959141808291_0
timestamp 1666199351
transform 1 0 11538 0 1 4629
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808291  sky130_fd_pr__via_l1m1__example_55959141808291_1
timestamp 1666199351
transform 1 0 11538 0 1 4771
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_0
timestamp 1666199351
transform 0 1 13498 1 0 3638
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_1
timestamp 1666199351
transform 0 1 16657 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_2
timestamp 1666199351
transform 0 1 15068 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_3
timestamp 1666199351
transform 0 1 17956 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_4
timestamp 1666199351
transform 0 -1 12994 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_0
timestamp 1666199351
transform -1 0 16515 0 1 2948
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_1
timestamp 1666199351
transform 1 0 13951 0 1 3032
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_2
timestamp 1666199351
transform -1 0 17944 0 1 3026
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808325  sky130_fd_pr__via_l1m1__example_55959141808325_0
timestamp 1666199351
transform 1 0 17719 0 1 4304
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1666199351
transform 1 0 11623 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1666199351
transform -1 0 11651 0 1 4623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1666199351
transform -1 0 11651 0 1 3546
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1666199351
transform -1 0 13344 0 1 4556
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1666199351
transform -1 0 12600 0 1 4381
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1666199351
transform -1 0 11740 0 1 3466
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1666199351
transform -1 0 11740 0 1 4543
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1666199351
transform -1 0 13264 0 1 4143
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1666199351
transform -1 0 11651 0 1 3386
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1666199351
transform 1 0 17190 0 1 3330
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1666199351
transform 0 1 13292 -1 0 3598
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1666199351
transform -1 0 17318 0 1 3020
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_11
timestamp 1666199351
transform -1 0 12600 0 1 3856
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1666199351
transform 0 -1 12293 1 0 5605
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1666199351
transform 1 0 13438 0 -1 4804
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1666199351
transform 0 -1 12739 -1 0 4279
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1666199351
transform 0 -1 12904 1 0 4543
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1666199351
transform 0 -1 13091 -1 0 4279
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1666199351
transform 0 -1 13256 1 0 4543
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1666199351
transform 0 -1 13855 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_7
timestamp 1666199351
transform 0 -1 13429 -1 0 4279
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_8
timestamp 1666199351
transform 1 0 11368 0 -1 4786
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1666199351
transform -1 0 12402 0 1 3252
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1666199351
transform 0 -1 13357 1 0 4105
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_0
timestamp 1666199351
transform 0 -1 18799 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_1
timestamp 1666199351
transform 0 -1 19423 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1666199351
transform 0 1 19583 1 0 4110
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808320  sky130_fd_pr__via_pol1__example_55959141808320_0
timestamp 1666199351
transform 0 -1 19265 -1 0 4354
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808321  sky130_fd_pr__via_pol1__example_55959141808321_0
timestamp 1666199351
transform 0 -1 15082 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808321  sky130_fd_pr__via_pol1__example_55959141808321_1
timestamp 1666199351
transform 0 -1 16527 -1 0 2996
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808321  sky130_fd_pr__via_pol1__example_55959141808321_2
timestamp 1666199351
transform 0 -1 17971 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808322  sky130_fd_pr__via_pol1__example_55959141808322_0
timestamp 1666199351
transform 0 1 11590 -1 0 4279
box 0 0 1 1
<< labels >>
flabel locali s 13805 2996 13855 3030 7 FreeSans 300 0 0 0 EN_H
port 1 nsew
flabel metal1 s 11364 4223 11400 4353 3 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 19989 4223 20025 4353 7 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 19949 3626 19985 3828 7 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 13146 4143 13191 4195 8 FreeSans 300 0 0 0 DRVLO_H_N
port 4 nsew
flabel metal1 s 11364 5251 11400 5453 3 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 11364 4839 11400 4969 3 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 13475 5251 13508 5453 7 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 13475 4839 13508 4969 7 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 19756 3100 19792 3302 7 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 11364 3100 11400 3302 3 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 11364 3626 11400 3828 3 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 11428 3856 11464 3908 3 FreeSans 300 180 0 0 PBIAS
port 5 nsew
flabel metal1 s 19927 3856 19963 3908 8 FreeSans 300 180 0 0 PBIAS
port 5 nsew
flabel metal1 s 13294 3470 13346 3514 3 FreeSans 300 270 0 0 EN_H_N
port 6 nsew
flabel metal1 s 13475 4636 13508 4682 3 FreeSans 300 0 0 0 PDEN_H_N
port 7 nsew
flabel metal1 s 12352 3401 12386 3435 7 FreeSans 300 180 0 0 PD_H
port 8 nsew
flabel comment s 13808 3895 13808 3895 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 18487 4363 18487 4363 0 FreeSans 300 0 0 0 VGND_IO
flabel comment s 17627 4233 17627 4233 0 FreeSans 300 90 0 0 VCC_IO
flabel comment s 19328 4220 19328 4220 0 FreeSans 300 90 0 0 2VTP
flabel comment s 13078 3951 13078 3951 0 FreeSans 300 90 0 0 BIAS_G
flabel comment s 12545 4128 12545 4128 0 FreeSans 300 0 0 0 M1 OPT TO BIAS_G
flabel comment s 11940 4227 11940 4227 0 FreeSans 300 0 0 0 BIAS_G
flabel comment s 12950 3166 12950 3166 0 FreeSans 300 0 0 0 VCC_IO
flabel comment s 12922 4076 12922 4076 0 FreeSans 300 0 0 0 M1 OPT TO PBIAS
flabel comment s 13215 4218 13215 4218 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 13765 4162 13765 4162 0 FreeSans 300 180 0 0 DRVLO_I_H
flabel comment s 13500 4753 13500 4753 0 FreeSans 300 90 0 0 N<1>
flabel comment s 12740 3563 12740 3563 0 FreeSans 300 180 0 0 N<0>
flabel comment s 11514 4821 11514 4821 0 FreeSans 300 180 0 0 N<1>
flabel comment s 11491 4653 11491 4653 0 FreeSans 300 180 0 0 N<0>
flabel comment s 12221 5593 12221 5593 0 FreeSans 300 0 0 0 BIAS_G
flabel comment s 12114 4991 12114 4991 0 FreeSans 300 90 0 0 NET157 OF I31
flabel comment s 11805 4403 11805 4403 0 FreeSans 300 180 0 0 M1 OPT TO PBIAS
flabel comment s 12201 4397 12201 4397 0 FreeSans 300 180 0 0 PBIAS
flabel comment s 12749 4500 12749 4500 0 FreeSans 300 180 0 0 N<1>
flabel comment s 13067 4540 13067 4540 0 FreeSans 300 270 0 0 BIAS_G
flabel comment s 13205 4614 13205 4614 0 FreeSans 300 0 0 0 EN_H_N
flabel comment s 13034 4279 13034 4279 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 12838 4609 12838 4609 0 FreeSans 300 0 0 0 PDEN_H_N
flabel comment s 14349 2974 14349 2974 0 FreeSans 300 180 0 0 PBIAS1
flabel comment s 15914 2974 15914 2974 0 FreeSans 300 180 0 0 PBIAS
flabel comment s 17404 2982 17404 2982 0 FreeSans 300 0 0 0 2VTP
flabel comment s 18516 2989 18516 2989 0 FreeSans 300 0 0 0 NET157 GT & DR TIED
flabel comment s 19133 2989 19133 2989 0 FreeSans 300 0 0 0 NET161 GT & DR TIED
flabel comment s 19723 4170 19723 4170 0 FreeSans 300 0 0 0 DRVLO_I_H
flabel comment s 19076 3586 19076 3586 0 FreeSans 300 0 0 0 NET161
flabel comment s 19225 3369 19225 3369 0 FreeSans 300 0 0 0 2VTP
flabel comment s 18593 3455 18593 3455 0 FreeSans 300 0 0 0 NET157
flabel comment s 16136 3566 16136 3566 0 FreeSans 300 180 0 0 PBIAS1
flabel comment s 13061 3380 13061 3380 0 FreeSans 300 90 0 0 BIAS_G
flabel comment s 18462 3871 18462 3871 0 FreeSans 300 180 0 0 PBIAS
flabel comment s 15965 3895 15965 3895 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 12082 3895 12082 3895 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 12105 3483 12105 3483 0 FreeSans 300 180 0 0 NET157 OF I31
<< properties >>
string GDS_END 32285534
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32244144
<< end >>
