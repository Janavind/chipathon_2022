magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 35 67 905 203
rect 35 21 789 67
rect 35 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 122 47 152 177
rect 227 47 257 177
rect 303 47 333 177
rect 418 47 448 177
rect 504 47 534 177
rect 590 47 620 177
rect 676 47 706 177
rect 778 93 808 177
<< scpmoshvt >>
rect 122 297 152 497
rect 227 297 257 497
rect 317 297 347 497
rect 418 297 448 497
rect 506 297 536 497
rect 590 297 620 497
rect 676 297 706 497
rect 778 345 808 429
<< ndiff >>
rect 61 161 122 177
rect 61 127 77 161
rect 111 127 122 161
rect 61 93 122 127
rect 61 59 77 93
rect 111 59 122 93
rect 61 47 122 59
rect 152 47 227 177
rect 257 47 303 177
rect 333 89 418 177
rect 333 55 372 89
rect 406 55 418 89
rect 333 47 418 55
rect 448 153 504 177
rect 448 119 459 153
rect 493 119 504 153
rect 448 47 504 119
rect 534 89 590 177
rect 534 55 545 89
rect 579 55 590 89
rect 534 47 590 55
rect 620 169 676 177
rect 620 135 631 169
rect 665 135 676 169
rect 620 101 676 135
rect 620 67 631 101
rect 665 67 676 101
rect 620 47 676 67
rect 706 93 778 177
rect 808 135 879 177
rect 808 101 833 135
rect 867 101 879 135
rect 808 93 879 101
rect 706 89 763 93
rect 706 55 717 89
rect 751 55 763 89
rect 706 47 763 55
<< pdiff >>
rect 56 417 122 497
rect 56 383 68 417
rect 102 383 122 417
rect 56 349 122 383
rect 56 315 68 349
rect 102 315 122 349
rect 56 297 122 315
rect 152 489 227 497
rect 152 455 176 489
rect 210 455 227 489
rect 152 297 227 455
rect 257 339 317 497
rect 257 305 272 339
rect 306 305 317 339
rect 257 297 317 305
rect 347 489 418 497
rect 347 455 365 489
rect 399 455 418 489
rect 347 297 418 455
rect 448 341 506 497
rect 448 307 461 341
rect 495 307 506 341
rect 448 297 506 307
rect 536 489 590 497
rect 536 455 546 489
rect 580 455 590 489
rect 536 297 590 455
rect 620 341 676 497
rect 620 307 631 341
rect 665 307 676 341
rect 620 297 676 307
rect 706 489 763 497
rect 706 455 717 489
rect 751 455 763 489
rect 706 429 763 455
rect 706 345 778 429
rect 808 421 865 429
rect 808 387 819 421
rect 853 387 865 421
rect 808 345 865 387
rect 706 297 763 345
<< ndiffc >>
rect 77 127 111 161
rect 77 59 111 93
rect 372 55 406 89
rect 459 119 493 153
rect 545 55 579 89
rect 631 135 665 169
rect 631 67 665 101
rect 833 101 867 135
rect 717 55 751 89
<< pdiffc >>
rect 68 383 102 417
rect 68 315 102 349
rect 176 455 210 489
rect 272 305 306 339
rect 365 455 399 489
rect 461 307 495 341
rect 546 455 580 489
rect 631 307 665 341
rect 717 455 751 489
rect 819 387 853 421
<< poly >>
rect 122 497 152 523
rect 227 497 257 523
rect 317 497 347 523
rect 418 497 448 523
rect 506 497 536 523
rect 590 497 620 523
rect 676 497 706 523
rect 778 429 808 523
rect 122 265 152 297
rect 227 265 257 297
rect 317 265 347 297
rect 418 265 448 297
rect 506 265 536 297
rect 590 265 620 297
rect 676 265 706 297
rect 778 265 808 345
rect 98 249 152 265
rect 98 215 108 249
rect 142 215 152 249
rect 98 199 152 215
rect 194 249 257 265
rect 194 215 204 249
rect 238 215 257 249
rect 194 199 257 215
rect 299 249 353 265
rect 299 215 309 249
rect 343 215 353 249
rect 299 199 353 215
rect 418 249 706 265
rect 418 215 434 249
rect 468 215 502 249
rect 536 215 570 249
rect 604 215 706 249
rect 418 199 706 215
rect 753 249 808 265
rect 753 215 763 249
rect 797 215 808 249
rect 753 199 808 215
rect 122 177 152 199
rect 227 177 257 199
rect 303 177 333 199
rect 418 177 448 199
rect 504 177 534 199
rect 590 177 620 199
rect 676 177 706 199
rect 778 177 808 199
rect 122 21 152 47
rect 227 21 257 47
rect 303 21 333 47
rect 418 21 448 47
rect 504 21 534 47
rect 590 21 620 47
rect 676 21 706 47
rect 778 27 808 93
<< polycont >>
rect 108 215 142 249
rect 204 215 238 249
rect 309 215 343 249
rect 434 215 468 249
rect 502 215 536 249
rect 570 215 604 249
rect 763 215 797 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 146 489 236 527
rect 146 455 176 489
rect 210 455 236 489
rect 349 489 415 527
rect 349 455 365 489
rect 399 455 415 489
rect 529 489 596 527
rect 529 455 546 489
rect 580 455 596 489
rect 701 489 767 527
rect 701 455 717 489
rect 751 455 767 489
rect 30 417 102 433
rect 30 383 68 417
rect 30 349 102 383
rect 30 315 68 349
rect 30 299 102 315
rect 136 387 819 421
rect 853 387 889 421
rect 136 375 889 387
rect 30 161 74 299
rect 136 265 170 375
rect 256 305 272 339
rect 306 305 411 339
rect 445 307 461 341
rect 495 307 631 341
rect 665 307 707 341
rect 377 271 411 305
rect 108 249 170 265
rect 142 215 170 249
rect 108 199 170 215
rect 204 249 247 268
rect 238 215 247 249
rect 30 127 77 161
rect 111 127 127 161
rect 204 145 247 215
rect 305 249 343 268
rect 305 215 309 249
rect 305 199 343 215
rect 377 249 620 271
rect 377 215 434 249
rect 468 215 502 249
rect 536 215 570 249
rect 604 215 620 249
rect 377 204 620 215
rect 377 161 423 204
rect 654 169 707 307
rect 30 109 127 127
rect 284 123 423 161
rect 457 153 631 169
rect 284 109 320 123
rect 30 93 320 109
rect 457 119 459 153
rect 493 135 631 153
rect 665 135 707 169
rect 493 123 707 135
rect 743 249 799 341
rect 743 215 763 249
rect 797 215 799 249
rect 743 123 799 215
rect 833 135 889 375
rect 493 119 495 123
rect 457 103 495 119
rect 30 59 77 93
rect 111 71 320 93
rect 629 101 667 123
rect 111 59 127 71
rect 30 51 127 59
rect 356 55 372 89
rect 406 55 422 89
rect 356 17 422 55
rect 529 55 545 89
rect 579 55 595 89
rect 529 17 595 55
rect 629 67 631 101
rect 665 67 667 101
rect 867 101 889 135
rect 629 51 667 67
rect 701 55 717 89
rect 751 55 767 89
rect 833 85 889 101
rect 701 17 767 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 765 221 799 255 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 673 153 707 187 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 305 221 339 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and3b_4
rlabel metal1 s 0 -48 920 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 3897976
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3891392
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 23.000 0.000 
<< end >>
