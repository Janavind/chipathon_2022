magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1907 203
rect 30 -17 64 21
<< locali >>
rect 115 323 165 425
rect 283 323 333 425
rect 115 289 341 323
rect 719 289 1159 323
rect 301 255 341 289
rect 719 265 753 289
rect 18 215 267 255
rect 301 219 649 255
rect 301 181 341 219
rect 107 145 341 181
rect 107 51 173 145
rect 275 51 341 145
rect 615 164 649 219
rect 683 199 753 265
rect 787 199 1057 255
rect 1093 215 1159 289
rect 1193 289 1653 323
rect 1193 215 1259 289
rect 1619 255 1653 289
rect 1295 215 1577 255
rect 1619 215 1915 255
rect 1102 164 1292 181
rect 615 147 1553 164
rect 615 129 1136 147
rect 1258 129 1553 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 18 459 425 493
rect 18 289 81 459
rect 199 357 249 459
rect 375 323 425 459
rect 463 443 1201 493
rect 1235 443 1637 527
rect 463 359 513 443
rect 1151 409 1201 443
rect 1671 409 1705 493
rect 547 367 1117 409
rect 547 323 606 367
rect 1151 357 1721 409
rect 1755 359 1789 527
rect 1687 323 1721 357
rect 1831 323 1881 493
rect 375 289 606 323
rect 23 17 73 179
rect 207 17 241 111
rect 375 129 581 185
rect 1687 289 1881 323
rect 1587 145 1805 181
rect 375 17 409 129
rect 547 119 581 129
rect 447 85 522 95
rect 607 85 1117 95
rect 447 51 1117 85
rect 1167 17 1201 111
rect 1587 95 1637 145
rect 1235 51 1637 95
rect 1671 17 1705 111
rect 1739 51 1805 145
rect 1839 17 1873 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 1295 215 1577 255 6 A1
port 1 nsew signal input
rlabel locali s 1619 215 1915 255 6 A2
port 2 nsew signal input
rlabel locali s 1619 255 1653 289 6 A2
port 2 nsew signal input
rlabel locali s 1193 215 1259 289 6 A2
port 2 nsew signal input
rlabel locali s 1193 289 1653 323 6 A2
port 2 nsew signal input
rlabel locali s 787 199 1057 255 6 B1
port 3 nsew signal input
rlabel locali s 1093 215 1159 289 6 B2
port 4 nsew signal input
rlabel locali s 683 199 753 265 6 B2
port 4 nsew signal input
rlabel locali s 719 265 753 289 6 B2
port 4 nsew signal input
rlabel locali s 719 289 1159 323 6 B2
port 4 nsew signal input
rlabel locali s 18 215 267 255 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1907 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1258 129 1553 147 6 Y
port 10 nsew signal output
rlabel locali s 615 129 1136 147 6 Y
port 10 nsew signal output
rlabel locali s 615 147 1553 164 6 Y
port 10 nsew signal output
rlabel locali s 1102 164 1292 181 6 Y
port 10 nsew signal output
rlabel locali s 615 164 649 219 6 Y
port 10 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 10 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 10 nsew signal output
rlabel locali s 107 145 341 181 6 Y
port 10 nsew signal output
rlabel locali s 301 181 341 219 6 Y
port 10 nsew signal output
rlabel locali s 301 219 649 255 6 Y
port 10 nsew signal output
rlabel locali s 301 255 341 289 6 Y
port 10 nsew signal output
rlabel locali s 115 289 341 323 6 Y
port 10 nsew signal output
rlabel locali s 283 323 333 425 6 Y
port 10 nsew signal output
rlabel locali s 115 323 165 425 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1932 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3687728
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3674506
<< end >>
